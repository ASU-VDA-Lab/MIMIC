module fake_jpeg_12683_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx4_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_36),
.B1(n_35),
.B2(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_48),
.B1(n_27),
.B2(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_21),
.B1(n_26),
.B2(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_16),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_31),
.B1(n_21),
.B2(n_27),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_27),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_63),
.B1(n_57),
.B2(n_59),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_51),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_72),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_23),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_51),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx11_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_56),
.B(n_67),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_78),
.B1(n_79),
.B2(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_104),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_61),
.C(n_66),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_62),
.B1(n_76),
.B2(n_73),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_76),
.B(n_94),
.C(n_90),
.D(n_92),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_110),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_41),
.C(n_65),
.Y(n_113)
);

FAx1_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_99),
.CI(n_100),
.CON(n_115),
.SN(n_115)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_112),
.B(n_107),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_53),
.B(n_56),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_119),
.A3(n_116),
.B1(n_84),
.B2(n_107),
.C1(n_82),
.C2(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_123),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_122),
.B(n_56),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_41),
.C(n_64),
.Y(n_123)
);

AOI21x1_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_43),
.B(n_10),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_4),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_10),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_125),
.Y(n_130)
);


endmodule