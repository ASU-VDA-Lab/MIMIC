module fake_netlist_6_3013_n_1872 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1872);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1872;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g177 ( 
.A(n_80),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_64),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_47),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_37),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_40),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_91),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_18),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_6),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_60),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_40),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_8),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_135),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_20),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_3),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_70),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_42),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_69),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_118),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_62),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_12),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_13),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_51),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_153),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_106),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_107),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_0),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_26),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_23),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_125),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_145),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_11),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_87),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_65),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_75),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_109),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_33),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_146),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_113),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_85),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_124),
.Y(n_253)
);

BUFx2_ASAP7_75t_SL g254 ( 
.A(n_137),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_15),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_168),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_79),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_52),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_22),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_35),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_20),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_77),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_53),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_61),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_55),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_24),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_101),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_59),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_152),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_89),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_158),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_51),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_83),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_57),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_155),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_149),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_52),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_39),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_88),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_10),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_66),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_136),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_98),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_174),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_78),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_129),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_58),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_17),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_117),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_1),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_12),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_36),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_44),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_94),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_133),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_121),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_140),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_130),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_17),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_13),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_123),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_43),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_36),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_43),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_76),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_126),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_150),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_166),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_41),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_160),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_49),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_58),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_39),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_21),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_59),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_1),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_81),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_84),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_93),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_96),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_16),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_5),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_47),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_54),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_116),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_41),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_56),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_2),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_24),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_112),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_55),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_71),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_156),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_2),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_165),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_54),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_224),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_188),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_182),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_213),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_300),
.B(n_0),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_235),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_204),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_312),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_215),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_184),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_253),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_178),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_188),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_218),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_224),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_178),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_279),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_184),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_187),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_7),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_187),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_308),
.B(n_7),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_193),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_331),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_226),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_193),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_189),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_231),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_313),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_196),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_233),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_322),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_224),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_234),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_248),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_269),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_277),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_236),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_285),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_294),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_287),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_237),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_290),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_240),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_243),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_249),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_257),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_291),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_292),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_262),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_263),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_301),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_314),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_221),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_196),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_273),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_317),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_276),
.B(n_9),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_276),
.B(n_10),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_259),
.B(n_14),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_278),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_190),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_280),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_282),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_203),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_210),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_284),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_259),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_288),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_247),
.B(n_14),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_289),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_177),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_203),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_251),
.B(n_16),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_357),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_355),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_361),
.B(n_195),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_359),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_433),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_363),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_436),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_353),
.B(n_180),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_190),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_368),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_216),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_356),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_385),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_397),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_402),
.B(n_216),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_353),
.A2(n_198),
.B(n_183),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_366),
.B(n_195),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_406),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_408),
.B(n_409),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_353),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_360),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_410),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

XNOR2x2_ASAP7_75t_L g477 ( 
.A(n_358),
.B(n_264),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_179),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_369),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_324),
.C(n_319),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_414),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_427),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_399),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_369),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_431),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_207),
.C(n_206),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_429),
.B(n_201),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_217),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_437),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_439),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_415),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_361),
.B(n_195),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_420),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_365),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_372),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_404),
.B(n_179),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_R g511 ( 
.A(n_430),
.B(n_295),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_392),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_395),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_398),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_364),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_375),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_373),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_457),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_511),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_481),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_472),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_457),
.B(n_371),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_458),
.B(n_393),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_457),
.B(n_362),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_491),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_494),
.A2(n_422),
.B1(n_424),
.B2(n_425),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_386),
.Y(n_532)
);

BUFx8_ASAP7_75t_SL g533 ( 
.A(n_444),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_472),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_478),
.B(n_370),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_381),
.C(n_377),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_455),
.B(n_412),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_481),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_491),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_443),
.B(n_422),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_494),
.A2(n_424),
.B1(n_425),
.B2(n_440),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_496),
.B(n_296),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_451),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_481),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_519),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_210),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_499),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_L g550 ( 
.A(n_493),
.B(n_419),
.C(n_387),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_481),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_499),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_500),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_451),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_500),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_455),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_471),
.B(n_210),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_501),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_464),
.B(n_432),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_455),
.B(n_297),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_501),
.Y(n_568)
);

NOR2x1p5_ASAP7_75t_L g569 ( 
.A(n_446),
.B(n_206),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_375),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_494),
.B(n_298),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_448),
.B(n_386),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_456),
.B(n_461),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_501),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_467),
.B(n_388),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_503),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_501),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_462),
.B(n_388),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_468),
.B(n_389),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_460),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_501),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_447),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_467),
.B(n_309),
.Y(n_584)
);

AND2x6_ASAP7_75t_L g585 ( 
.A(n_459),
.B(n_210),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_465),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_475),
.B(n_389),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_480),
.B(n_403),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_447),
.B(n_311),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_447),
.B(n_316),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_459),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_447),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_484),
.B(n_403),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_454),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_454),
.B(n_320),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

BUFx6f_ASAP7_75t_SL g597 ( 
.A(n_453),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_465),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_474),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_465),
.B(n_210),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_512),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_485),
.B(n_181),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_453),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_492),
.B(n_181),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_454),
.B(n_223),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_466),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_463),
.B(n_321),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_463),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_466),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_463),
.B(n_470),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_470),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_473),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_449),
.B(n_354),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_449),
.B(n_354),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_445),
.B(n_212),
.C(n_211),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_470),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_450),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_506),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_477),
.A2(n_376),
.B1(n_380),
.B2(n_254),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_450),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_509),
.B(n_352),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_476),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_518),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_498),
.B(n_185),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_504),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_502),
.B(n_185),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_479),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_482),
.Y(n_634)
);

BUFx10_ASAP7_75t_L g635 ( 
.A(n_469),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_486),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_486),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_487),
.B(n_367),
.Y(n_639)
);

INVx4_ASAP7_75t_SL g640 ( 
.A(n_487),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_488),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_488),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_489),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_489),
.B(n_186),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_490),
.A2(n_376),
.B1(n_380),
.B2(n_268),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_495),
.B(n_186),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_452),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_495),
.B(n_191),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_497),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_452),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_497),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_505),
.B(n_325),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_505),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_510),
.B(n_514),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_510),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_514),
.B(n_367),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_517),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_507),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_517),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

AND3x2_ASAP7_75t_L g663 ( 
.A(n_508),
.B(n_228),
.C(n_227),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_472),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_457),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_451),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_458),
.B(n_191),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_472),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_494),
.B(n_378),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_481),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_491),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_472),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_457),
.B(n_232),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_593),
.B(n_527),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_562),
.B(n_238),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_562),
.B(n_239),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_638),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_633),
.B(n_63),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_641),
.B(n_244),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_570),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_605),
.A2(n_539),
.B1(n_532),
.B2(n_575),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_560),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_641),
.B(n_246),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_646),
.B(n_255),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_646),
.B(n_261),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

O2A1O1Ixp5_ASAP7_75t_L g687 ( 
.A1(n_586),
.A2(n_271),
.B(n_293),
.C(n_299),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_661),
.B(n_266),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_605),
.A2(n_346),
.B1(n_333),
.B2(n_323),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_669),
.A2(n_310),
.B1(n_304),
.B2(n_224),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_650),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_601),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_560),
.B(n_413),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_654),
.B(n_223),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_669),
.A2(n_224),
.B1(n_252),
.B2(n_230),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_521),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_654),
.B(n_223),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_588),
.B(n_435),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_660),
.B(n_223),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_650),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_566),
.B(n_192),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_537),
.B(n_192),
.Y(n_702)
);

AND2x2_ASAP7_75t_SL g703 ( 
.A(n_622),
.B(n_223),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_660),
.B(n_230),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_538),
.B(n_435),
.C(n_428),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_413),
.Y(n_706)
);

AND3x1_ASAP7_75t_L g707 ( 
.A(n_550),
.B(n_428),
.C(n_426),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_532),
.A2(n_224),
.B1(n_252),
.B2(n_230),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_660),
.B(n_230),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_614),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_572),
.B(n_579),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_524),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_524),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_624),
.A2(n_241),
.B1(n_197),
.B2(n_315),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_530),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_530),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_SL g717 ( 
.A(n_630),
.B(n_340),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_539),
.B(n_416),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_580),
.B(n_587),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_614),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_633),
.B(n_230),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_536),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_630),
.B(n_194),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_539),
.B(n_426),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_667),
.B(n_194),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_543),
.B(n_200),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_536),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_584),
.B(n_200),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_522),
.B(n_202),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_633),
.B(n_252),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_586),
.B(n_224),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_618),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_664),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_636),
.B(n_252),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_664),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_618),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_625),
.B(n_416),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_625),
.B(n_423),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_636),
.B(n_252),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_570),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_636),
.B(n_268),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_525),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_521),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_SL g744 ( 
.A1(n_624),
.A2(n_342),
.B1(n_207),
.B2(n_209),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_643),
.B(n_268),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_628),
.B(n_202),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_268),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_643),
.B(n_268),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_531),
.B(n_205),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_668),
.Y(n_750)
);

AND2x2_ASAP7_75t_SL g751 ( 
.A(n_600),
.B(n_396),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_629),
.B(n_205),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_544),
.B(n_208),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_620),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_629),
.B(n_208),
.Y(n_755)
);

AOI22x1_ASAP7_75t_L g756 ( 
.A1(n_596),
.A2(n_598),
.B1(n_634),
.B2(n_632),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_551),
.B(n_332),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_668),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_632),
.B(n_332),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_634),
.A2(n_224),
.B1(n_209),
.B2(n_345),
.Y(n_760)
);

BUFx8_ASAP7_75t_L g761 ( 
.A(n_597),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_672),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_637),
.B(n_334),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_617),
.A2(n_221),
.B1(n_256),
.B2(n_347),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_528),
.B(n_334),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_637),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_642),
.B(n_335),
.Y(n_767)
);

AND2x6_ASAP7_75t_SL g768 ( 
.A(n_649),
.B(n_417),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_642),
.B(n_335),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_522),
.B(n_341),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_652),
.B(n_341),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_588),
.B(n_348),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_665),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_652),
.B(n_348),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_656),
.A2(n_339),
.B1(n_265),
.B2(n_345),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_602),
.B(n_349),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_596),
.A2(n_423),
.B(n_421),
.C(n_417),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_656),
.B(n_349),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_542),
.B(n_603),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_658),
.A2(n_330),
.B1(n_339),
.B2(n_265),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_672),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_658),
.B(n_421),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_604),
.B(n_631),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_598),
.A2(n_330),
.B1(n_343),
.B2(n_267),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_665),
.B(n_219),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_529),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_620),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_607),
.B(n_220),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_547),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_529),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_603),
.B(n_225),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_601),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_610),
.B(n_229),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_610),
.B(n_242),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_541),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_541),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_620),
.B(n_623),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_639),
.B(n_378),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_549),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_549),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_653),
.B(n_245),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_620),
.B(n_250),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_553),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_600),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_591),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_567),
.B(n_258),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_533),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_620),
.B(n_302),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_571),
.B(n_286),
.Y(n_809)
);

NAND2x1_ASAP7_75t_L g810 ( 
.A(n_546),
.B(n_384),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_655),
.B(n_303),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_623),
.B(n_305),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_623),
.B(n_283),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_553),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_671),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_671),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_591),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_673),
.A2(n_384),
.B(n_382),
.C(n_379),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_639),
.B(n_382),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_594),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_623),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_623),
.B(n_281),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_576),
.Y(n_823)
);

AND2x6_ASAP7_75t_SL g824 ( 
.A(n_657),
.B(n_379),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_592),
.B(n_260),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_645),
.B(n_275),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_609),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_644),
.B(n_274),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_554),
.A2(n_306),
.B(n_270),
.C(n_272),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_661),
.B(n_326),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_662),
.B(n_626),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_657),
.A2(n_344),
.B1(n_343),
.B2(n_329),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_540),
.B(n_267),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_SL g834 ( 
.A1(n_581),
.A2(n_344),
.B1(n_329),
.B2(n_347),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_595),
.A2(n_151),
.B(n_68),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_615),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_647),
.B(n_347),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_615),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_556),
.B(n_148),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_594),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_556),
.B(n_154),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_616),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_777),
.A2(n_548),
.B(n_616),
.C(n_608),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_797),
.A2(n_670),
.B(n_546),
.Y(n_844)
);

AND2x6_ASAP7_75t_SL g845 ( 
.A(n_702),
.B(n_576),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_711),
.B(n_559),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_703),
.A2(n_221),
.B1(n_256),
.B2(n_597),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_797),
.A2(n_546),
.B(n_565),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_789),
.B(n_626),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_742),
.B(n_561),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_751),
.A2(n_597),
.B1(n_589),
.B2(n_590),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_742),
.B(n_561),
.Y(n_852)
);

CKINVDCx6p67_ASAP7_75t_R g853 ( 
.A(n_807),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_751),
.B(n_563),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_751),
.A2(n_573),
.B1(n_569),
.B2(n_627),
.Y(n_855)
);

OAI22x1_ASAP7_75t_L g856 ( 
.A1(n_674),
.A2(n_621),
.B1(n_627),
.B2(n_599),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_721),
.A2(n_734),
.B(n_730),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_754),
.A2(n_787),
.B(n_731),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_753),
.B(n_563),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_696),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_746),
.B(n_564),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_731),
.A2(n_582),
.B(n_564),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_789),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_675),
.A2(n_582),
.B(n_554),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_710),
.B(n_555),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_L g866 ( 
.A1(n_703),
.A2(n_621),
.B(n_613),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_678),
.A2(n_552),
.B(n_565),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_701),
.B(n_662),
.C(n_663),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_804),
.A2(n_578),
.B1(n_574),
.B2(n_568),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_703),
.A2(n_574),
.B(n_578),
.C(n_555),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_676),
.A2(n_568),
.B(n_611),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_677),
.Y(n_872)
);

BUFx12f_ASAP7_75t_L g873 ( 
.A(n_761),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_710),
.B(n_640),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_795),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_792),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_678),
.A2(n_651),
.B(n_648),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_706),
.B(n_659),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_804),
.A2(n_651),
.B(n_648),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_804),
.B(n_583),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_804),
.A2(n_651),
.B(n_648),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_720),
.B(n_640),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_696),
.A2(n_651),
.B(n_648),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_743),
.A2(n_651),
.B(n_648),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_743),
.A2(n_666),
.B(n_534),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_773),
.A2(n_666),
.B(n_534),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_795),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_756),
.A2(n_545),
.B(n_557),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_756),
.A2(n_545),
.B(n_557),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_686),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_640),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_773),
.A2(n_666),
.B(n_534),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_783),
.A2(n_640),
.B1(n_583),
.B2(n_545),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_687),
.A2(n_594),
.B(n_619),
.C(n_535),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_698),
.Y(n_895)
);

OAI21xp33_ASAP7_75t_SL g896 ( 
.A1(n_732),
.A2(n_619),
.B(n_557),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_732),
.B(n_535),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_686),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_682),
.B(n_583),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_779),
.A2(n_666),
.B(n_534),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_680),
.B(n_635),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_691),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_692),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_681),
.B(n_583),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_SL g905 ( 
.A1(n_829),
.A2(n_619),
.B(n_558),
.C(n_535),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_757),
.B(n_548),
.C(n_583),
.Y(n_906)
);

O2A1O1Ixp5_ASAP7_75t_L g907 ( 
.A1(n_679),
.A2(n_558),
.B(n_585),
.C(n_606),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_836),
.A2(n_558),
.B(n_585),
.C(n_606),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_796),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_736),
.B(n_666),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_691),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_680),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_836),
.A2(n_585),
.B(n_606),
.C(n_256),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_682),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_693),
.Y(n_915)
);

O2A1O1Ixp5_ASAP7_75t_L g916 ( 
.A1(n_683),
.A2(n_585),
.B(n_606),
.C(n_534),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_821),
.A2(n_808),
.B(n_802),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_796),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_776),
.A2(n_577),
.B(n_526),
.C(n_523),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_799),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_693),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_740),
.B(n_577),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_736),
.B(n_577),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_821),
.A2(n_577),
.B(n_523),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_812),
.A2(n_577),
.B(n_523),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_801),
.A2(n_606),
.B1(n_585),
.B2(n_635),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_766),
.B(n_526),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_799),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_700),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_740),
.B(n_635),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_700),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_813),
.A2(n_526),
.B(n_523),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_766),
.B(n_526),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_765),
.B(n_526),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_800),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_806),
.A2(n_606),
.B1(n_585),
.B2(n_523),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_681),
.A2(n_612),
.B1(n_173),
.B2(n_172),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_838),
.A2(n_19),
.B(n_21),
.C(n_23),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_822),
.A2(n_612),
.B(n_170),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_739),
.A2(n_612),
.B(n_164),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_838),
.B(n_612),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_842),
.B(n_612),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_693),
.Y(n_943)
);

NOR2x1_ASAP7_75t_R g944 ( 
.A(n_823),
.B(n_19),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_817),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_791),
.B(n_25),
.C(n_26),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_698),
.B(n_25),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_706),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_807),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_842),
.B(n_161),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_772),
.B(n_27),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_718),
.B(n_28),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_718),
.B(n_28),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_800),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_724),
.B(n_29),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_724),
.B(n_159),
.Y(n_956)
);

OAI21xp33_ASAP7_75t_L g957 ( 
.A1(n_837),
.A2(n_29),
.B(n_30),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_824),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_823),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_741),
.A2(n_747),
.B(n_745),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_803),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_749),
.A2(n_111),
.B1(n_108),
.B2(n_103),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_798),
.B(n_819),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_748),
.A2(n_100),
.B(n_99),
.Y(n_964)
);

OAI21xp33_ASAP7_75t_L g965 ( 
.A1(n_775),
.A2(n_30),
.B(n_31),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_803),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_798),
.B(n_31),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_744),
.B(n_32),
.C(n_34),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_831),
.B(n_820),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_786),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_819),
.B(n_737),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_737),
.B(n_32),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_SL g973 ( 
.A1(n_744),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_717),
.A2(n_73),
.B1(n_72),
.B2(n_67),
.Y(n_974)
);

NOR2x1_ASAP7_75t_L g975 ( 
.A(n_729),
.B(n_38),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_825),
.A2(n_38),
.B(n_42),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_738),
.B(n_44),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_820),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_833),
.A2(n_45),
.B(n_46),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_785),
.A2(n_45),
.B(n_46),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_786),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_784),
.A2(n_53),
.B1(n_48),
.B2(n_50),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_684),
.A2(n_48),
.B(n_685),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_SL g984 ( 
.A(n_761),
.B(n_714),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_828),
.A2(n_717),
.B(n_752),
.C(n_763),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_840),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_738),
.B(n_755),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_834),
.B(n_770),
.C(n_689),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_793),
.B(n_726),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_759),
.A2(n_767),
.B(n_771),
.C(n_774),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_712),
.A2(n_750),
.B(n_758),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_780),
.A2(n_832),
.B(n_760),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_712),
.A2(n_750),
.B(n_758),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_840),
.A2(n_709),
.B(n_694),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_840),
.B(n_816),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_761),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_697),
.A2(n_699),
.B(n_704),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_708),
.A2(n_695),
.B1(n_778),
.B2(n_769),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_790),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_707),
.B(n_689),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_790),
.B(n_816),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_707),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_832),
.B(n_688),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_814),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_841),
.A2(n_839),
.B(n_815),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_814),
.A2(n_815),
.B(n_810),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_725),
.B(n_782),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_713),
.B(n_781),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_713),
.B(n_781),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_688),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_715),
.A2(n_733),
.B(n_762),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_728),
.A2(n_690),
.B1(n_788),
.B2(n_688),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_715),
.B(n_733),
.Y(n_1013)
);

OAI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_764),
.A2(n_705),
.B(n_723),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_827),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_810),
.A2(n_827),
.B(n_716),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_809),
.A2(n_811),
.B1(n_688),
.B2(n_794),
.Y(n_1017)
);

OAI321xp33_ASAP7_75t_L g1018 ( 
.A1(n_834),
.A2(n_826),
.A3(n_830),
.B1(n_818),
.B2(n_768),
.C(n_835),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_716),
.B(n_722),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_805),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_722),
.A2(n_727),
.B(n_735),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_762),
.B(n_805),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_805),
.A2(n_777),
.B(n_676),
.C(n_675),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_768),
.A2(n_719),
.B(n_711),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_824),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_876),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_875),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_858),
.A2(n_867),
.B(n_848),
.Y(n_1028)
);

AO21x1_ASAP7_75t_L g1029 ( 
.A1(n_950),
.A2(n_989),
.B(n_1012),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_870),
.A2(n_854),
.B(n_1023),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_990),
.B(n_864),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_887),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_857),
.A2(n_960),
.B(n_889),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1024),
.B(n_895),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_844),
.A2(n_963),
.B(n_917),
.Y(n_1035)
);

INVx3_ASAP7_75t_SL g1036 ( 
.A(n_853),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_909),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_1016),
.A2(n_994),
.B(n_888),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_919),
.A2(n_905),
.B(n_1005),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_971),
.B(n_921),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_918),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_959),
.Y(n_1042)
);

AO21x2_ASAP7_75t_L g1043 ( 
.A1(n_862),
.A2(n_997),
.B(n_871),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_894),
.A2(n_925),
.B(n_932),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_987),
.B(n_948),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_894),
.A2(n_1006),
.B(n_993),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_912),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_948),
.B(n_846),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_L g1049 ( 
.A(n_921),
.B(n_914),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_921),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_934),
.A2(n_859),
.B(n_861),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_895),
.B(n_878),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_921),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1001),
.A2(n_886),
.B(n_885),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_991),
.A2(n_1021),
.B(n_1011),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_907),
.A2(n_869),
.B(n_892),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_985),
.A2(n_943),
.B1(n_915),
.B2(n_860),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_907),
.A2(n_933),
.B(n_927),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_924),
.A2(n_916),
.B(n_877),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_998),
.A2(n_843),
.B(n_896),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_863),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_879),
.A2(n_881),
.B(n_910),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_915),
.A2(n_943),
.B1(n_860),
.B2(n_851),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_923),
.A2(n_995),
.B(n_850),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_956),
.B(n_899),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_916),
.A2(n_904),
.B(n_900),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_995),
.A2(n_852),
.B(n_969),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_969),
.A2(n_1022),
.B(n_978),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_920),
.Y(n_1069)
);

AOI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_992),
.A2(n_1014),
.B(n_951),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_904),
.A2(n_865),
.B(n_843),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_928),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_849),
.B(n_1003),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_897),
.A2(n_1009),
.B(n_1013),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_903),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_951),
.A2(n_965),
.B(n_847),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_873),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_947),
.B(n_1002),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_947),
.A2(n_957),
.B(n_982),
.C(n_988),
.Y(n_1079)
);

NAND2x1_ASAP7_75t_L g1080 ( 
.A(n_1020),
.B(n_986),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1008),
.A2(n_1019),
.B(n_874),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_914),
.B(n_899),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1002),
.B(n_912),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_906),
.A2(n_1007),
.B(n_967),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_935),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_880),
.A2(n_884),
.B(n_883),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_958),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_882),
.A2(n_891),
.B(n_942),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_855),
.A2(n_1025),
.B1(n_1000),
.B2(n_1017),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_972),
.B(n_954),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_961),
.B(n_966),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_880),
.A2(n_1020),
.B(n_941),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_872),
.A2(n_911),
.B(n_902),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_952),
.B(n_953),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_950),
.A2(n_956),
.B(n_981),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_901),
.B(n_930),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_975),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_914),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_L g1100 ( 
.A1(n_866),
.A2(n_847),
.B(n_1018),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_977),
.B(n_955),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_901),
.B(n_930),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_914),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_988),
.A2(n_938),
.B(n_968),
.C(n_946),
.Y(n_1104)
);

HAxp5_ASAP7_75t_L g1105 ( 
.A(n_973),
.B(n_968),
.CON(n_1105),
.SN(n_1105)
);

INVx5_ASAP7_75t_L g1106 ( 
.A(n_986),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_L g1107 ( 
.A1(n_982),
.A2(n_984),
.B1(n_973),
.B2(n_856),
.C(n_938),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1010),
.B(n_868),
.Y(n_1108)
);

OA22x2_ASAP7_75t_L g1109 ( 
.A1(n_974),
.A2(n_937),
.B1(n_922),
.B2(n_926),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_962),
.A2(n_983),
.B(n_976),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_R g1111 ( 
.A(n_996),
.B(n_922),
.Y(n_1111)
);

OA21x2_ASAP7_75t_L g1112 ( 
.A1(n_970),
.A2(n_1004),
.B(n_999),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_890),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_SL g1114 ( 
.A1(n_908),
.A2(n_913),
.B(n_939),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_845),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_SL g1116 ( 
.A1(n_908),
.A2(n_980),
.B(n_979),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_986),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_986),
.B(n_898),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1015),
.A2(n_929),
.B(n_931),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_893),
.B(n_936),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_944),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_913),
.B(n_940),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_964),
.B(n_711),
.Y(n_1123)
);

AOI21x1_ASAP7_75t_L g1124 ( 
.A1(n_857),
.A2(n_917),
.B(n_1016),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_878),
.B(n_849),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_963),
.B(n_711),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_853),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_858),
.A2(n_751),
.B(n_754),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_858),
.A2(n_751),
.B(n_754),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_978),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_921),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_963),
.B(n_711),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_858),
.A2(n_751),
.B(n_754),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_963),
.A2(n_804),
.B1(n_751),
.B2(n_711),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_878),
.B(n_849),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_921),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_858),
.A2(n_751),
.B(n_754),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_963),
.B(n_711),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_945),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_963),
.B(n_804),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_963),
.B(n_711),
.Y(n_1141)
);

AOI221x1_ASAP7_75t_L g1142 ( 
.A1(n_988),
.A2(n_1024),
.B1(n_985),
.B2(n_960),
.C(n_1014),
.Y(n_1142)
);

AND3x4_ASAP7_75t_L g1143 ( 
.A(n_968),
.B(n_550),
.C(n_988),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_854),
.A2(n_908),
.B(n_967),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1024),
.A2(n_719),
.B1(n_711),
.B2(n_674),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_945),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_878),
.B(n_849),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_963),
.B(n_711),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_875),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_963),
.B(n_711),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_SL g1151 ( 
.A1(n_874),
.A2(n_676),
.B(n_675),
.Y(n_1151)
);

AOI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_1024),
.A2(n_719),
.B(n_711),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_915),
.B(n_943),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_963),
.B(n_711),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_963),
.B(n_711),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_857),
.A2(n_917),
.B(n_1016),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1024),
.A2(n_719),
.B1(n_711),
.B2(n_674),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_870),
.A2(n_751),
.B(n_854),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_875),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_858),
.A2(n_751),
.B(n_754),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_L g1161 ( 
.A(n_853),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_945),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_978),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_963),
.B(n_711),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_878),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_854),
.A2(n_908),
.B(n_967),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_870),
.A2(n_751),
.B(n_854),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_857),
.A2(n_960),
.B(n_889),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_870),
.A2(n_751),
.B(n_854),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_857),
.A2(n_960),
.B(n_889),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_857),
.A2(n_917),
.B(n_1016),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_876),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_971),
.A2(n_963),
.B1(n_605),
.B2(n_948),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1026),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_1165),
.B(n_1075),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1143),
.A2(n_1076),
.B1(n_1100),
.B2(n_1070),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_1127),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1027),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1090),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1172),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1028),
.A2(n_1051),
.B(n_1035),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1053),
.B(n_1106),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1123),
.A2(n_1129),
.B(n_1128),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1152),
.B(n_1138),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1050),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1141),
.B(n_1148),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1053),
.B(n_1106),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1032),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_1049),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1150),
.B(n_1154),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1133),
.A2(n_1160),
.B(n_1137),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1037),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_1155),
.B1(n_1164),
.B2(n_1145),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1079),
.A2(n_1104),
.B(n_1105),
.C(n_1173),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1090),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1031),
.A2(n_1043),
.B(n_1062),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1122),
.A2(n_1060),
.B(n_1034),
.C(n_1084),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1157),
.B(n_1142),
.C(n_1107),
.Y(n_1200)
);

AOI222xp33_ASAP7_75t_L g1201 ( 
.A1(n_1105),
.A2(n_1078),
.B1(n_1165),
.B2(n_1073),
.C1(n_1045),
.C2(n_1089),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_L g1202 ( 
.A(n_1050),
.B(n_1131),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1054),
.A2(n_1096),
.B(n_1081),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1061),
.B(n_1052),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1034),
.B(n_1101),
.C(n_1095),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1047),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1147),
.B(n_1097),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1029),
.A2(n_1068),
.B(n_1030),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1041),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1069),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1064),
.A2(n_1067),
.B(n_1170),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1127),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1048),
.B(n_1134),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1091),
.A2(n_1108),
.B1(n_1042),
.B2(n_1098),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1033),
.A2(n_1168),
.B(n_1170),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1072),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1047),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1065),
.B(n_1103),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1065),
.B(n_1083),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1085),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1143),
.A2(n_1092),
.B1(n_1149),
.B2(n_1159),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1102),
.B(n_1065),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1153),
.B(n_1099),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1053),
.B(n_1106),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1117),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1161),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1117),
.Y(n_1227)
);

AO22x1_ASAP7_75t_L g1228 ( 
.A1(n_1115),
.A2(n_1036),
.B1(n_1153),
.B2(n_1077),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1036),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1161),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1153),
.B(n_1082),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_SL g1232 ( 
.A(n_1121),
.B(n_1087),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1077),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1173),
.A2(n_1116),
.B(n_1040),
.C(n_1144),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1140),
.B(n_1040),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1158),
.B(n_1167),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1109),
.A2(n_1110),
.B1(n_1140),
.B2(n_1063),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1111),
.B(n_1087),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1082),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1131),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1106),
.B(n_1099),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1109),
.A2(n_1166),
.B1(n_1169),
.B2(n_1122),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1113),
.B(n_1146),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1113),
.B(n_1146),
.Y(n_1244)
);

AO22x1_ASAP7_75t_L g1245 ( 
.A1(n_1131),
.A2(n_1136),
.B1(n_1118),
.B2(n_1057),
.Y(n_1245)
);

NOR2x1_ASAP7_75t_L g1246 ( 
.A(n_1049),
.B(n_1118),
.Y(n_1246)
);

CKINVDCx8_ASAP7_75t_R g1247 ( 
.A(n_1131),
.Y(n_1247)
);

INVx3_ASAP7_75t_SL g1248 ( 
.A(n_1136),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1120),
.A2(n_1130),
.B1(n_1163),
.B2(n_1136),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1139),
.B(n_1162),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1136),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1118),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1121),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1071),
.A2(n_1088),
.B(n_1066),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1080),
.Y(n_1255)
);

INVx8_ASAP7_75t_L g1256 ( 
.A(n_1130),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1163),
.Y(n_1257)
);

NOR2xp67_ASAP7_75t_L g1258 ( 
.A(n_1119),
.B(n_1171),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1071),
.A2(n_1039),
.B1(n_1112),
.B2(n_1093),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1112),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1039),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1094),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1086),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1066),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1074),
.B(n_1055),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1059),
.B(n_1058),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1151),
.B(n_1114),
.C(n_1058),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1038),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1059),
.B(n_1056),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1056),
.A2(n_1046),
.B(n_1044),
.C(n_1114),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1028),
.A2(n_1051),
.B(n_1035),
.Y(n_1271)
);

CKINVDCx8_ASAP7_75t_R g1272 ( 
.A(n_1042),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1152),
.B(n_711),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1027),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1026),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1065),
.B(n_1082),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1143),
.A2(n_1076),
.B1(n_1024),
.B2(n_1100),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1027),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1053),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1028),
.A2(n_1051),
.B(n_1035),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1053),
.Y(n_1284)
);

AND2x2_ASAP7_75t_SL g1285 ( 
.A(n_1107),
.B(n_703),
.Y(n_1285)
);

OR2x6_ASAP7_75t_L g1286 ( 
.A(n_1065),
.B(n_1082),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1028),
.A2(n_1051),
.B(n_1035),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1042),
.Y(n_1288)
);

INVx8_ASAP7_75t_L g1289 ( 
.A(n_1053),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1026),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1079),
.A2(n_703),
.B1(n_1132),
.B2(n_1126),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1165),
.B(n_789),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1065),
.B(n_1103),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1152),
.A2(n_674),
.B(n_1024),
.C(n_719),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1027),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1027),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1026),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1073),
.A2(n_984),
.B1(n_831),
.B2(n_711),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_1165),
.B(n_789),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1052),
.B(n_581),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1026),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1065),
.B(n_1103),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1127),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1026),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1042),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1134),
.A2(n_804),
.B(n_1128),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1065),
.B(n_1082),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1065),
.B(n_1103),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1027),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1065),
.B(n_1103),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1028),
.A2(n_1051),
.B(n_1035),
.Y(n_1312)
);

O2A1O1Ixp5_ASAP7_75t_SL g1313 ( 
.A1(n_1100),
.A2(n_1070),
.B(n_1152),
.C(n_1140),
.Y(n_1313)
);

BUFx4f_ASAP7_75t_SL g1314 ( 
.A(n_1127),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1090),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1143),
.A2(n_719),
.B1(n_711),
.B2(n_1024),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1212),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1184),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1316),
.A2(n_1273),
.B1(n_1299),
.B2(n_1285),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1186),
.A2(n_1188),
.B1(n_1177),
.B2(n_1280),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1201),
.B(n_1195),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1192),
.A2(n_1297),
.B1(n_1175),
.B2(n_1191),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1179),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1178),
.A2(n_1272),
.B1(n_1233),
.B2(n_1314),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1190),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1194),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1209),
.Y(n_1327)
);

BUFx8_ASAP7_75t_SL g1328 ( 
.A(n_1288),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1210),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1289),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1216),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1220),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1276),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1304),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1276),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1289),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1260),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1275),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1281),
.Y(n_1339)
);

AO21x1_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1208),
.B(n_1291),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1246),
.B(n_1262),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1200),
.A2(n_1291),
.B1(n_1195),
.B2(n_1236),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1243),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1306),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1295),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1200),
.A2(n_1236),
.B1(n_1297),
.B2(n_1192),
.Y(n_1346)
);

CKINVDCx6p67_ASAP7_75t_R g1347 ( 
.A(n_1226),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1244),
.Y(n_1348)
);

BUFx2_ASAP7_75t_R g1349 ( 
.A(n_1253),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1201),
.B(n_1222),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1189),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1296),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1240),
.Y(n_1353)
);

INVx6_ASAP7_75t_L g1354 ( 
.A(n_1240),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1240),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1207),
.B(n_1180),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_SL g1357 ( 
.A(n_1294),
.B(n_1199),
.C(n_1205),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1181),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1205),
.A2(n_1221),
.B1(n_1279),
.B2(n_1278),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1274),
.B(n_1301),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1298),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1310),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1213),
.B(n_1235),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1242),
.B(n_1231),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1221),
.A2(n_1219),
.B1(n_1229),
.B2(n_1302),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1219),
.A2(n_1292),
.B1(n_1300),
.B2(n_1204),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1197),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1250),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1206),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1270),
.A2(n_1185),
.B(n_1193),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1225),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1251),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1227),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1203),
.A2(n_1271),
.B(n_1283),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1227),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1217),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1183),
.A2(n_1287),
.B(n_1312),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1268),
.Y(n_1379)
);

AOI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1245),
.A2(n_1258),
.B(n_1211),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1315),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1313),
.A2(n_1234),
.B(n_1249),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1254),
.A2(n_1263),
.B(n_1265),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1229),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1265),
.Y(n_1385)
);

INVxp33_ASAP7_75t_L g1386 ( 
.A(n_1182),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1176),
.A2(n_1302),
.B1(n_1290),
.B2(n_1237),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1305),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1269),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1218),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1266),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1239),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1202),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1252),
.B(n_1277),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1224),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1254),
.A2(n_1263),
.B(n_1264),
.Y(n_1396)
);

OAI22x1_ASAP7_75t_L g1397 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1267),
.B2(n_1266),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1218),
.A2(n_1293),
.B1(n_1303),
.B2(n_1309),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1187),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1261),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1257),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1257),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1257),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1293),
.A2(n_1311),
.B1(n_1309),
.B2(n_1303),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1267),
.A2(n_1307),
.B(n_1249),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1311),
.B(n_1223),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1252),
.B(n_1308),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1238),
.A2(n_1230),
.B1(n_1256),
.B2(n_1282),
.Y(n_1408)
);

INVx4_ASAP7_75t_SL g1409 ( 
.A(n_1277),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1286),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1187),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1241),
.A2(n_1255),
.B(n_1256),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1187),
.Y(n_1413)
);

INVx4_ASAP7_75t_SL g1414 ( 
.A(n_1286),
.Y(n_1414)
);

BUFx8_ASAP7_75t_L g1415 ( 
.A(n_1223),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1247),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1256),
.A2(n_1284),
.B1(n_1286),
.B2(n_1308),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1308),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1228),
.A2(n_1241),
.B(n_1284),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1248),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1232),
.B(n_1188),
.Y(n_1421)
);

AO21x1_ASAP7_75t_L g1422 ( 
.A1(n_1196),
.A2(n_1100),
.B(n_1208),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1273),
.B(n_355),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1191),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1215),
.A2(n_1156),
.B(n_1124),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1285),
.A2(n_984),
.B1(n_1273),
.B2(n_831),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1181),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1276),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1206),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1174),
.Y(n_1430)
);

BUFx8_ASAP7_75t_L g1431 ( 
.A(n_1182),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1270),
.A2(n_1185),
.B(n_1198),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1174),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1215),
.A2(n_1156),
.B(n_1124),
.Y(n_1434)
);

BUFx2_ASAP7_75t_SL g1435 ( 
.A(n_1240),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1177),
.B(n_1280),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1382),
.A2(n_1375),
.B(n_1378),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1321),
.B(n_1365),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1321),
.B(n_1365),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1328),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1376),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1376),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1379),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1385),
.B(n_1364),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1320),
.B(n_1322),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1429),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1364),
.B(n_1357),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1396),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1317),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1429),
.Y(n_1450)
);

INVx5_ASAP7_75t_SL g1451 ( 
.A(n_1347),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1436),
.B(n_1369),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1354),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1405),
.B(n_1340),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1400),
.B(n_1361),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1342),
.B(n_1350),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1426),
.A2(n_1423),
.B(n_1319),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1409),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1409),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1391),
.B(n_1337),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1380),
.A2(n_1397),
.B(n_1422),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1337),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1354),
.Y(n_1463)
);

INVxp67_ASAP7_75t_R g1464 ( 
.A(n_1324),
.Y(n_1464)
);

AOI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1422),
.A2(n_1434),
.B(n_1425),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1421),
.A2(n_1346),
.B(n_1424),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1391),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1389),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1389),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1362),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1328),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1360),
.B(n_1386),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1340),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1396),
.A2(n_1383),
.B(n_1345),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1341),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1350),
.B(n_1343),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1383),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1436),
.B(n_1356),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1323),
.Y(n_1479)
);

AOI21xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1317),
.A2(n_1334),
.B(n_1387),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1341),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1325),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1326),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1327),
.A2(n_1363),
.B(n_1338),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1359),
.A2(n_1366),
.B(n_1367),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1341),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1415),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1329),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1348),
.B(n_1331),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1430),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1332),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1339),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1352),
.A2(n_1418),
.B(n_1410),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1354),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1433),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1410),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1418),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1371),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1394),
.B(n_1407),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1432),
.A2(n_1412),
.B(n_1419),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1333),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1374),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1335),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1394),
.B(n_1407),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1355),
.A2(n_1393),
.B(n_1330),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1409),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1334),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1409),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1370),
.B(n_1372),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1414),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1388),
.B(n_1373),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1388),
.B(n_1428),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1419),
.A2(n_1392),
.B(n_1412),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1502),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1450),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1448),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1447),
.B(n_1377),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1447),
.B(n_1420),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1445),
.B(n_1386),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1457),
.A2(n_1456),
.B1(n_1486),
.B2(n_1478),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1476),
.B(n_1414),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1494),
.B(n_1420),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1443),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1448),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1472),
.B(n_1384),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1494),
.B(n_1384),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1448),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1476),
.B(n_1414),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1494),
.B(n_1414),
.Y(n_1530)
);

BUFx2_ASAP7_75t_SL g1531 ( 
.A(n_1488),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1448),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1494),
.B(n_1403),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1454),
.B(n_1390),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1475),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1454),
.B(n_1399),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1467),
.B(n_1401),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1467),
.B(n_1402),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1454),
.B(n_1413),
.Y(n_1540)
);

OAI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1456),
.A2(n_1408),
.B(n_1349),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1470),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1485),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1454),
.B(n_1411),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1441),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1465),
.A2(n_1416),
.B(n_1406),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_1431),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1454),
.B(n_1435),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1504),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1496),
.B(n_1431),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1469),
.B(n_1417),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1482),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1500),
.B(n_1318),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1482),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1500),
.B(n_1395),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1505),
.B(n_1395),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1444),
.B(n_1368),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1450),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1507),
.B(n_1509),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1479),
.B(n_1351),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1542),
.B(n_1442),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1518),
.B(n_1446),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1518),
.B(n_1503),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1545),
.B(n_1503),
.Y(n_1564)
);

NAND4xp25_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_1452),
.C(n_1466),
.D(n_1512),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1533),
.B(n_1474),
.Y(n_1566)
);

OAI21xp33_ASAP7_75t_L g1567 ( 
.A1(n_1521),
.A2(n_1480),
.B(n_1439),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1533),
.B(n_1474),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1455),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1519),
.B(n_1455),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1557),
.B(n_1512),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1557),
.B(n_1444),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1527),
.B(n_1480),
.C(n_1473),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1541),
.A2(n_1513),
.B1(n_1404),
.B2(n_1398),
.C(n_1488),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1520),
.B(n_1513),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1527),
.B(n_1473),
.C(n_1487),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1522),
.A2(n_1439),
.B1(n_1438),
.B2(n_1459),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1526),
.B(n_1449),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1536),
.B(n_1479),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1530),
.B(n_1477),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1483),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1483),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1522),
.B(n_1458),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1529),
.A2(n_1438),
.B1(n_1459),
.B2(n_1458),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1534),
.B(n_1487),
.C(n_1462),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1541),
.A2(n_1511),
.B(n_1509),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1530),
.B(n_1477),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1547),
.A2(n_1451),
.B1(n_1488),
.B2(n_1464),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1550),
.A2(n_1506),
.B(n_1514),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1515),
.B(n_1449),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1524),
.B(n_1497),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1539),
.B(n_1516),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1524),
.B(n_1497),
.Y(n_1593)
);

AOI211xp5_ASAP7_75t_L g1594 ( 
.A1(n_1537),
.A2(n_1464),
.B(n_1506),
.C(n_1510),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1549),
.B(n_1487),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1534),
.B(n_1508),
.C(n_1471),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1537),
.B(n_1487),
.C(n_1462),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1539),
.B(n_1484),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1543),
.A2(n_1501),
.B(n_1499),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1523),
.B(n_1510),
.C(n_1484),
.D(n_1489),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_L g1601 ( 
.A(n_1540),
.B(n_1487),
.C(n_1481),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1540),
.A2(n_1481),
.B(n_1460),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1516),
.B(n_1489),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1558),
.B(n_1492),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1551),
.A2(n_1493),
.B1(n_1492),
.B2(n_1490),
.C(n_1560),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1553),
.B(n_1498),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1553),
.B(n_1555),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1555),
.B(n_1461),
.Y(n_1608)
);

OAI21xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1529),
.A2(n_1459),
.B(n_1458),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1544),
.B(n_1437),
.C(n_1468),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1544),
.A2(n_1514),
.B(n_1501),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1567),
.A2(n_1551),
.B1(n_1559),
.B2(n_1531),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1591),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1567),
.A2(n_1559),
.B1(n_1531),
.B2(n_1556),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1591),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1599),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1607),
.B(n_1548),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1607),
.B(n_1548),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1599),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1548),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1608),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1593),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1563),
.B(n_1523),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1580),
.B(n_1548),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1562),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1587),
.B(n_1608),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1587),
.B(n_1548),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1573),
.A2(n_1546),
.B(n_1490),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1566),
.B(n_1546),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1517),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1568),
.B(n_1517),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1599),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1564),
.B(n_1535),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1568),
.B(n_1517),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1569),
.B(n_1535),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1594),
.B(n_1451),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1570),
.B(n_1546),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1571),
.B(n_1552),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1579),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1581),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1592),
.B(n_1552),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1582),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1572),
.B(n_1554),
.Y(n_1645)
);

NAND2x1p5_ASAP7_75t_SL g1646 ( 
.A(n_1595),
.B(n_1453),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1606),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1595),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1603),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1604),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1597),
.B(n_1525),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1652),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1617),
.B(n_1609),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1618),
.B(n_1621),
.Y(n_1656)
);

OR2x6_ASAP7_75t_L g1657 ( 
.A(n_1648),
.B(n_1459),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1629),
.B(n_1600),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1650),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1618),
.B(n_1609),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1626),
.B(n_1525),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1626),
.B(n_1525),
.Y(n_1662)
);

OAI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1625),
.A2(n_1586),
.B1(n_1565),
.B2(n_1588),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1619),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1652),
.B(n_1610),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1649),
.B(n_1578),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1650),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1630),
.B(n_1525),
.Y(n_1668)
);

INVxp33_ASAP7_75t_L g1669 ( 
.A(n_1649),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1528),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1628),
.B(n_1576),
.C(n_1561),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1651),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1651),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1613),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1623),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1613),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1632),
.B(n_1528),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1612),
.A2(n_1574),
.B1(n_1596),
.B2(n_1577),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1629),
.B(n_1638),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1632),
.B(n_1528),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1615),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1615),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1619),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1622),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1622),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1635),
.B(n_1528),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1635),
.B(n_1532),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1652),
.B(n_1611),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_SL g1690 ( 
.A(n_1648),
.B(n_1585),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1652),
.B(n_1620),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1658),
.B(n_1623),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1659),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1658),
.B(n_1636),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1657),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1666),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1691),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1664),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1659),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1655),
.B(n_1620),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1676),
.B(n_1636),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1676),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1655),
.B(n_1624),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1691),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1663),
.B(n_1640),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1660),
.B(n_1624),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1664),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1672),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1690),
.C(n_1675),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1639),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1680),
.B(n_1639),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1660),
.B(n_1627),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1672),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1653),
.B(n_1627),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1653),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1680),
.B(n_1645),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1673),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1669),
.B(n_1671),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1673),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1674),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1674),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1664),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_SL g1725 ( 
.A(n_1679),
.B(n_1614),
.C(n_1654),
.D(n_1628),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1657),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1653),
.B(n_1440),
.Y(n_1727)
);

NOR2xp67_ASAP7_75t_L g1728 ( 
.A(n_1665),
.B(n_1647),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1602),
.C(n_1584),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1679),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1665),
.B(n_1640),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1677),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1665),
.B(n_1641),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1697),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1691),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1702),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1717),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1696),
.B(n_1344),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1698),
.Y(n_1740)
);

BUFx4_ASAP7_75t_SL g1741 ( 
.A(n_1711),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1706),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1700),
.B(n_1691),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1706),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1701),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1707),
.Y(n_1746)
);

CKINVDCx16_ASAP7_75t_R g1747 ( 
.A(n_1727),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1730),
.B(n_1656),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1694),
.B(n_1682),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1697),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1705),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1703),
.B(n_1654),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1703),
.B(n_1665),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1694),
.B(n_1682),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1707),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1720),
.B(n_1656),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1701),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1712),
.B(n_1689),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1708),
.B(n_1714),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1708),
.B(n_1689),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1714),
.B(n_1689),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1725),
.B(n_1344),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1722),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1712),
.B(n_1689),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1723),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1692),
.B(n_1683),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1698),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1692),
.B(n_1683),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1729),
.B(n_1631),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1728),
.B(n_1657),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1733),
.B(n_1731),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1748),
.B(n_1713),
.Y(n_1772)
);

OAI31xp33_ASAP7_75t_L g1773 ( 
.A1(n_1762),
.A2(n_1704),
.A3(n_1695),
.B(n_1716),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1716),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_SL g1775 ( 
.A(n_1741),
.B(n_1695),
.C(n_1713),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1735),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1751),
.A2(n_1704),
.B(n_1590),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1750),
.B(n_1726),
.Y(n_1778)
);

NOR3xp33_ASAP7_75t_L g1779 ( 
.A(n_1747),
.B(n_1726),
.C(n_1699),
.Y(n_1779)
);

AOI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1735),
.A2(n_1710),
.B(n_1693),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1737),
.A2(n_1715),
.B1(n_1721),
.B2(n_1719),
.C(n_1726),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1756),
.A2(n_1718),
.B1(n_1657),
.B2(n_1732),
.C(n_1734),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1745),
.Y(n_1783)
);

AOI321xp33_ASAP7_75t_L g1784 ( 
.A1(n_1737),
.A2(n_1718),
.A3(n_1724),
.B1(n_1709),
.B2(n_1684),
.C(n_1631),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1757),
.B(n_1738),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1759),
.B(n_1685),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1759),
.B(n_1685),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1739),
.A2(n_1358),
.B1(n_1427),
.B2(n_1381),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1752),
.B(n_1758),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1742),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1764),
.B(n_1634),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1750),
.A2(n_1657),
.B1(n_1634),
.B2(n_1645),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1742),
.Y(n_1793)
);

NOR2x1_ASAP7_75t_L g1794 ( 
.A(n_1763),
.B(n_1709),
.Y(n_1794)
);

NAND2x1_ASAP7_75t_L g1795 ( 
.A(n_1770),
.B(n_1724),
.Y(n_1795)
);

OR4x1_ASAP7_75t_L g1796 ( 
.A(n_1763),
.B(n_1765),
.C(n_1746),
.D(n_1744),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1785),
.B(n_1752),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1783),
.B(n_1765),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1776),
.B(n_1753),
.Y(n_1799)
);

NAND2x1_ASAP7_75t_SL g1800 ( 
.A(n_1774),
.B(n_1770),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1790),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1789),
.B(n_1766),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1777),
.B(n_1753),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1775),
.B(n_1788),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1779),
.A2(n_1743),
.B1(n_1736),
.B2(n_1760),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1788),
.B(n_1736),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1793),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_L g1808 ( 
.A(n_1794),
.B(n_1744),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1796),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1780),
.Y(n_1810)
);

NOR3xp33_ASAP7_75t_L g1811 ( 
.A(n_1781),
.B(n_1755),
.C(n_1746),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1772),
.B(n_1755),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1784),
.B(n_1768),
.C(n_1766),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1786),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1787),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1778),
.Y(n_1816)
);

NAND4xp75_ASAP7_75t_L g1817 ( 
.A(n_1808),
.B(n_1773),
.C(n_1771),
.D(n_1784),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1797),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1806),
.B(n_1792),
.Y(n_1819)
);

NOR3x1_ASAP7_75t_L g1820 ( 
.A(n_1816),
.B(n_1782),
.C(n_1795),
.Y(n_1820)
);

AOI211xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1809),
.A2(n_1804),
.B(n_1810),
.C(n_1811),
.Y(n_1821)
);

AOI322xp5_ASAP7_75t_L g1822 ( 
.A1(n_1803),
.A2(n_1761),
.A3(n_1760),
.B1(n_1743),
.B2(n_1778),
.C1(n_1770),
.C2(n_1740),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1800),
.Y(n_1823)
);

A2O1A1Ixp33_ASAP7_75t_SL g1824 ( 
.A1(n_1801),
.A2(n_1767),
.B(n_1740),
.C(n_1761),
.Y(n_1824)
);

AOI311xp33_ASAP7_75t_L g1825 ( 
.A1(n_1814),
.A2(n_1686),
.A3(n_1791),
.B(n_1641),
.C(n_1644),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1815),
.B(n_1768),
.Y(n_1826)
);

OAI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1805),
.A2(n_1770),
.B(n_1754),
.Y(n_1827)
);

AOI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1813),
.A2(n_1754),
.B(n_1749),
.C(n_1767),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1823),
.A2(n_1798),
.B(n_1799),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_L g1830 ( 
.A(n_1817),
.B(n_1807),
.Y(n_1830)
);

NOR2xp67_ASAP7_75t_L g1831 ( 
.A(n_1818),
.B(n_1802),
.Y(n_1831)
);

NOR3x1_ASAP7_75t_L g1832 ( 
.A(n_1819),
.B(n_1798),
.C(n_1812),
.Y(n_1832)
);

AOI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1824),
.A2(n_1812),
.B(n_1749),
.C(n_1767),
.Y(n_1833)
);

NOR3x1_ASAP7_75t_L g1834 ( 
.A(n_1821),
.B(n_1686),
.C(n_1347),
.Y(n_1834)
);

NAND4xp25_ASAP7_75t_L g1835 ( 
.A(n_1821),
.B(n_1820),
.C(n_1828),
.D(n_1822),
.Y(n_1835)
);

AO22x2_ASAP7_75t_L g1836 ( 
.A1(n_1825),
.A2(n_1740),
.B1(n_1684),
.B2(n_1368),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1827),
.B(n_1358),
.Y(n_1837)
);

NOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1826),
.B(n_1381),
.Y(n_1838)
);

AOI22x1_ASAP7_75t_SL g1839 ( 
.A1(n_1818),
.A2(n_1431),
.B1(n_1684),
.B2(n_1451),
.Y(n_1839)
);

NAND5xp2_ASAP7_75t_L g1840 ( 
.A(n_1821),
.B(n_1451),
.C(n_1507),
.D(n_1511),
.E(n_1461),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1833),
.B(n_1451),
.C(n_1583),
.Y(n_1841)
);

AOI221xp5_ASAP7_75t_SL g1842 ( 
.A1(n_1835),
.A2(n_1661),
.B1(n_1662),
.B2(n_1681),
.C(n_1678),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_SL g1843 ( 
.A(n_1837),
.B(n_1583),
.C(n_1642),
.Y(n_1843)
);

AOI222xp33_ASAP7_75t_L g1844 ( 
.A1(n_1830),
.A2(n_1631),
.B1(n_1643),
.B2(n_1616),
.C1(n_1619),
.C2(n_1633),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1831),
.A2(n_1427),
.B(n_1668),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1838),
.B(n_1644),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1842),
.B(n_1832),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1845),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1846),
.A2(n_1839),
.B1(n_1836),
.B2(n_1829),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1843),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1841),
.A2(n_1836),
.B1(n_1834),
.B2(n_1840),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1844),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1848),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1850),
.B(n_1661),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1847),
.A2(n_1330),
.B(n_1336),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1852),
.B(n_1662),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_SL g1857 ( 
.A1(n_1851),
.A2(n_1849),
.B(n_1643),
.C(n_1616),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1853),
.B(n_1435),
.Y(n_1858)
);

AO22x2_ASAP7_75t_L g1859 ( 
.A1(n_1854),
.A2(n_1616),
.B1(n_1643),
.B2(n_1633),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1856),
.B(n_1854),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1855),
.B1(n_1857),
.B2(n_1631),
.Y(n_1861)
);

XNOR2xp5_ASAP7_75t_L g1862 ( 
.A(n_1861),
.B(n_1858),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1862),
.Y(n_1863)
);

AO22x2_ASAP7_75t_L g1864 ( 
.A1(n_1862),
.A2(n_1859),
.B1(n_1616),
.B2(n_1643),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1863),
.A2(n_1688),
.B(n_1670),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1864),
.B(n_1668),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1866),
.A2(n_1336),
.B(n_1353),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1865),
.B(n_1353),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1868),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1869),
.Y(n_1870)
);

OAI221xp5_ASAP7_75t_R g1871 ( 
.A1(n_1870),
.A2(n_1867),
.B1(n_1646),
.B2(n_1354),
.C(n_1687),
.Y(n_1871)
);

AOI211xp5_ASAP7_75t_L g1872 ( 
.A1(n_1871),
.A2(n_1463),
.B(n_1495),
.C(n_1453),
.Y(n_1872)
);


endmodule