module fake_jpeg_27585_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_22),
.Y(n_24)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_16),
.B1(n_12),
.B2(n_13),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_16),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_12),
.B(n_17),
.C(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_14),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_10),
.B(n_9),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_23),
.B1(n_28),
.B2(n_5),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_35),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_31),
.B1(n_32),
.B2(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_42),
.C(n_48),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_29),
.B1(n_2),
.B2(n_6),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_42),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_47),
.C(n_6),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_55),
.C(n_44),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_4),
.B1(n_43),
.B2(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);


endmodule