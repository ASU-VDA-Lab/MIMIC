module fake_jpeg_26547_n_64 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

INVx4_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_20),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_10),
.C(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_54),
.B(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_12),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_13),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_49),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_48),
.B(n_57),
.Y(n_63)
);

OAI31xp33_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_51),
.A3(n_17),
.B(n_19),
.Y(n_64)
);


endmodule