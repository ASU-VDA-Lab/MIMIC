module fake_aes_11232_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_7), .B(n_4), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_15), .B(n_0), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVxp67_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
OA21x2_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_14), .B(n_13), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_17), .A2(n_16), .B1(n_2), .B2(n_3), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_21), .B(n_17), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_19), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_24), .B(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_27), .Y(n_28) );
OAI32xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_20), .A3(n_18), .B1(n_16), .B2(n_25), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_26), .B(n_25), .Y(n_30) );
XNOR2x1_ASAP7_75t_L g31 ( .A(n_29), .B(n_24), .Y(n_31) );
OAI21xp5_ASAP7_75t_L g32 ( .A1(n_28), .A2(n_25), .B(n_24), .Y(n_32) );
INVxp67_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_30), .B(n_25), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
OR5x1_ASAP7_75t_L g36 ( .A(n_33), .B(n_1), .C(n_2), .D(n_3), .E(n_5), .Y(n_36) );
AOI22x1_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_24), .B1(n_1), .B2(n_22), .Y(n_37) );
OAI21xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_34), .B(n_24), .Y(n_38) );
AOI22x1_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_36), .B1(n_8), .B2(n_9), .Y(n_39) );
endmodule