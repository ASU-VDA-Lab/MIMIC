module fake_ariane_1776_n_1979 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1979);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1979;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g191 ( 
.A(n_64),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_35),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_49),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_125),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_37),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_85),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_91),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_113),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_84),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_29),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_156),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_15),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_43),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_108),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_63),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_56),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_58),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_80),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_133),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_71),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_163),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_70),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_82),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_50),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_22),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_137),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_65),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_78),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_28),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_86),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_97),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_185),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_30),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_53),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_130),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_183),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_101),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_144),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_59),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_29),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_73),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_53),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_123),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_79),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_36),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_61),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_117),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_83),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_52),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_120),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_72),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_160),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_127),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_105),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_161),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_175),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_81),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_149),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_159),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_1),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_112),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_138),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_28),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_1),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_166),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_140),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_162),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_42),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_48),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_164),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_65),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_189),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_99),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_44),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_56),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_184),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_109),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_93),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_176),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_141),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_88),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_168),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_4),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_50),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_119),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_19),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_32),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_173),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_147),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_17),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_136),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_107),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_32),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_36),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_181),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_158),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_40),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_129),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_18),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_139),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_68),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_95),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_61),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_18),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_76),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_87),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_69),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_187),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_92),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_51),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_110),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_131),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_26),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_146),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_188),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_67),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_150),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_126),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_24),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_75),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_14),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_62),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_142),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_21),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_169),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_41),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_103),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_102),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_182),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_57),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_55),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_62),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_44),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_23),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_60),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_116),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_3),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_115),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_114),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_20),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_45),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_70),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_5),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_71),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_172),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_7),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_46),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_52),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_128),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_177),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_27),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_376),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_297),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_199),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_325),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_288),
.B(n_0),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_325),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_215),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_194),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_345),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_345),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_232),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_191),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_191),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_212),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_201),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_201),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_223),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_206),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_248),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_259),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_223),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_206),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_252),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_346),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_210),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_210),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_195),
.B(n_203),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_219),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_272),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_198),
.B(n_2),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_254),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_275),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_323),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_358),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_255),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_219),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_196),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_215),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_249),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_249),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_371),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_215),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_192),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_195),
.B(n_3),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_371),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_198),
.B(n_4),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_207),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_262),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_262),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_214),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_265),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_217),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_227),
.B(n_5),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_374),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_310),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_203),
.B(n_8),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_218),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_220),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_296),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_310),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_296),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_230),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_231),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_371),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_227),
.B(n_10),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_313),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_215),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_313),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_317),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_310),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_233),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_317),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_236),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_321),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_321),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_205),
.B(n_10),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_289),
.B(n_11),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_333),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_333),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_336),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_243),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_336),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_237),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_205),
.B(n_221),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_239),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_221),
.B(n_11),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_193),
.B(n_12),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_222),
.B(n_13),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_215),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_348),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_240),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_348),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_355),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_242),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_355),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_278),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_362),
.B(n_13),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_278),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_278),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_362),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_245),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_385),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_429),
.A2(n_225),
.B(n_222),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_390),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_455),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_455),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_455),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_395),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_413),
.B(n_193),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_404),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_405),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_414),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_450),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_417),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_460),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_485),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_460),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_468),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_427),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_473),
.A2(n_234),
.B(n_225),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_382),
.B(n_224),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_427),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_409),
.B(n_209),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_408),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_384),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_386),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_234),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_453),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_418),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_408),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_470),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_478),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_474),
.B(n_200),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_419),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_383),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_478),
.Y(n_540)
);

AND2x2_ASAP7_75t_SL g541 ( 
.A(n_388),
.B(n_200),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_409),
.A2(n_401),
.B1(n_400),
.B2(n_485),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_398),
.B(n_407),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_410),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_411),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_424),
.B(n_289),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_453),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_422),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_435),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_476),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_425),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_416),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_437),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_447),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_443),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_454),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_444),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_416),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_400),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_448),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_459),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_420),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_458),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_428),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_500),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_526),
.A2(n_484),
.B1(n_396),
.B2(n_403),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_502),
.B(n_401),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_493),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_530),
.A2(n_432),
.B1(n_481),
.B2(n_486),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_541),
.B(n_486),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_541),
.B(n_428),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_518),
.B(n_391),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_528),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_493),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_516),
.B(n_432),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_527),
.B(n_533),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_500),
.B(n_412),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_481),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_555),
.B(n_420),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_543),
.B(n_397),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_537),
.A2(n_471),
.B1(n_520),
.B2(n_490),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_549),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_550),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_507),
.B(n_510),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_510),
.B(n_488),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_558),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_537),
.A2(n_520),
.B1(n_490),
.B2(n_463),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_559),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_489),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_558),
.B(n_488),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_574),
.B(n_562),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_568),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_574),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_567),
.B(n_536),
.Y(n_608)
);

INVx4_ASAP7_75t_SL g609 ( 
.A(n_537),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_495),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_537),
.B(n_472),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_574),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_537),
.A2(n_475),
.B1(n_441),
.B2(n_431),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_537),
.B(n_399),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_537),
.B(n_402),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_497),
.B(n_434),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_498),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_571),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_499),
.Y(n_619)
);

BUFx4f_ASAP7_75t_L g620 ( 
.A(n_490),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_490),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_567),
.B(n_518),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_544),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_544),
.B(n_406),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_498),
.Y(n_625)
);

AND2x6_ASAP7_75t_SL g626 ( 
.A(n_547),
.B(n_365),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_545),
.B(n_466),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_542),
.B(n_244),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_529),
.Y(n_629)
);

CKINVDCx11_ASAP7_75t_R g630 ( 
.A(n_566),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_545),
.B(n_467),
.Y(n_631)
);

AND2x2_ASAP7_75t_SL g632 ( 
.A(n_520),
.B(n_241),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_235),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_543),
.B(n_244),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_536),
.B(n_445),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_522),
.A2(n_438),
.B1(n_451),
.B2(n_415),
.Y(n_636)
);

AND2x4_ASAP7_75t_SL g637 ( 
.A(n_513),
.B(n_440),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_543),
.B(n_452),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_520),
.A2(n_464),
.B1(n_469),
.B2(n_465),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_505),
.B(n_371),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_501),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_546),
.B(n_477),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_491),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_491),
.Y(n_646)
);

BUFx4f_ASAP7_75t_L g647 ( 
.A(n_546),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_506),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_SL g649 ( 
.A1(n_552),
.A2(n_332),
.B1(n_350),
.B2(n_295),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_547),
.B(n_440),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_SL g651 ( 
.A(n_509),
.B(n_241),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_547),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_552),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_512),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_570),
.A2(n_439),
.B1(n_387),
.B2(n_392),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_532),
.B(n_479),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_556),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_556),
.B(n_563),
.Y(n_659)
);

AO22x2_ASAP7_75t_L g660 ( 
.A1(n_547),
.A2(n_389),
.B1(n_392),
.B2(n_387),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_539),
.Y(n_661)
);

OAI221xp5_ASAP7_75t_L g662 ( 
.A1(n_563),
.A2(n_365),
.B1(n_378),
.B2(n_257),
.C(n_373),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_538),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_565),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_565),
.B(n_247),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_517),
.B(n_480),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_560),
.B(n_247),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_569),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_560),
.B(n_260),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_521),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_534),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_492),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_501),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_540),
.B(n_482),
.Y(n_675)
);

AND3x2_ASAP7_75t_L g676 ( 
.A(n_572),
.B(n_378),
.C(n_257),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_560),
.B(n_260),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_572),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_551),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_561),
.B(n_487),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_561),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_494),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_494),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_561),
.B(n_264),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_501),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_515),
.B(n_264),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_515),
.B(n_204),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_523),
.B(n_202),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_523),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_524),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_494),
.B(n_270),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_501),
.B(n_270),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_501),
.B(n_279),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_524),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_496),
.B(n_279),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_524),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_504),
.B(n_389),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_524),
.A2(n_269),
.B1(n_246),
.B2(n_381),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_504),
.B(n_446),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_548),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_503),
.B(n_280),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_496),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_496),
.A2(n_347),
.B1(n_309),
.B2(n_280),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_511),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_511),
.B(n_315),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_525),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_525),
.B(n_446),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_553),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_553),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_578),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_591),
.B(n_300),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_598),
.A2(n_357),
.B(n_557),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_687),
.B(n_304),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_578),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_668),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_653),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_575),
.B(n_305),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_575),
.B(n_305),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_580),
.B(n_251),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_623),
.B(n_308),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_587),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_581),
.B(n_253),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_681),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_394),
.B1(n_457),
.B2(n_347),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_457),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_577),
.B(n_394),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_623),
.B(n_308),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_585),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_632),
.A2(n_665),
.B1(n_639),
.B2(n_576),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_603),
.A2(n_554),
.B(n_553),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_681),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_594),
.B(n_263),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_585),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_589),
.B(n_639),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_668),
.B(n_326),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_592),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_670),
.Y(n_737)
);

AOI22x1_ASAP7_75t_L g738 ( 
.A1(n_690),
.A2(n_335),
.B1(n_379),
.B2(n_326),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_589),
.B(n_331),
.Y(n_739)
);

OAI221xp5_ASAP7_75t_L g740 ( 
.A1(n_628),
.A2(n_271),
.B1(n_291),
.B2(n_320),
.C(n_377),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_671),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_SL g742 ( 
.A(n_602),
.B(n_439),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_665),
.A2(n_341),
.B1(n_331),
.B2(n_352),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_610),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_610),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_576),
.A2(n_613),
.B1(n_647),
.B2(n_643),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_657),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_581),
.B(n_268),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_588),
.B(n_335),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_652),
.A2(n_302),
.B1(n_285),
.B2(n_329),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_665),
.A2(n_349),
.B1(n_352),
.B2(n_379),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_661),
.B(n_274),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_647),
.B(n_343),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_666),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_659),
.B(n_343),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_659),
.B(n_349),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_635),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_620),
.B(n_643),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_584),
.B(n_368),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_680),
.B(n_290),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_622),
.B(n_298),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_582),
.B(n_301),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_625),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_680),
.B(n_311),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_584),
.B(n_224),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_665),
.A2(n_316),
.B1(n_213),
.B2(n_287),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_625),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_584),
.B(n_612),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_680),
.B(n_314),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_591),
.B(n_322),
.Y(n_771)
);

BUFx5_ASAP7_75t_L g772 ( 
.A(n_665),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_628),
.A2(n_316),
.B1(n_258),
.B2(n_380),
.Y(n_773)
);

NAND2x1_ASAP7_75t_L g774 ( 
.A(n_601),
.B(n_548),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_591),
.B(n_213),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_666),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_648),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_654),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_703),
.A2(n_287),
.B1(n_261),
.B2(n_229),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_658),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_619),
.B(n_663),
.C(n_595),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_638),
.B(n_327),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_584),
.B(n_204),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_655),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_664),
.B(n_330),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_666),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_673),
.B(n_678),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_583),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_642),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_586),
.B(n_339),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_600),
.B(n_261),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_612),
.B(n_342),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_597),
.B(n_351),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_596),
.B(n_353),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_586),
.B(n_359),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_633),
.A2(n_294),
.B1(n_216),
.B2(n_375),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_608),
.B(n_226),
.Y(n_797)
);

AND2x2_ASAP7_75t_SL g798 ( 
.A(n_633),
.B(n_226),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_629),
.B(n_360),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_707),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_703),
.A2(n_229),
.B1(n_273),
.B2(n_303),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_634),
.B(n_361),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_634),
.B(n_364),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_600),
.B(n_273),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_688),
.B(n_367),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_606),
.B(n_372),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_611),
.B(n_604),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_612),
.B(n_303),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_593),
.A2(n_366),
.B1(n_356),
.B2(n_328),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_645),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_636),
.A2(n_366),
.B1(n_369),
.B2(n_197),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_612),
.B(n_235),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_653),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_689),
.B(n_208),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_651),
.B(n_650),
.C(n_675),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_627),
.B(n_211),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_631),
.B(n_228),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_644),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_646),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_624),
.A2(n_554),
.B(n_557),
.C(n_20),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_614),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_605),
.B(n_618),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_651),
.A2(n_557),
.B(n_554),
.C(n_306),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_615),
.Y(n_825)
);

BUFx5_ASAP7_75t_L g826 ( 
.A(n_686),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_694),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_593),
.B(n_235),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_605),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_621),
.A2(n_686),
.B1(n_599),
.B2(n_662),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_599),
.B(n_235),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_608),
.B(n_14),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_696),
.Y(n_833)
);

BUFx6f_ASAP7_75t_SL g834 ( 
.A(n_661),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_618),
.B(n_699),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_SL g836 ( 
.A(n_670),
.B(n_238),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_621),
.B(n_16),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_704),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_608),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_601),
.B(n_235),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_679),
.B(n_250),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_672),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_621),
.B(n_21),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_601),
.B(n_235),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_607),
.B(n_235),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_607),
.B(n_235),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_590),
.B(n_23),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_682),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_667),
.A2(n_328),
.B1(n_356),
.B2(n_548),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_741),
.B(n_656),
.Y(n_850)
);

OAI321xp33_ASAP7_75t_L g851 ( 
.A1(n_729),
.A2(n_677),
.A3(n_669),
.B1(n_667),
.B2(n_684),
.C(n_698),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_778),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_734),
.A2(n_640),
.B(n_669),
.C(n_684),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_819),
.B(n_677),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_723),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_780),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_731),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_739),
.B(n_579),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_788),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_747),
.B(n_637),
.Y(n_860)
);

AOI21x1_ASAP7_75t_L g861 ( 
.A1(n_831),
.A2(n_706),
.B(n_708),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_715),
.B(n_609),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_736),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_777),
.B(n_637),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_823),
.B(n_609),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_784),
.B(n_697),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_730),
.A2(n_709),
.B(n_682),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_746),
.A2(n_649),
.B(n_692),
.C(n_701),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_719),
.B(n_749),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_729),
.A2(n_660),
.B1(n_697),
.B2(n_705),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_735),
.A2(n_701),
.B(n_693),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_719),
.B(n_626),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_829),
.B(n_609),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_837),
.A2(n_709),
.B(n_702),
.Y(n_874)
);

BUFx4f_ASAP7_75t_L g875 ( 
.A(n_755),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_798),
.A2(n_697),
.B1(n_653),
.B2(n_660),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_794),
.B(n_722),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_787),
.A2(n_702),
.B(n_683),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_831),
.A2(n_700),
.B(n_685),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_758),
.B(n_660),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_751),
.A2(n_700),
.B(n_27),
.C(n_30),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_722),
.B(n_676),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_837),
.A2(n_695),
.B(n_691),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_748),
.B(n_691),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_710),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_713),
.B(n_691),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_790),
.B(n_630),
.C(n_641),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_843),
.A2(n_319),
.B(n_256),
.C(n_266),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_807),
.B(n_691),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_751),
.A2(n_795),
.B(n_790),
.C(n_740),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_716),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_795),
.A2(n_25),
.B(n_31),
.C(n_33),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_835),
.B(n_674),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_807),
.B(n_695),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_756),
.A2(n_25),
.B(n_31),
.C(n_33),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_843),
.A2(n_844),
.B(n_840),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_714),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_716),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_737),
.Y(n_899)
);

AO21x1_ASAP7_75t_L g900 ( 
.A1(n_828),
.A2(n_695),
.B(n_328),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_789),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_725),
.B(n_630),
.C(n_318),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_841),
.A2(n_324),
.B(n_276),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_716),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_728),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_840),
.A2(n_344),
.B(n_277),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_844),
.A2(n_267),
.B(n_281),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_SL g908 ( 
.A1(n_757),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_733),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_845),
.A2(n_334),
.B(n_283),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_798),
.A2(n_337),
.B1(n_284),
.B2(n_286),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_809),
.A2(n_282),
.B1(n_292),
.B2(n_293),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_845),
.A2(n_354),
.B(n_307),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_809),
.B(n_299),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_782),
.A2(n_34),
.B(n_38),
.C(n_39),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_SL g916 ( 
.A(n_742),
.B(n_312),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_846),
.A2(n_338),
.B(n_340),
.Y(n_917)
);

OAI321xp33_ASAP7_75t_L g918 ( 
.A1(n_724),
.A2(n_328),
.A3(n_356),
.B1(n_503),
.B2(n_508),
.C(n_514),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_846),
.A2(n_328),
.B(n_356),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_762),
.B(n_39),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_822),
.B(n_825),
.Y(n_921)
);

AO32x1_ASAP7_75t_L g922 ( 
.A1(n_744),
.A2(n_548),
.A3(n_535),
.B1(n_531),
.B2(n_514),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_711),
.B(n_535),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_755),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_716),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_745),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_750),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_743),
.A2(n_535),
.B(n_531),
.C(n_514),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_764),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_711),
.B(n_531),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_793),
.A2(n_46),
.B(n_47),
.C(n_54),
.Y(n_931)
);

NOR2xp67_ASAP7_75t_L g932 ( 
.A(n_776),
.B(n_121),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_SL g933 ( 
.A(n_753),
.B(n_47),
.C(n_54),
.Y(n_933)
);

AND2x2_ASAP7_75t_SL g934 ( 
.A(n_724),
.B(n_55),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_768),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_711),
.B(n_514),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_743),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_783),
.A2(n_514),
.B(n_508),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_814),
.Y(n_939)
);

OAI321xp33_ASAP7_75t_L g940 ( 
.A1(n_752),
.A2(n_503),
.A3(n_508),
.B1(n_68),
.B2(n_69),
.C(n_66),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_814),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_726),
.B(n_63),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_711),
.B(n_508),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_755),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_813),
.A2(n_508),
.B(n_503),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_816),
.B(n_66),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_752),
.A2(n_77),
.B1(n_89),
.B2(n_90),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_839),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_830),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_814),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_R g951 ( 
.A(n_834),
.B(n_111),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_791),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_834),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_838),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_817),
.A2(n_132),
.B(n_135),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_818),
.A2(n_148),
.B(n_152),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_827),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_806),
.B(n_157),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_833),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_800),
.B(n_174),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_786),
.B(n_178),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_814),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_L g963 ( 
.A(n_836),
.B(n_773),
.C(n_781),
.Y(n_963)
);

BUFx4f_ASAP7_75t_L g964 ( 
.A(n_804),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_830),
.A2(n_179),
.B1(n_186),
.B2(n_190),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_774),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_754),
.A2(n_712),
.B(n_815),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_791),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_797),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_804),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_754),
.A2(n_727),
.B(n_720),
.C(n_718),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_805),
.B(n_775),
.Y(n_972)
);

BUFx8_ASAP7_75t_L g973 ( 
.A(n_832),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_L g974 ( 
.A1(n_771),
.A2(n_785),
.B(n_799),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_810),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_L g976 ( 
.A(n_732),
.B(n_763),
.C(n_721),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_820),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_775),
.B(n_717),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_761),
.B(n_770),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_769),
.A2(n_842),
.B(n_848),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_802),
.B(n_803),
.C(n_811),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_765),
.B(n_811),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_801),
.A2(n_767),
.B1(n_779),
.B2(n_738),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_772),
.B(n_826),
.Y(n_985)
);

AOI21xp33_ASAP7_75t_L g986 ( 
.A1(n_767),
.A2(n_801),
.B(n_779),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_824),
.A2(n_821),
.B(n_808),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_796),
.A2(n_797),
.B1(n_847),
.B2(n_849),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_808),
.A2(n_766),
.B(n_792),
.Y(n_989)
);

AOI31xp33_ASAP7_75t_L g990 ( 
.A1(n_849),
.A2(n_753),
.A3(n_760),
.B(n_797),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_772),
.A2(n_729),
.B1(n_809),
.B2(n_734),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_826),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_772),
.A2(n_576),
.B(n_739),
.C(n_746),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_826),
.B(n_734),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_826),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_741),
.B(n_616),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_831),
.A2(n_828),
.B(n_759),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_996),
.B(n_850),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_867),
.A2(n_879),
.B(n_997),
.Y(n_999)
);

OAI22x1_ASAP7_75t_L g1000 ( 
.A1(n_876),
.A2(n_946),
.B1(n_872),
.B2(n_934),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_899),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_869),
.A2(n_877),
.B(n_987),
.C(n_896),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_945),
.A2(n_861),
.B(n_938),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_852),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_875),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_985),
.A2(n_981),
.B(n_874),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_863),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_994),
.A2(n_989),
.B(n_884),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_856),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_890),
.A2(n_993),
.B(n_982),
.C(n_983),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_859),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_921),
.B(n_991),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_942),
.B(n_866),
.Y(n_1013)
);

OAI22x1_ASAP7_75t_L g1014 ( 
.A1(n_969),
.A2(n_963),
.B1(n_880),
.B2(n_968),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_860),
.B(n_864),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_991),
.B(n_854),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_974),
.A2(n_868),
.B(n_851),
.C(n_853),
.Y(n_1017)
);

OAI22x1_ASAP7_75t_L g1018 ( 
.A1(n_920),
.A2(n_858),
.B1(n_958),
.B2(n_887),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_952),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_916),
.B(n_964),
.Y(n_1020)
);

AO31x2_ASAP7_75t_L g1021 ( 
.A1(n_900),
.A2(n_971),
.A3(n_870),
.B(n_889),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_870),
.A2(n_894),
.A3(n_889),
.B(n_949),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_976),
.A2(n_988),
.B1(n_972),
.B2(n_984),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_875),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_954),
.Y(n_1025)
);

OAI22x1_ASAP7_75t_L g1026 ( 
.A1(n_902),
.A2(n_882),
.B1(n_957),
.B2(n_959),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_964),
.B(n_970),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_980),
.B(n_885),
.Y(n_1028)
);

INVx8_ASAP7_75t_L g1029 ( 
.A(n_970),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_979),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_924),
.B(n_944),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_897),
.B(n_905),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_909),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_948),
.Y(n_1034)
);

OA21x2_ASAP7_75t_L g1035 ( 
.A1(n_987),
.A2(n_894),
.B(n_878),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_953),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_953),
.B(n_988),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_926),
.B(n_927),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_919),
.A2(n_995),
.B(n_992),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_929),
.B(n_935),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_855),
.B(n_857),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_975),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_901),
.B(n_978),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_965),
.A2(n_928),
.A3(n_886),
.B(n_984),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_955),
.A2(n_956),
.B(n_930),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_871),
.A2(n_906),
.B(n_888),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_923),
.A2(n_936),
.B(n_930),
.Y(n_1047)
);

NOR2xp67_ASAP7_75t_L g1048 ( 
.A(n_961),
.B(n_960),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_970),
.B(n_865),
.Y(n_1049)
);

AND2x2_ASAP7_75t_SL g1050 ( 
.A(n_914),
.B(n_918),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_906),
.A2(n_940),
.B(n_892),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_977),
.B(n_986),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_937),
.B(n_951),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_891),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_986),
.B(n_939),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_937),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_990),
.B(n_893),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_914),
.A2(n_947),
.A3(n_912),
.B(n_936),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_898),
.B(n_939),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_881),
.A2(n_931),
.B(n_915),
.C(n_895),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_898),
.B(n_904),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_923),
.A2(n_943),
.B(n_904),
.Y(n_1062)
);

AO31x2_ASAP7_75t_L g1063 ( 
.A1(n_947),
.A2(n_912),
.A3(n_943),
.B(n_922),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_862),
.A2(n_903),
.B(n_873),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_908),
.Y(n_1065)
);

CKINVDCx11_ASAP7_75t_R g1066 ( 
.A(n_891),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_SL g1067 ( 
.A1(n_891),
.A2(n_950),
.B(n_925),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_911),
.B(n_932),
.Y(n_1068)
);

OAI22x1_ASAP7_75t_L g1069 ( 
.A1(n_973),
.A2(n_933),
.B1(n_922),
.B2(n_950),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_922),
.A2(n_941),
.B(n_962),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_925),
.A2(n_941),
.B(n_962),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_907),
.A2(n_910),
.B(n_913),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_925),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_917),
.A2(n_966),
.B(n_950),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_941),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_962),
.A2(n_966),
.B(n_973),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_966),
.A2(n_867),
.B(n_879),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_852),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_SL g1079 ( 
.A1(n_993),
.A2(n_890),
.B(n_949),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_869),
.B(n_734),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_993),
.B(n_869),
.C(n_946),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_875),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_852),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_996),
.B(n_616),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_869),
.A2(n_729),
.B1(n_934),
.B2(n_734),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_869),
.B(n_734),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_875),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_875),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_852),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_872),
.B(n_385),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_890),
.A2(n_993),
.B(n_869),
.C(n_946),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_L g1092 ( 
.A1(n_869),
.A2(n_877),
.B(n_604),
.C(n_987),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_869),
.B(n_734),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_869),
.B(n_734),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_869),
.B(n_734),
.Y(n_1095)
);

AO21x2_ASAP7_75t_L g1096 ( 
.A1(n_874),
.A2(n_987),
.B(n_883),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_867),
.A2(n_874),
.B(n_896),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_934),
.B(n_798),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_896),
.A2(n_843),
.B(n_837),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_991),
.A2(n_900),
.A3(n_994),
.B(n_853),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_924),
.B(n_944),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_869),
.B(n_734),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_869),
.B(n_734),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_890),
.A2(n_993),
.B(n_869),
.C(n_946),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_852),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_896),
.A2(n_843),
.B(n_837),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_869),
.B(n_734),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_869),
.B(n_734),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_867),
.A2(n_879),
.B(n_997),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_875),
.Y(n_1110)
);

BUFx8_ASAP7_75t_L g1111 ( 
.A(n_996),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_869),
.B(n_734),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_869),
.B(n_734),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_875),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_890),
.A2(n_993),
.B(n_869),
.C(n_946),
.Y(n_1115)
);

AO221x2_ASAP7_75t_L g1116 ( 
.A1(n_937),
.A2(n_576),
.B1(n_746),
.B2(n_870),
.C(n_751),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_869),
.A2(n_877),
.B(n_967),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_852),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_890),
.A2(n_993),
.B(n_869),
.C(n_946),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_869),
.A2(n_526),
.B(n_549),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_867),
.A2(n_879),
.B(n_997),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_890),
.A2(n_993),
.B(n_934),
.Y(n_1122)
);

NOR2x1_ASAP7_75t_L g1123 ( 
.A(n_887),
.B(n_600),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_852),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_869),
.A2(n_877),
.B(n_967),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_867),
.A2(n_879),
.B(n_997),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_896),
.A2(n_843),
.B(n_837),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_890),
.A2(n_993),
.B(n_869),
.C(n_946),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_875),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_1066),
.Y(n_1130)
);

CKINVDCx11_ASAP7_75t_R g1131 ( 
.A(n_1001),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1007),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1005),
.B(n_1110),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1111),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1055),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1120),
.B(n_1053),
.C(n_1090),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1111),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1005),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1084),
.B(n_1028),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1004),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1055),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1116),
.A2(n_1098),
.B1(n_1085),
.B2(n_1000),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1054),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1012),
.Y(n_1144)
);

INVxp67_ASAP7_75t_SL g1145 ( 
.A(n_1012),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1019),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1081),
.A2(n_1104),
.B(n_1091),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1028),
.B(n_1080),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1115),
.A2(n_1128),
.B(n_1119),
.C(n_1010),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_SL g1150 ( 
.A(n_1110),
.B(n_1114),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1114),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1021),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1009),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1080),
.B(n_1086),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_1029),
.B(n_1076),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1086),
.B(n_1093),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1054),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1011),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1082),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1098),
.B(n_1015),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1025),
.Y(n_1162)
);

O2A1O1Ixp5_ASAP7_75t_L g1163 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.C(n_1122),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_998),
.B(n_1013),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1093),
.B(n_1094),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1060),
.A2(n_1079),
.B(n_1122),
.C(n_1017),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1078),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1095),
.B(n_1102),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1002),
.A2(n_1085),
.B(n_1051),
.C(n_1023),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1021),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1116),
.B(n_1056),
.C(n_1051),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1083),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1102),
.A2(n_1113),
.B1(n_1107),
.B2(n_1108),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1089),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1105),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1037),
.B(n_1118),
.Y(n_1177)
);

AO21x1_ASAP7_75t_L g1178 ( 
.A1(n_1016),
.A2(n_1046),
.B(n_1107),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1031),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_SL g1180 ( 
.A1(n_1046),
.A2(n_1117),
.B(n_1125),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1103),
.B(n_1108),
.Y(n_1181)
);

NOR4xp25_ASAP7_75t_L g1182 ( 
.A(n_1065),
.B(n_1103),
.C(n_1113),
.D(n_1112),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1112),
.B(n_1030),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1048),
.B(n_1092),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1041),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1032),
.A2(n_1040),
.B1(n_1038),
.B2(n_1034),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1032),
.A2(n_1040),
.B1(n_1038),
.B2(n_1123),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_1020),
.B1(n_1068),
.B2(n_1018),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1124),
.B(n_1033),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1021),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1031),
.B(n_1101),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1050),
.A2(n_1096),
.B1(n_1042),
.B2(n_1022),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1101),
.B(n_1129),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1024),
.B(n_1129),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1024),
.B(n_1087),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1088),
.B(n_1027),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1100),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1027),
.B(n_1029),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1036),
.B(n_1049),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1059),
.B(n_1061),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1036),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1026),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1029),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1073),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1069),
.B(n_1074),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1049),
.B(n_1075),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1096),
.B(n_1043),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1014),
.Y(n_1208)
);

OR2x2_ASAP7_75t_SL g1209 ( 
.A(n_1035),
.B(n_1052),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1022),
.B(n_1052),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_SL g1211 ( 
.A(n_1064),
.B(n_1008),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1062),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1047),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1077),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1074),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_999),
.A2(n_1126),
.B(n_1121),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1022),
.B(n_1058),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1071),
.B(n_1100),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1058),
.B(n_1044),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1058),
.B(n_1067),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1039),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1070),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1072),
.B(n_1044),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1044),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1097),
.A2(n_1072),
.B1(n_1045),
.B2(n_1006),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1063),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1063),
.B(n_1109),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1003),
.B(n_1084),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1066),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1004),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1004),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1005),
.B(n_1110),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1055),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1066),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1084),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1001),
.Y(n_1236)
);

OR2x6_ASAP7_75t_SL g1237 ( 
.A(n_998),
.B(n_385),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1001),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_998),
.B(n_1084),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1120),
.B(n_934),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1005),
.B(n_1110),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1066),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1084),
.B(n_996),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_1084),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1005),
.B(n_594),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_869),
.B1(n_1127),
.B2(n_1106),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1081),
.A2(n_890),
.B(n_1104),
.C(n_1091),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1001),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1005),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1099),
.A2(n_869),
.B1(n_1127),
.B2(n_1106),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1084),
.B(n_996),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1066),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1084),
.B(n_996),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1005),
.B(n_1110),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1120),
.B(n_934),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1111),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1120),
.B(n_934),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1004),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1084),
.B(n_996),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1066),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1084),
.B(n_996),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1084),
.B(n_996),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1066),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1084),
.B(n_996),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1084),
.B(n_996),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1005),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1029),
.B(n_755),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_998),
.B(n_1084),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1001),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1116),
.A2(n_934),
.B1(n_724),
.B2(n_1098),
.Y(n_1275)
);

OAI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1120),
.A2(n_526),
.B(n_869),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1111),
.Y(n_1277)
);

O2A1O1Ixp5_ASAP7_75t_L g1278 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.C(n_1081),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1066),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1106),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1203),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1248),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1139),
.B(n_1148),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1209),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1143),
.Y(n_1286)
);

NOR2x1_ASAP7_75t_SL g1287 ( 
.A(n_1187),
.B(n_1184),
.Y(n_1287)
);

CKINVDCx11_ASAP7_75t_R g1288 ( 
.A(n_1131),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1144),
.Y(n_1289)
);

CKINVDCx14_ASAP7_75t_R g1290 ( 
.A(n_1131),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1218),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_1229),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1177),
.B(n_1142),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1145),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1189),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_1156),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1218),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1145),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1215),
.B(n_1228),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1156),
.B(n_1147),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1135),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1135),
.Y(n_1302)
);

AO21x2_ASAP7_75t_L g1303 ( 
.A1(n_1180),
.A2(n_1220),
.B(n_1205),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1275),
.A2(n_1261),
.B1(n_1240),
.B2(n_1259),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1201),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1199),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1156),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1275),
.A2(n_1240),
.B1(n_1261),
.B2(n_1259),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1247),
.A2(n_1149),
.B1(n_1246),
.B2(n_1250),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1141),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1214),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1214),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1141),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1233),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1272),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1205),
.B(n_1184),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1136),
.A2(n_1172),
.B1(n_1188),
.B2(n_1235),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1161),
.A2(n_1186),
.B1(n_1142),
.B2(n_1276),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1130),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1233),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1192),
.B(n_1219),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1192),
.B(n_1182),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1207),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1207),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1229),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1210),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1152),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1152),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1247),
.A2(n_1167),
.B(n_1278),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1225),
.A2(n_1221),
.B(n_1213),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1243),
.A2(n_1263),
.B1(n_1256),
.B2(n_1265),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1217),
.B(n_1171),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1269),
.A2(n_1202),
.B1(n_1208),
.B2(n_1266),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1223),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1171),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1200),
.B(n_1155),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1146),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1234),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1170),
.A2(n_1281),
.B1(n_1270),
.B2(n_1258),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1251),
.A2(n_1268),
.B1(n_1174),
.B2(n_1244),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1200),
.B(n_1253),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1234),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1190),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1235),
.A2(n_1244),
.B1(n_1239),
.B2(n_1273),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1164),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1254),
.B(n_1255),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1223),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1140),
.B(n_1153),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1224),
.Y(n_1349)
);

CKINVDCx16_ASAP7_75t_R g1350 ( 
.A(n_1242),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1170),
.A2(n_1279),
.B1(n_1165),
.B2(n_1169),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1190),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_SL g1353 ( 
.A(n_1242),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1237),
.A2(n_1181),
.B1(n_1157),
.B2(n_1166),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1183),
.A2(n_1161),
.B1(n_1185),
.B2(n_1154),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1191),
.B(n_1179),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1159),
.B(n_1176),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1224),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1197),
.Y(n_1359)
);

BUFx4_ASAP7_75t_R g1360 ( 
.A(n_1252),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1178),
.A2(n_1211),
.B(n_1197),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1216),
.A2(n_1227),
.B(n_1278),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_1229),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1226),
.A2(n_1168),
.B(n_1262),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1134),
.A2(n_1137),
.B1(n_1277),
.B2(n_1260),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1162),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1173),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1132),
.A2(n_1230),
.B1(n_1175),
.B2(n_1231),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1163),
.B(n_1226),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1216),
.A2(n_1163),
.B(n_1206),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1236),
.B(n_1274),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1206),
.A2(n_1138),
.B(n_1151),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1238),
.B(n_1160),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1138),
.A2(n_1271),
.B1(n_1249),
.B2(n_1151),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1222),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1204),
.A2(n_1193),
.B1(n_1267),
.B2(n_1252),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1143),
.B(n_1133),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1249),
.A2(n_1271),
.B(n_1198),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1212),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1143),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1196),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1194),
.A2(n_1133),
.B(n_1257),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1267),
.A2(n_1280),
.B1(n_1229),
.B2(n_1264),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1264),
.Y(n_1384)
);

BUFx2_ASAP7_75t_R g1385 ( 
.A(n_1158),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1264),
.B(n_1280),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1158),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1272),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1245),
.A2(n_1150),
.B(n_1241),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1195),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1264),
.B(n_1280),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1280),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1195),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1232),
.A2(n_1116),
.B1(n_934),
.B2(n_660),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1232),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1257),
.B(n_1210),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1209),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1240),
.A2(n_1116),
.B1(n_934),
.B2(n_1098),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1144),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1156),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1177),
.B(n_1142),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1144),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1144),
.Y(n_1403)
);

OR2x2_ASAP7_75t_SL g1404 ( 
.A(n_1136),
.B(n_1172),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1209),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1144),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1209),
.Y(n_1407)
);

AO21x1_ASAP7_75t_L g1408 ( 
.A1(n_1147),
.A2(n_1122),
.B(n_1106),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1209),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1209),
.Y(n_1410)
);

CKINVDCx6p67_ASAP7_75t_R g1411 ( 
.A(n_1130),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1143),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1144),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1240),
.A2(n_1116),
.B1(n_934),
.B2(n_1098),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1144),
.Y(n_1415)
);

NAND2x1_ASAP7_75t_L g1416 ( 
.A(n_1213),
.B(n_1180),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1177),
.B(n_1142),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1209),
.Y(n_1418)
);

INVx5_ASAP7_75t_L g1419 ( 
.A(n_1156),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1240),
.A2(n_1053),
.B1(n_1261),
.B2(n_1259),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1144),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1156),
.B(n_1037),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1209),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1144),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1275),
.A2(n_1116),
.B1(n_934),
.B2(n_660),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1144),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1214),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1177),
.B(n_1142),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1144),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1144),
.Y(n_1430)
);

CKINVDCx6p67_ASAP7_75t_R g1431 ( 
.A(n_1130),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1209),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1156),
.B(n_1037),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1336),
.B(n_1341),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1311),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1305),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1295),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1318),
.A2(n_1398),
.B1(n_1414),
.B2(n_1309),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1336),
.B(n_1341),
.Y(n_1440)
);

AOI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1416),
.A2(n_1339),
.B(n_1408),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1366),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1329),
.A2(n_1351),
.B(n_1354),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1346),
.B(n_1369),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1367),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1282),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1425),
.A2(n_1394),
.B1(n_1304),
.B2(n_1308),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1337),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1311),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1348),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1364),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1364),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1348),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1346),
.B(n_1369),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1332),
.B(n_1347),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1282),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1321),
.B(n_1347),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1289),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1294),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1298),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1298),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1382),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1399),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1322),
.B(n_1334),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1334),
.B(n_1293),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1288),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1334),
.B(n_1293),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1399),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1345),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1348),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1311),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1402),
.Y(n_1474)
);

OAI21xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1389),
.A2(n_1392),
.B(n_1372),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1357),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1325),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1402),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1401),
.B(n_1417),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1403),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1403),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1357),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1325),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1357),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1301),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1332),
.B(n_1301),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1302),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1302),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1300),
.B(n_1422),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1310),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1310),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1313),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1428),
.B(n_1291),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1283),
.B(n_1305),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1313),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1284),
.B(n_1355),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1314),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1382),
.Y(n_1498)
);

BUFx12f_ASAP7_75t_L g1499 ( 
.A(n_1384),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1406),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1362),
.A2(n_1370),
.B(n_1330),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1406),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1428),
.B(n_1291),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1413),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1314),
.B(n_1320),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1413),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1320),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1415),
.Y(n_1508)
);

BUFx12f_ASAP7_75t_L g1509 ( 
.A(n_1319),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1317),
.A2(n_1396),
.B1(n_1316),
.B2(n_1350),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1349),
.B(n_1359),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1415),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1300),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1381),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1312),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1381),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1333),
.A2(n_1300),
.B1(n_1432),
.B2(n_1423),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1359),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1421),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1421),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1424),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1424),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1338),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1306),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1422),
.B(n_1433),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1340),
.B(n_1344),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1349),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1422),
.B(n_1433),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1426),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1426),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1429),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1326),
.B(n_1285),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1373),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1312),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1429),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1312),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1427),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1430),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1430),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1371),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1433),
.B(n_1296),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1327),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1316),
.A2(n_1420),
.B(n_1378),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1427),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1316),
.A2(n_1378),
.B(n_1372),
.Y(n_1547)
);

AO21x1_ASAP7_75t_SL g1548 ( 
.A1(n_1287),
.A2(n_1335),
.B(n_1343),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1299),
.B(n_1397),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1327),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1427),
.Y(n_1551)
);

AOI21xp33_ASAP7_75t_L g1552 ( 
.A1(n_1397),
.A2(n_1409),
.B(n_1423),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1328),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1511),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1519),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1450),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1445),
.B(n_1303),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1434),
.B(n_1405),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1445),
.B(n_1303),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1527),
.B(n_1407),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1455),
.B(n_1361),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1439),
.A2(n_1432),
.B1(n_1407),
.B2(n_1409),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1455),
.B(n_1434),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1444),
.A2(n_1331),
.B1(n_1376),
.B2(n_1383),
.C(n_1404),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1440),
.B(n_1466),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1466),
.B(n_1361),
.Y(n_1566)
);

AOI221x1_ASAP7_75t_L g1567 ( 
.A1(n_1552),
.A2(n_1375),
.B1(n_1387),
.B2(n_1410),
.C(n_1418),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1450),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1501),
.Y(n_1569)
);

NOR2xp67_ASAP7_75t_L g1570 ( 
.A(n_1464),
.B(n_1375),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1544),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_1419),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1511),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1544),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1460),
.B(n_1379),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1467),
.B(n_1343),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1550),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1550),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1467),
.B(n_1469),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1456),
.B(n_1352),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1435),
.B(n_1442),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1493),
.B(n_1382),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1503),
.B(n_1358),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1435),
.B(n_1358),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1486),
.B(n_1396),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1514),
.B(n_1382),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1498),
.B(n_1391),
.Y(n_1590)
);

OAI33xp33_ASAP7_75t_L g1591 ( 
.A1(n_1443),
.A2(n_1365),
.A3(n_1356),
.B1(n_1387),
.B2(n_1388),
.B3(n_1404),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1498),
.B(n_1391),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1479),
.B(n_1386),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1548),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1529),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1507),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1442),
.B(n_1368),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1516),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1459),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_L g1600 ( 
.A(n_1547),
.B(n_1374),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1459),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1509),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1530),
.B(n_1489),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1505),
.B(n_1307),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1548),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1461),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1462),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1448),
.A2(n_1390),
.B1(n_1393),
.B2(n_1400),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1501),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1583),
.B(n_1438),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1600),
.B(n_1545),
.C(n_1449),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1565),
.B(n_1520),
.Y(n_1612)
);

XNOR2xp5_ASAP7_75t_L g1613 ( 
.A(n_1602),
.B(n_1525),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1471),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1596),
.B(n_1451),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1564),
.A2(n_1510),
.B1(n_1528),
.B2(n_1518),
.C(n_1496),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1596),
.B(n_1454),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1600),
.B(n_1517),
.C(n_1515),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1565),
.B(n_1538),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1564),
.B(n_1468),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_L g1621 ( 
.A(n_1555),
.B(n_1487),
.C(n_1485),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1562),
.A2(n_1535),
.B1(n_1542),
.B2(n_1484),
.C(n_1482),
.Y(n_1622)
);

AND2x2_ASAP7_75t_SL g1623 ( 
.A(n_1603),
.B(n_1530),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1555),
.B(n_1491),
.C(n_1488),
.Y(n_1624)
);

NAND4xp25_ASAP7_75t_L g1625 ( 
.A(n_1556),
.B(n_1494),
.C(n_1457),
.D(n_1447),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1579),
.B(n_1472),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1563),
.A2(n_1525),
.B1(n_1437),
.B2(n_1290),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1563),
.B(n_1476),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1595),
.B(n_1497),
.C(n_1495),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1446),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1599),
.B(n_1492),
.C(n_1490),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1554),
.B(n_1573),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1591),
.A2(n_1470),
.B1(n_1474),
.B2(n_1478),
.C(n_1480),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1554),
.B(n_1463),
.Y(n_1634)
);

OAI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1561),
.A2(n_1441),
.B(n_1505),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1599),
.B(n_1470),
.C(n_1465),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1579),
.B(n_1530),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1554),
.B(n_1573),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1557),
.A2(n_1489),
.B1(n_1513),
.B2(n_1549),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1579),
.B(n_1447),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1573),
.B(n_1465),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1581),
.B(n_1539),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1597),
.A2(n_1475),
.B1(n_1534),
.B2(n_1481),
.C(n_1508),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1591),
.A2(n_1499),
.B1(n_1468),
.B2(n_1315),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1581),
.B(n_1546),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1584),
.B(n_1546),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1584),
.B(n_1549),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1588),
.B(n_1436),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1588),
.B(n_1436),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1601),
.B(n_1500),
.C(n_1512),
.Y(n_1650)
);

AND2x2_ASAP7_75t_SL g1651 ( 
.A(n_1603),
.B(n_1489),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1567),
.A2(n_1452),
.B(n_1453),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1594),
.A2(n_1353),
.B1(n_1292),
.B2(n_1338),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1597),
.A2(n_1532),
.B1(n_1512),
.B2(n_1508),
.C(n_1531),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1601),
.B(n_1500),
.C(n_1506),
.Y(n_1655)
);

AND2x2_ASAP7_75t_SL g1656 ( 
.A(n_1603),
.B(n_1543),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1575),
.B(n_1480),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1608),
.A2(n_1534),
.B1(n_1521),
.B2(n_1502),
.C(n_1522),
.Y(n_1658)
);

NAND4xp25_ASAP7_75t_L g1659 ( 
.A(n_1556),
.B(n_1457),
.C(n_1477),
.D(n_1483),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1593),
.B(n_1473),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1587),
.B(n_1502),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1560),
.A2(n_1315),
.B1(n_1395),
.B2(n_1513),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1593),
.B(n_1473),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1606),
.B(n_1524),
.C(n_1504),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1586),
.B(n_1504),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1586),
.B(n_1506),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1594),
.A2(n_1441),
.B(n_1360),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1557),
.A2(n_1531),
.B1(n_1521),
.B2(n_1541),
.C(n_1540),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1593),
.B(n_1477),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_SL g1670 ( 
.A(n_1572),
.B(n_1499),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1606),
.B(n_1522),
.C(n_1523),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1571),
.Y(n_1672)
);

NAND4xp25_ASAP7_75t_L g1673 ( 
.A(n_1568),
.B(n_1483),
.C(n_1551),
.D(n_1536),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1558),
.B(n_1533),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_SL g1675 ( 
.A(n_1598),
.B(n_1526),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1590),
.B(n_1592),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1557),
.A2(n_1541),
.B1(n_1540),
.B2(n_1533),
.C(n_1537),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1676),
.B(n_1559),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1672),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1652),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1676),
.B(n_1559),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1652),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1636),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1615),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1610),
.B(n_1674),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1646),
.B(n_1561),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1675),
.B(n_1570),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1619),
.B(n_1561),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1612),
.B(n_1566),
.Y(n_1691)
);

AND2x4_ASAP7_75t_SL g1692 ( 
.A(n_1642),
.B(n_1572),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1677),
.B(n_1607),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1668),
.B(n_1607),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1650),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1655),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1617),
.B(n_1582),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1654),
.B(n_1571),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1664),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1635),
.B(n_1574),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1648),
.B(n_1570),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1665),
.B(n_1574),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1645),
.B(n_1589),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1577),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1671),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1649),
.B(n_1605),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1645),
.B(n_1589),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1634),
.B(n_1577),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1647),
.B(n_1576),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1641),
.B(n_1578),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1618),
.B(n_1578),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1623),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1630),
.B(n_1580),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1647),
.B(n_1660),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1623),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1651),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1656),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1631),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1657),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1661),
.B(n_1633),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1621),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1712),
.B(n_1637),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1718),
.B(n_1685),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1712),
.B(n_1640),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1679),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1693),
.B(n_1614),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1712),
.B(n_1663),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1692),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1718),
.B(n_1411),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1632),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1679),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1711),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1694),
.B(n_1638),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1720),
.A2(n_1620),
.B(n_1611),
.C(n_1616),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1721),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1721),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1694),
.B(n_1628),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1720),
.B(n_1624),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1682),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1715),
.B(n_1626),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1711),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1682),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1685),
.B(n_1629),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1680),
.A2(n_1716),
.B1(n_1682),
.B2(n_1683),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1686),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1695),
.B(n_1558),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1698),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1695),
.B(n_1643),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1696),
.B(n_1585),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1683),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1698),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1696),
.B(n_1585),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1669),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1713),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1708),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1699),
.B(n_1585),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1699),
.B(n_1411),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1705),
.B(n_1604),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1683),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1708),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1680),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1691),
.B(n_1669),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1710),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1710),
.Y(n_1767)
);

NOR2x1_ASAP7_75t_SL g1768 ( 
.A(n_1716),
.B(n_1667),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1697),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1680),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1748),
.B(n_1686),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1735),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1723),
.B(n_1687),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1729),
.B(n_1431),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1753),
.B(n_1700),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1725),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1731),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1768),
.B(n_1692),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1736),
.B(n_1700),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1768),
.B(n_1692),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1764),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1727),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1769),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1760),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1728),
.B(n_1692),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1742),
.B(n_1717),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1760),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1746),
.B(n_1687),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1732),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1741),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1738),
.B(n_1687),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1742),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1764),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1751),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1751),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1727),
.B(n_1678),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1770),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1755),
.B(n_1717),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1762),
.B(n_1759),
.C(n_1744),
.D(n_1738),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1754),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1749),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1770),
.Y(n_1803)
);

INVx1_ASAP7_75t_SL g1804 ( 
.A(n_1744),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1754),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1722),
.B(n_1678),
.Y(n_1806)
);

AOI21xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1749),
.A2(n_1613),
.B(n_1627),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1739),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1722),
.B(n_1678),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1739),
.Y(n_1810)
);

OAI21xp33_ASAP7_75t_L g1811 ( 
.A1(n_1734),
.A2(n_1680),
.B(n_1625),
.Y(n_1811)
);

NAND2x2_ASAP7_75t_L g1812 ( 
.A(n_1726),
.B(n_1431),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1726),
.B(n_1719),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1745),
.A2(n_1644),
.B(n_1717),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1758),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1765),
.B(n_1681),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1743),
.Y(n_1817)
);

NOR2x1_ASAP7_75t_L g1818 ( 
.A(n_1800),
.B(n_1755),
.Y(n_1818)
);

INVx3_ASAP7_75t_SL g1819 ( 
.A(n_1804),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1792),
.B(n_1737),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1792),
.B(n_1750),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1774),
.B(n_1737),
.Y(n_1822)
);

INVx4_ASAP7_75t_L g1823 ( 
.A(n_1773),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1773),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_SL g1825 ( 
.A(n_1787),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1774),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1793),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1793),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1789),
.B(n_1730),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1778),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1775),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1772),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1779),
.B(n_1724),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1778),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1790),
.B(n_1756),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1785),
.B(n_1730),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1779),
.B(n_1724),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1771),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1807),
.B(n_1319),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1783),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1785),
.B(n_1733),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1771),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1783),
.Y(n_1843)
);

NAND3x1_ASAP7_75t_L g1844 ( 
.A(n_1781),
.B(n_1717),
.C(n_1740),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1788),
.B(n_1733),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1781),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1777),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1802),
.B(n_1757),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1787),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1788),
.B(n_1767),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1791),
.B(n_1807),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1811),
.A2(n_1761),
.B1(n_1752),
.B2(n_1743),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1786),
.B(n_1806),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1777),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1791),
.Y(n_1855)
);

INVx4_ASAP7_75t_L g1856 ( 
.A(n_1787),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1852),
.A2(n_1811),
.B1(n_1814),
.B2(n_1776),
.C(n_1780),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1852),
.A2(n_1784),
.B(n_1808),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1842),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1842),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1818),
.A2(n_1752),
.B1(n_1761),
.B2(n_1810),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1828),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1819),
.A2(n_1812),
.B1(n_1717),
.B2(n_1809),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1784),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1839),
.B(n_1509),
.Y(n_1865)
);

AND2x2_ASAP7_75t_SL g1866 ( 
.A(n_1823),
.B(n_1644),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1839),
.B(n_1813),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1828),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1831),
.B(n_1787),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1840),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1826),
.B(n_1843),
.Y(n_1871)
);

OAI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1851),
.A2(n_1812),
.B1(n_1716),
.B2(n_1758),
.Y(n_1872)
);

AOI32xp33_ASAP7_75t_L g1873 ( 
.A1(n_1832),
.A2(n_1799),
.A3(n_1796),
.B1(n_1815),
.B2(n_1795),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1823),
.B(n_1816),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1820),
.A2(n_1812),
.B1(n_1846),
.B2(n_1822),
.Y(n_1875)
);

OAI21xp33_ASAP7_75t_L g1876 ( 
.A1(n_1821),
.A2(n_1796),
.B(n_1795),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1838),
.Y(n_1877)
);

OAI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1848),
.A2(n_1801),
.B1(n_1815),
.B2(n_1805),
.C(n_1794),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1853),
.B(n_1833),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1844),
.A2(n_1809),
.B(n_1806),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1847),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1854),
.Y(n_1882)
);

OAI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1823),
.A2(n_1829),
.B1(n_1824),
.B2(n_1836),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1856),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1824),
.B(n_1816),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1862),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1864),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1870),
.B(n_1827),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1873),
.A2(n_1849),
.B(n_1837),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1868),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1879),
.B(n_1856),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1883),
.B(n_1827),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1871),
.B(n_1841),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1883),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1880),
.B(n_1856),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1865),
.B(n_1825),
.Y(n_1896)
);

NOR2x1_ASAP7_75t_L g1897 ( 
.A(n_1859),
.B(n_1855),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1874),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1869),
.B(n_1825),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1876),
.B(n_1845),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1884),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1860),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1868),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1885),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1857),
.A2(n_1817),
.B1(n_1810),
.B2(n_1794),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1877),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1881),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1875),
.Y(n_1908)
);

AOI31xp33_ASAP7_75t_L g1909 ( 
.A1(n_1894),
.A2(n_1867),
.A3(n_1861),
.B(n_1863),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1890),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1891),
.Y(n_1911)
);

NAND3xp33_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1858),
.C(n_1878),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1892),
.Y(n_1913)
);

NOR2x1_ASAP7_75t_L g1914 ( 
.A(n_1897),
.B(n_1882),
.Y(n_1914)
);

NOR3xp33_ASAP7_75t_L g1915 ( 
.A(n_1887),
.B(n_1872),
.C(n_1834),
.Y(n_1915)
);

NAND4xp25_ASAP7_75t_L g1916 ( 
.A(n_1899),
.B(n_1835),
.C(n_1830),
.D(n_1850),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1898),
.B(n_1866),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1889),
.A2(n_1866),
.B(n_1798),
.Y(n_1918)
);

AOI322xp5_ASAP7_75t_L g1919 ( 
.A1(n_1908),
.A2(n_1803),
.A3(n_1794),
.B1(n_1798),
.B2(n_1817),
.C1(n_1810),
.C2(n_1782),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1905),
.A2(n_1844),
.B1(n_1798),
.B2(n_1803),
.Y(n_1920)
);

OAI322xp33_ASAP7_75t_L g1921 ( 
.A1(n_1890),
.A2(n_1805),
.A3(n_1801),
.B1(n_1803),
.B2(n_1817),
.C1(n_1782),
.C2(n_1747),
.Y(n_1921)
);

AOI21xp33_ASAP7_75t_SL g1922 ( 
.A1(n_1893),
.A2(n_1342),
.B(n_1653),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1891),
.B(n_1786),
.Y(n_1923)
);

NAND2x1_ASAP7_75t_L g1924 ( 
.A(n_1895),
.B(n_1797),
.Y(n_1924)
);

AOI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1900),
.A2(n_1766),
.B1(n_1763),
.B2(n_1622),
.C(n_1797),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1914),
.Y(n_1926)
);

NOR3xp33_ASAP7_75t_L g1927 ( 
.A(n_1912),
.B(n_1903),
.C(n_1888),
.Y(n_1927)
);

NAND3xp33_ASAP7_75t_L g1928 ( 
.A(n_1910),
.B(n_1886),
.C(n_1902),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1911),
.B(n_1904),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1917),
.B(n_1893),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1918),
.B(n_1901),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1909),
.A2(n_1895),
.B(n_1896),
.Y(n_1932)
);

NOR2x1_ASAP7_75t_L g1933 ( 
.A(n_1924),
.B(n_1907),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_SL g1934 ( 
.A(n_1923),
.B(n_1907),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1913),
.Y(n_1935)
);

AND4x1_ASAP7_75t_L g1936 ( 
.A(n_1915),
.B(n_1906),
.C(n_1670),
.D(n_1342),
.Y(n_1936)
);

AND5x1_ASAP7_75t_L g1937 ( 
.A(n_1919),
.B(n_1662),
.C(n_1659),
.D(n_1363),
.E(n_1385),
.Y(n_1937)
);

NOR2x1p5_ASAP7_75t_L g1938 ( 
.A(n_1916),
.B(n_1763),
.Y(n_1938)
);

NOR3xp33_ASAP7_75t_L g1939 ( 
.A(n_1921),
.B(n_1922),
.C(n_1920),
.Y(n_1939)
);

OAI21xp33_ASAP7_75t_L g1940 ( 
.A1(n_1925),
.A2(n_1766),
.B(n_1740),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1921),
.B(n_1389),
.C(n_1689),
.Y(n_1941)
);

NAND2x1_ASAP7_75t_SL g1942 ( 
.A(n_1933),
.B(n_1765),
.Y(n_1942)
);

NAND4xp25_ASAP7_75t_L g1943 ( 
.A(n_1932),
.B(n_1673),
.C(n_1363),
.D(n_1605),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1939),
.A2(n_1689),
.B1(n_1701),
.B2(n_1691),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1934),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1935),
.B(n_1719),
.Y(n_1946)
);

NOR3xp33_ASAP7_75t_L g1947 ( 
.A(n_1931),
.B(n_1689),
.C(n_1412),
.Y(n_1947)
);

NAND4xp25_ASAP7_75t_L g1948 ( 
.A(n_1927),
.B(n_1701),
.C(n_1706),
.D(n_1689),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1926),
.B(n_1702),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1944),
.A2(n_1941),
.B1(n_1930),
.B2(n_1940),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1945),
.B(n_1929),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1948),
.A2(n_1928),
.B1(n_1938),
.B2(n_1937),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1947),
.A2(n_1928),
.B1(n_1936),
.B2(n_1689),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1942),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1949),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1946),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1943),
.A2(n_1658),
.B1(n_1609),
.B2(n_1569),
.Y(n_1957)
);

NAND2xp33_ASAP7_75t_SL g1958 ( 
.A(n_1954),
.B(n_1714),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1951),
.B(n_1697),
.Y(n_1959)
);

AND3x4_ASAP7_75t_L g1960 ( 
.A(n_1952),
.B(n_1701),
.C(n_1706),
.Y(n_1960)
);

NAND3x1_ASAP7_75t_L g1961 ( 
.A(n_1956),
.B(n_1714),
.C(n_1709),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1955),
.B(n_1697),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1950),
.Y(n_1963)
);

XNOR2x1_ASAP7_75t_SL g1964 ( 
.A(n_1953),
.B(n_1714),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1958),
.Y(n_1965)
);

XNOR2xp5_ASAP7_75t_L g1966 ( 
.A(n_1960),
.B(n_1957),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1964),
.Y(n_1967)
);

OAI22x1_ASAP7_75t_L g1968 ( 
.A1(n_1967),
.A2(n_1963),
.B1(n_1959),
.B2(n_1962),
.Y(n_1968)
);

AOI22x1_ASAP7_75t_L g1969 ( 
.A1(n_1968),
.A2(n_1965),
.B1(n_1966),
.B2(n_1961),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1969),
.A2(n_1691),
.B1(n_1681),
.B2(n_1701),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1969),
.A2(n_1681),
.B1(n_1701),
.B2(n_1688),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1970),
.A2(n_1971),
.B(n_1704),
.Y(n_1972)
);

NOR3xp33_ASAP7_75t_L g1973 ( 
.A(n_1970),
.B(n_1412),
.C(n_1286),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1973),
.A2(n_1688),
.B1(n_1703),
.B2(n_1707),
.Y(n_1974)
);

XNOR2x1_ASAP7_75t_L g1975 ( 
.A(n_1972),
.B(n_1377),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1975),
.B(n_1684),
.Y(n_1976)
);

BUFx2_ASAP7_75t_L g1977 ( 
.A(n_1976),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_R g1978 ( 
.A1(n_1977),
.A2(n_1974),
.B1(n_1639),
.B2(n_1706),
.C(n_1709),
.Y(n_1978)
);

AOI211xp5_ASAP7_75t_L g1979 ( 
.A1(n_1978),
.A2(n_1688),
.B(n_1380),
.C(n_1690),
.Y(n_1979)
);


endmodule