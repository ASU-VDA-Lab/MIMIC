module fake_jpeg_8459_n_168 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_6),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx12_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_38),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_39),
.B(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_22),
.B1(n_13),
.B2(n_12),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_20),
.C(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_46),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_30),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_49),
.B1(n_41),
.B2(n_33),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_31),
.B1(n_23),
.B2(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_25),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_31),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_29),
.B1(n_23),
.B2(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_45),
.B1(n_51),
.B2(n_32),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_49),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_55),
.B1(n_57),
.B2(n_49),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_69),
.B1(n_49),
.B2(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_44),
.B1(n_55),
.B2(n_35),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_45),
.B1(n_56),
.B2(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_77),
.B(n_81),
.Y(n_97)
);

BUFx12f_ASAP7_75t_SL g77 ( 
.A(n_70),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_66),
.C(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_72),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_52),
.B(n_48),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_89),
.B(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_48),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_62),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_99),
.C(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_60),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_46),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_35),
.B1(n_13),
.B2(n_15),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_61),
.Y(n_100)
);

OAI322xp33_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_85),
.A3(n_69),
.B1(n_77),
.B2(n_81),
.C1(n_12),
.C2(n_16),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_114),
.C(n_116),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_80),
.B1(n_77),
.B2(n_66),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_101),
.B1(n_97),
.B2(n_99),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_20),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_46),
.C(n_28),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_28),
.C(n_11),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_126),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_0),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_109),
.B(n_107),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_20),
.C(n_18),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_127),
.B(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_125),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_20),
.C(n_18),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_110),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_106),
.C(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_133),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_118),
.B1(n_127),
.B2(n_111),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_117),
.C(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_117),
.C(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_9),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_19),
.C(n_14),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_0),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_133),
.B1(n_19),
.B2(n_14),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_146),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_14),
.A3(n_6),
.B1(n_7),
.B2(n_10),
.C1(n_5),
.C2(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_152),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_5),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_158),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_142),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_148),
.B(n_141),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

AOI21x1_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_5),
.B(n_8),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_164),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_2),
.C(n_3),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);


endmodule