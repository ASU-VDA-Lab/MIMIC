module fake_jpeg_6285_n_331 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_50),
.Y(n_74)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_47),
.Y(n_72)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_53),
.B(n_54),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_57),
.B(n_63),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_17),
.B1(n_15),
.B2(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_83),
.B1(n_27),
.B2(n_25),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_15),
.B1(n_17),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_60),
.B1(n_32),
.B2(n_28),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_16),
.B1(n_15),
.B2(n_17),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_25),
.B1(n_30),
.B2(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_70),
.Y(n_113)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_82),
.Y(n_132)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_91),
.Y(n_131)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_88),
.Y(n_114)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_31),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_18),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_19),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_19),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_36),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_24),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_36),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_36),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_107),
.B1(n_86),
.B2(n_56),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_59),
.A2(n_30),
.B1(n_9),
.B2(n_12),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_59),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_92),
.B1(n_98),
.B2(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_100),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_84),
.B(n_97),
.C(n_89),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_23),
.B(n_9),
.C(n_12),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_10),
.B(n_9),
.C(n_8),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_59),
.B(n_23),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_60),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_139),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_136),
.A2(n_165),
.B1(n_122),
.B2(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_146),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_104),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_148),
.B1(n_154),
.B2(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_64),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_156),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_72),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_147),
.B(n_150),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_84),
.B1(n_86),
.B2(n_90),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_74),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_71),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_71),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_162),
.B(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_64),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_103),
.A2(n_23),
.B(n_67),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_117),
.B(n_115),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_113),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_158),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_88),
.B1(n_28),
.B2(n_32),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_122),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_68),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_168),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_70),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_23),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_125),
.C(n_124),
.Y(n_183)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_123),
.B(n_125),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_173),
.A2(n_174),
.B(n_186),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_177),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_180),
.B(n_203),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_139),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_126),
.B(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_162),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_140),
.A2(n_154),
.B1(n_148),
.B2(n_135),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_193),
.A2(n_198),
.B1(n_175),
.B2(n_142),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_121),
.B1(n_118),
.B2(n_106),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_133),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_201),
.Y(n_212)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_69),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_133),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_130),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_170),
.C(n_137),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_139),
.B(n_10),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_158),
.B(n_157),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_115),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_3),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_142),
.A2(n_109),
.B1(n_117),
.B2(n_130),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_167),
.B1(n_166),
.B2(n_161),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_231),
.B1(n_186),
.B2(n_187),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_228),
.B(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_149),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_222),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_178),
.B(n_188),
.C(n_176),
.Y(n_255)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_156),
.B(n_109),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_234),
.B(n_237),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_196),
.B1(n_177),
.B2(n_175),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_198),
.B1(n_190),
.B2(n_209),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_194),
.C(n_183),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_141),
.B(n_165),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_236),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_193),
.A2(n_111),
.B1(n_108),
.B2(n_159),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_232),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_172),
.Y(n_236)
);

OAI22x1_ASAP7_75t_SL g237 ( 
.A1(n_174),
.A2(n_69),
.B1(n_62),
.B2(n_61),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_111),
.B(n_28),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_202),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_257),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_229),
.B1(n_222),
.B2(n_212),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_251),
.C(n_258),
.Y(n_276)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_252),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_238),
.B(n_228),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_206),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_190),
.B1(n_195),
.B2(n_178),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_253),
.A2(n_211),
.B1(n_218),
.B2(n_213),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_214),
.B(n_233),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_182),
.A3(n_195),
.B1(n_176),
.B2(n_188),
.C1(n_208),
.C2(n_184),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_182),
.C(n_189),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_179),
.B1(n_191),
.B2(n_200),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_231),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_224),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_277),
.C(n_251),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_264),
.B(n_265),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_224),
.B(n_226),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_230),
.B(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_268),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_261),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_275),
.B1(n_247),
.B2(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_246),
.A2(n_248),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_279),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_225),
.C(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.C(n_279),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_240),
.C(n_244),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_290),
.C(n_294),
.Y(n_298)
);

AOI321xp33_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_240),
.A3(n_249),
.B1(n_217),
.B2(n_260),
.C(n_226),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_271),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_260),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_278),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_265),
.B(n_274),
.C(n_263),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_249),
.C(n_239),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_260),
.C(n_254),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_296),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_267),
.C(n_268),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_299),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_232),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_304),
.B(n_291),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_271),
.C(n_269),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_284),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_273),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_217),
.C(n_252),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_294),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_293),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_314),
.B(n_243),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_311),
.B(n_313),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_281),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_298),
.C(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_215),
.C(n_179),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_243),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_308),
.A2(n_191),
.B1(n_8),
.B2(n_197),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_197),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_310),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_320),
.B(n_315),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_323),
.B(n_324),
.Y(n_330)
);

XOR2x1_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_328),
.Y(n_331)
);


endmodule