module fake_netlist_6_3583_n_4405 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4405);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4405;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3813;
wire n_3660;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_700;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_798;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2974;
wire n_2886;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4026;
wire n_4065;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_544;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_835;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_539;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_1986;
wire n_2300;
wire n_699;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_1909;
wire n_2080;
wire n_813;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_606;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_792;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_2714;
wire n_1289;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_1236;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_586;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_3337;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3431;
wire n_3450;
wire n_3253;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_2693;
wire n_1293;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_791;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3348;
wire n_3229;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_738;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_3580;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_947;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_2403;
wire n_1070;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1178;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_716;
wire n_2354;
wire n_2682;
wire n_3103;
wire n_3032;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_683;
wire n_2442;
wire n_1207;
wire n_811;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_1837;
wire n_831;
wire n_2218;
wire n_964;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_2250;
wire n_1951;
wire n_3090;
wire n_4299;
wire n_3724;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1286;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3364;
wire n_3226;
wire n_3323;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_3646;
wire n_2801;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4056;
wire n_4034;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2289;
wire n_2315;
wire n_1733;
wire n_688;
wire n_1077;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4030;
wire n_1129;
wire n_3870;
wire n_4003;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_952;
wire n_725;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_4234;
wire n_4304;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_710;
wire n_1108;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_1601;
wire n_609;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_662;
wire n_3501;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2760;
wire n_1940;
wire n_1979;
wire n_2560;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_1823;
wire n_776;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3439;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_3858;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_3292;
wire n_1271;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_799;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_4369;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3932;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_786;
wire n_706;
wire n_3506;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2787;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_3268;
wire n_2149;
wire n_1754;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_3486;
wire n_1414;
wire n_4086;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_839;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_779;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_709;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4105;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_570;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_756;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_2477;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_629;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g509 ( 
.A(n_255),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_28),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_289),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_493),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_398),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_275),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_360),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_376),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_21),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_127),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_306),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_32),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_273),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_208),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_213),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_298),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_53),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_400),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_424),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_465),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_289),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_104),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_94),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_464),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_432),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_223),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_176),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_102),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_72),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_121),
.Y(n_539)
);

BUFx5_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_110),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_354),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_197),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_119),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_476),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_208),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_358),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_137),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_20),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_447),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_268),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_255),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_204),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_53),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_66),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_237),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_337),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_18),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_138),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_66),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_108),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_343),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_345),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_318),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_470),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_280),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_317),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_501),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_410),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_346),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_386),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_363),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_478),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_78),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_263),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_3),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_497),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_197),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_483),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_77),
.Y(n_580)
);

BUFx5_ASAP7_75t_L g581 ( 
.A(n_431),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_199),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_244),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_140),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_204),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_202),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_185),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_334),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_89),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_131),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_214),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_25),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_389),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_438),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_48),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_49),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_108),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_420),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_147),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_395),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_246),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_347),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_139),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_262),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_222),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_140),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_239),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_158),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_193),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_351),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_192),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_100),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_361),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_428),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_404),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_149),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_403),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_107),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_70),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_250),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_82),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_212),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_216),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_169),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_199),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_149),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_231),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_162),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_183),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_83),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_391),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_128),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_302),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_281),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_418),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_68),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_118),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_407),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_61),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_4),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_109),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_59),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_384),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_189),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_25),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_225),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_301),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_433),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_171),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_183),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_250),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_502),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_85),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_72),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_405),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_132),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_392),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_35),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_40),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_335),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_75),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_121),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_318),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_416),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_181),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_308),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_122),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_17),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_408),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_397),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_257),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_124),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_307),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_417),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_375),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_412),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_322),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_472),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_33),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_174),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_48),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_311),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_215),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_9),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_150),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_31),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_12),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_390),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_5),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_339),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_482),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_65),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_242),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_369),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_381),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_304),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_344),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_122),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_456),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_132),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_460),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_100),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_223),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_4),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_103),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_42),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_363),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_406),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_80),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_260),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_291),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_263),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_336),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_361),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_224),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_22),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_139),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_189),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_207),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_176),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_1),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_155),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_73),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_342),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_180),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_278),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_224),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_196),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_468),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_92),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_254),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_333),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_57),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_459),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_8),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_244),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_328),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_429),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_351),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_146),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_136),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_158),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_365),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_287),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_328),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_168),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_16),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_368),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_181),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_11),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_327),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_28),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_24),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_162),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_481),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_200),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_59),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_173),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_475),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_47),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_37),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_141),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_73),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_164),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_360),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_343),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_415),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_495),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_217),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_50),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_90),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_257),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_299),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_27),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_58),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_437),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_445),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_461),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_430),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_505),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_18),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_494),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_164),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_115),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_321),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_138),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_41),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_54),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_284),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_269),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_36),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_254),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_147),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_249),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_427),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_253),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_38),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_443),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_492),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_266),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_458),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_143),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_409),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_362),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_89),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_42),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_14),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_81),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_330),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_151),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_36),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_195),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_348),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_127),
.Y(n_816)
);

BUFx10_ASAP7_75t_L g817 ( 
.A(n_95),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_50),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_98),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_51),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_348),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_490),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_388),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_785),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_785),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_785),
.Y(n_826)
);

INVxp33_ASAP7_75t_L g827 ( 
.A(n_695),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_689),
.Y(n_828)
);

BUFx5_ASAP7_75t_L g829 ( 
.A(n_522),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_785),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_785),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_511),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_550),
.Y(n_833)
);

BUFx2_ASAP7_75t_SL g834 ( 
.A(n_569),
.Y(n_834)
);

INVx4_ASAP7_75t_R g835 ( 
.A(n_645),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_785),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_785),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_678),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_785),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_785),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_511),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_524),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_511),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_576),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_645),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_511),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_511),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_511),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_562),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_576),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_689),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_562),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_562),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_603),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_562),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_562),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_562),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_662),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_662),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_730),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_532),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_603),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_517),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_662),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_751),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_569),
.B(n_0),
.Y(n_866)
);

INVxp33_ASAP7_75t_L g867 ( 
.A(n_730),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_662),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_662),
.Y(n_869)
);

INVxp33_ASAP7_75t_SL g870 ( 
.A(n_518),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_662),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_519),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_521),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_682),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_682),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_682),
.Y(n_876)
);

CKINVDCx14_ASAP7_75t_R g877 ( 
.A(n_532),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_663),
.B(n_0),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_522),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_528),
.Y(n_880)
);

INVxp33_ASAP7_75t_SL g881 ( 
.A(n_525),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_528),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_529),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_616),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_682),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_529),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_533),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_533),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_571),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_534),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_539),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_514),
.B(n_1),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_514),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_701),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_534),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_545),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_545),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_579),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_530),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_579),
.Y(n_900)
);

INVxp33_ASAP7_75t_SL g901 ( 
.A(n_542),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_543),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_701),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_582),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_582),
.Y(n_905)
);

CKINVDCx14_ASAP7_75t_R g906 ( 
.A(n_532),
.Y(n_906)
);

CKINVDCx16_ASAP7_75t_R g907 ( 
.A(n_784),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_587),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_587),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_659),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_659),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_532),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_530),
.B(n_2),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_671),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_682),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_617),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_745),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_671),
.Y(n_918)
);

INVxp33_ASAP7_75t_L g919 ( 
.A(n_535),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_682),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_690),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_626),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_515),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_571),
.Y(n_924)
);

CKINVDCx14_ASAP7_75t_R g925 ( 
.A(n_556),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_690),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_703),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_703),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_757),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_784),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_757),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_769),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_626),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_769),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_770),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_770),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_782),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_626),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_782),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_515),
.Y(n_940)
);

CKINVDCx14_ASAP7_75t_R g941 ( 
.A(n_556),
.Y(n_941)
);

INVxp33_ASAP7_75t_SL g942 ( 
.A(n_544),
.Y(n_942)
);

INVxp67_ASAP7_75t_SL g943 ( 
.A(n_626),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_520),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_520),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_523),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_523),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_585),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_546),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_585),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_656),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_656),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_626),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_722),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_571),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_722),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_535),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_509),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_788),
.Y(n_959)
);

INVxp33_ASAP7_75t_SL g960 ( 
.A(n_548),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_509),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_510),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_510),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_541),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_541),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_611),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_611),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_621),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_549),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_621),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_643),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_540),
.Y(n_972)
);

INVxp33_ASAP7_75t_SL g973 ( 
.A(n_551),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_858),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_858),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_864),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_864),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_832),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_844),
.A2(n_618),
.B1(n_627),
.B2(n_567),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_834),
.B(n_513),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_832),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_842),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_832),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_933),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_940),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_933),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_953),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_867),
.A2(n_748),
.B1(n_553),
.B2(n_554),
.Y(n_988)
);

CKINVDCx11_ASAP7_75t_R g989 ( 
.A(n_833),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_844),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_959),
.B(n_788),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_829),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_876),
.B(n_595),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_850),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_829),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_922),
.Y(n_996)
);

INVx6_ASAP7_75t_L g997 ( 
.A(n_829),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_885),
.B(n_595),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_953),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_841),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_841),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_843),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_843),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_846),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_846),
.Y(n_1005)
);

INVxp33_ASAP7_75t_SL g1006 ( 
.A(n_842),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_850),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_884),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_847),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_847),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_848),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_889),
.Y(n_1012)
);

INVx5_ASAP7_75t_L g1013 ( 
.A(n_972),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_848),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_854),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_829),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_916),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_915),
.B(n_731),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_972),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_938),
.Y(n_1020)
);

INVx5_ASAP7_75t_L g1021 ( 
.A(n_889),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_849),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_920),
.B(n_731),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_943),
.B(n_573),
.Y(n_1024)
);

AOI22x1_ASAP7_75t_SL g1025 ( 
.A1(n_917),
.A2(n_684),
.B1(n_686),
.B2(n_660),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_849),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_852),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_923),
.Y(n_1028)
);

OAI22x1_ASAP7_75t_SL g1029 ( 
.A1(n_854),
.A2(n_737),
.B1(n_767),
.B2(n_708),
.Y(n_1029)
);

BUFx8_ASAP7_75t_SL g1030 ( 
.A(n_862),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_862),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_852),
.A2(n_820),
.B(n_537),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_853),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_828),
.A2(n_804),
.B1(n_814),
.B2(n_795),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_853),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_894),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_855),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_855),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_856),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_845),
.B(n_823),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_834),
.B(n_512),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_856),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_879),
.B(n_573),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_857),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_924),
.B(n_822),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_857),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_825),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_880),
.B(n_573),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_825),
.Y(n_1050)
);

BUFx8_ASAP7_75t_L g1051 ( 
.A(n_861),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_859),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_829),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_860),
.A2(n_526),
.B1(n_634),
.B2(n_555),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_882),
.B(n_573),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_944),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_863),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_945),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_863),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_868),
.Y(n_1060)
);

CKINVDCx6p67_ASAP7_75t_R g1061 ( 
.A(n_903),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_868),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_869),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_826),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_869),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_871),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_946),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_907),
.Y(n_1068)
);

OAI22x1_ASAP7_75t_R g1069 ( 
.A1(n_872),
.A2(n_559),
.B1(n_561),
.B2(n_552),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_871),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_947),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_872),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_883),
.B(n_573),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_948),
.B(n_704),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_826),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_874),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_874),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_924),
.B(n_516),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_875),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_873),
.Y(n_1080)
);

OA22x2_ASAP7_75t_SL g1081 ( 
.A1(n_838),
.A2(n_537),
.B1(n_538),
.B2(n_536),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_875),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_839),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_824),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_839),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_886),
.B(n_573),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_830),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_831),
.Y(n_1088)
);

BUFx8_ASAP7_75t_SL g1089 ( 
.A(n_873),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_891),
.Y(n_1090)
);

CKINVDCx11_ASAP7_75t_R g1091 ( 
.A(n_930),
.Y(n_1091)
);

NOR2x1_ASAP7_75t_L g1092 ( 
.A(n_955),
.B(n_577),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_955),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_887),
.B(n_619),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_891),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_836),
.Y(n_1096)
);

INVx5_ASAP7_75t_L g1097 ( 
.A(n_923),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1083),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1056),
.B(n_888),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1083),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1085),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_996),
.B(n_1020),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_987),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_L g1104 ( 
.A(n_1092),
.B(n_902),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1085),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1047),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_986),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_986),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_987),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1028),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1047),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_974),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1047),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_974),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_975),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1047),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_975),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_976),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1050),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_976),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1024),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1000),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_996),
.B(n_829),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1050),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1024),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_977),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1050),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1050),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_1026),
.A2(n_837),
.B(n_840),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_977),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1040),
.B(n_870),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1097),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_982),
.B(n_1006),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1024),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_SL g1136 ( 
.A(n_982),
.B(n_750),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1001),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1000),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1064),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1024),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1001),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1064),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1002),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_1036),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1020),
.B(n_829),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1000),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_986),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_986),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1064),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1000),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1064),
.Y(n_1151)
);

BUFx8_ASAP7_75t_L g1152 ( 
.A(n_1015),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1075),
.A2(n_840),
.B(n_890),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_991),
.B(n_895),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1002),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1003),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_991),
.B(n_896),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1003),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_986),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1075),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1097),
.B(n_980),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1027),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1084),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_1026),
.A2(n_898),
.B(n_897),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1075),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1075),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1097),
.B(n_870),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1084),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1084),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1097),
.B(n_900),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1056),
.B(n_904),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1097),
.B(n_905),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1037),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1037),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1038),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1038),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1042),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1027),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1097),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1042),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1089),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_993),
.B(n_829),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1092),
.B(n_881),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1030),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1044),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1046),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_993),
.B(n_998),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_993),
.B(n_866),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_993),
.B(n_908),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_998),
.B(n_909),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1039),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_1032),
.B(n_892),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1084),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1004),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1046),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1039),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1060),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1091),
.Y(n_1199)
);

AND2x2_ASAP7_75t_SL g1200 ( 
.A(n_1032),
.B(n_892),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1012),
.B(n_881),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1084),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_998),
.B(n_1018),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1060),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1074),
.B(n_910),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1087),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1066),
.Y(n_1207)
);

XNOR2xp5_ASAP7_75t_L g1208 ( 
.A(n_1029),
.B(n_851),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1049),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1007),
.Y(n_1210)
);

AND2x6_ASAP7_75t_L g1211 ( 
.A(n_998),
.B(n_643),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_L g1212 ( 
.A(n_1041),
.B(n_902),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1066),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_978),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_978),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1074),
.B(n_911),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_978),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_978),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_981),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_981),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1049),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1007),
.Y(n_1222)
);

AND2x6_ASAP7_75t_L g1223 ( 
.A(n_1018),
.B(n_648),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_981),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1004),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1052),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1052),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1034),
.A2(n_906),
.B1(n_925),
.B2(n_877),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1018),
.B(n_914),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1087),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1018),
.B(n_918),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1004),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_1080),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1076),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1076),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1087),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1094),
.B(n_921),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_981),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1032),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1023),
.B(n_926),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1032),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1023),
.B(n_927),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1023),
.B(n_928),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1023),
.B(n_929),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1021),
.B(n_931),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1021),
.B(n_932),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_984),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1056),
.B(n_934),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_988),
.B(n_861),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1087),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_984),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1087),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1088),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1021),
.B(n_935),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1088),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1088),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_984),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1088),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1088),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1096),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1096),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1096),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1094),
.B(n_1012),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_984),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1096),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_985),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1096),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1004),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_999),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_999),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1004),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1043),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1043),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1043),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1005),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1043),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1094),
.B(n_936),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1094),
.B(n_985),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1017),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1005),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_990),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_999),
.Y(n_1282)
);

BUFx8_ASAP7_75t_L g1283 ( 
.A(n_1015),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1080),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1058),
.B(n_937),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1005),
.Y(n_1286)
);

AND2x6_ASAP7_75t_L g1287 ( 
.A(n_1048),
.B(n_648),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1021),
.B(n_1093),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_999),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1005),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1058),
.B(n_939),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1048),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1005),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1034),
.A2(n_941),
.B1(n_531),
.B2(n_691),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1067),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1067),
.B(n_950),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1048),
.Y(n_1297)
);

XNOR2xp5_ASAP7_75t_L g1298 ( 
.A(n_1029),
.B(n_827),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1071),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1048),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1057),
.B(n_913),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1051),
.B(n_901),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1055),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1051),
.B(n_901),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1021),
.B(n_1093),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1055),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1071),
.B(n_951),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1021),
.B(n_949),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1045),
.B(n_942),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1055),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1093),
.B(n_949),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1093),
.B(n_969),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1055),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1073),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1009),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1009),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1009),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1078),
.A2(n_913),
.B(n_952),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1073),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1009),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1073),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1009),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1154),
.B(n_912),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1132),
.B(n_1095),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1122),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1279),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1263),
.B(n_1051),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1122),
.B(n_1126),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1098),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1126),
.B(n_1135),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1098),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1100),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1210),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1185),
.Y(n_1334)
);

NAND2xp33_ASAP7_75t_L g1335 ( 
.A(n_1211),
.B(n_1095),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1100),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1130),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1135),
.B(n_1093),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1101),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1249),
.A2(n_1054),
.B1(n_979),
.B2(n_1059),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1301),
.B(n_1057),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1140),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1263),
.B(n_1051),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1185),
.B(n_1008),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1266),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1140),
.B(n_1093),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1130),
.Y(n_1347)
);

NOR2x1p5_ASAP7_75t_L g1348 ( 
.A(n_1249),
.B(n_1061),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1101),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1200),
.A2(n_1073),
.B1(n_1086),
.B2(n_878),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1106),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1266),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1130),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1211),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1200),
.A2(n_1086),
.B1(n_979),
.B2(n_1054),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1106),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1211),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1210),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1200),
.Y(n_1359)
);

BUFx8_ASAP7_75t_SL g1360 ( 
.A(n_1199),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1130),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1272),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1272),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1309),
.B(n_1072),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1188),
.B(n_983),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1273),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1173),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1193),
.A2(n_1086),
.B1(n_960),
.B2(n_973),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1173),
.Y(n_1369)
);

INVx5_ASAP7_75t_L g1370 ( 
.A(n_1211),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1174),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1174),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1273),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1203),
.B(n_983),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1154),
.B(n_1157),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1111),
.B(n_942),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1274),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1274),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1276),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1175),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1153),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1175),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1189),
.B(n_983),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1176),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1111),
.B(n_960),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1176),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1276),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1292),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1278),
.B(n_1068),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1177),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1301),
.B(n_1090),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1153),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1183),
.B(n_973),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1177),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1301),
.B(n_1090),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1193),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1180),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1170),
.B(n_983),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1180),
.Y(n_1399)
);

NAND2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1228),
.B(n_994),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1222),
.B(n_969),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1211),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1237),
.A2(n_1086),
.B1(n_803),
.B2(n_640),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1292),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1297),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1157),
.B(n_912),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1184),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1184),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1211),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1297),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1186),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1300),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1300),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1211),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1278),
.B(n_1068),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1170),
.B(n_995),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1186),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1187),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1303),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1172),
.B(n_995),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1201),
.B(n_1031),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1187),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1303),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1172),
.B(n_1306),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1190),
.A2(n_1061),
.B1(n_865),
.B2(n_1031),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1306),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1310),
.B(n_992),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1295),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1237),
.B(n_527),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1196),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1310),
.B(n_992),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1196),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1277),
.B(n_565),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1198),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1284),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1313),
.B(n_992),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1198),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1222),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1313),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1204),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1102),
.B(n_1008),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_SL g1442 ( 
.A(n_1301),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1223),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1204),
.Y(n_1444)
);

INVx5_ASAP7_75t_L g1445 ( 
.A(n_1223),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1314),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1233),
.B(n_989),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1314),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1163),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1277),
.B(n_568),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1319),
.B(n_992),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1296),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1319),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1295),
.B(n_919),
.Y(n_1454)
);

AND2x6_ASAP7_75t_L g1455 ( 
.A(n_1239),
.B(n_536),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1321),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1296),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1321),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1207),
.Y(n_1459)
);

INVx5_ASAP7_75t_L g1460 ( 
.A(n_1223),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1223),
.A2(n_540),
.B1(n_581),
.B2(n_704),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1207),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1299),
.B(n_653),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1223),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1223),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1299),
.B(n_596),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1223),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1191),
.B(n_995),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1213),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1214),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1213),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1205),
.B(n_954),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1205),
.B(n_956),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1214),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1229),
.B(n_602),
.C(n_600),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1216),
.B(n_893),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1215),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1215),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1287),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1103),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1103),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1285),
.B(n_633),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1217),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1217),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1287),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1218),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1218),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1163),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1110),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1219),
.Y(n_1490)
);

INVxp33_ASAP7_75t_L g1491 ( 
.A(n_1281),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1110),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1113),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1113),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1167),
.B(n_664),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1163),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1219),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1284),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1287),
.A2(n_540),
.B1(n_581),
.B2(n_714),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1285),
.B(n_637),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_L g1501 ( 
.A(n_1287),
.B(n_540),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1285),
.B(n_650),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1115),
.Y(n_1503)
);

BUFx10_ASAP7_75t_L g1504 ( 
.A(n_1287),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1220),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1294),
.A2(n_1025),
.B1(n_571),
.B2(n_729),
.Y(n_1506)
);

AND3x2_ASAP7_75t_L g1507 ( 
.A(n_1134),
.B(n_759),
.C(n_733),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1287),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1296),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1287),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1220),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1115),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1224),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1116),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1104),
.B(n_789),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1116),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1224),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1231),
.B(n_657),
.C(n_654),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1099),
.B(n_666),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1239),
.A2(n_961),
.B(n_958),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1238),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1118),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1307),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1240),
.B(n_1016),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1118),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1238),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1107),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1318),
.B(n_714),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1242),
.B(n_995),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1216),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1119),
.Y(n_1531)
);

AND2x2_ASAP7_75t_SL g1532 ( 
.A(n_1241),
.B(n_733),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1119),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1121),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1121),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1107),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1112),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1127),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1307),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1127),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1307),
.Y(n_1541)
);

BUFx10_ASAP7_75t_L g1542 ( 
.A(n_1099),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1131),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1112),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1114),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1131),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1144),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1241),
.A2(n_540),
.B1(n_581),
.B2(n_734),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_L g1549 ( 
.A(n_1179),
.B(n_540),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1163),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1137),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1137),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1141),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1163),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1168),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1099),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1141),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1136),
.A2(n_1025),
.B1(n_729),
.B2(n_809),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1291),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1114),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1143),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1117),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1243),
.B(n_1016),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1182),
.A2(n_540),
.B1(n_581),
.B2(n_734),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1291),
.Y(n_1565)
);

INVxp67_ASAP7_75t_SL g1566 ( 
.A(n_1168),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1212),
.B(n_793),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1333),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1362),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1530),
.B(n_1171),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1362),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1359),
.B(n_1124),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1479),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1342),
.Y(n_1574)
);

BUFx10_ASAP7_75t_L g1575 ( 
.A(n_1334),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1345),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1367),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1171),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1479),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1556),
.B(n_1171),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1359),
.A2(n_1532),
.B1(n_1396),
.B2(n_1455),
.Y(n_1581)
);

AO22x2_ASAP7_75t_L g1582 ( 
.A1(n_1396),
.A2(n_1302),
.B1(n_1304),
.B2(n_758),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1363),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1556),
.B(n_1248),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1542),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1363),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1370),
.B(n_1145),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1323),
.B(n_1248),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1345),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1367),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1366),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1366),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1369),
.Y(n_1593)
);

CKINVDCx8_ASAP7_75t_R g1594 ( 
.A(n_1334),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1369),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1324),
.B(n_1441),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1323),
.B(n_1248),
.Y(n_1597)
);

BUFx4f_ASAP7_75t_L g1598 ( 
.A(n_1341),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1373),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1352),
.B(n_1318),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1364),
.B(n_1244),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1373),
.Y(n_1602)
);

INVx8_ASAP7_75t_L g1603 ( 
.A(n_1455),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1547),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1370),
.B(n_1133),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1377),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1479),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1377),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1333),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1567),
.B(n_1208),
.C(n_1298),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1532),
.B(n_1117),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1378),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1479),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1371),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1340),
.B(n_1161),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1523),
.B(n_1120),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1325),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1378),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1379),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1360),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1371),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1379),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1387),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1479),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1372),
.Y(n_1625)
);

INVx5_ASAP7_75t_L g1626 ( 
.A(n_1504),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1387),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1342),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1485),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1485),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1388),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1388),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1372),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1498),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1406),
.B(n_1144),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1435),
.B(n_1181),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1404),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1404),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1380),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1406),
.B(n_899),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1405),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1405),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1352),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1485),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1375),
.B(n_957),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1485),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_SL g1647 ( 
.A1(n_1515),
.A2(n_758),
.B1(n_1081),
.B2(n_547),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1376),
.B(n_1120),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1532),
.A2(n_547),
.B1(n_557),
.B2(n_538),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1455),
.A2(n_557),
.B1(n_575),
.B2(n_560),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1341),
.B(n_1152),
.Y(n_1651)
);

OAI22x1_ASAP7_75t_SL g1652 ( 
.A1(n_1326),
.A2(n_1199),
.B1(n_558),
.B2(n_564),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1368),
.A2(n_1128),
.B1(n_1129),
.B2(n_1125),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1355),
.A2(n_560),
.B1(n_583),
.B2(n_575),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1375),
.B(n_1208),
.Y(n_1655)
);

INVx5_ASAP7_75t_L g1656 ( 
.A(n_1504),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1380),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1382),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1410),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1382),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1384),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1370),
.B(n_1125),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1506),
.A2(n_1298),
.B1(n_594),
.B2(n_607),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_SL g1664 ( 
.A(n_1435),
.B(n_1152),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1385),
.B(n_1128),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1498),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1428),
.B(n_1523),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1370),
.B(n_1129),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1370),
.B(n_1139),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1358),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1344),
.Y(n_1671)
);

CKINVDCx8_ASAP7_75t_R g1672 ( 
.A(n_1341),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1370),
.B(n_1139),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1485),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1428),
.B(n_1308),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1329),
.B(n_1142),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1329),
.B(n_1142),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1410),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1510),
.Y(n_1679)
);

INVxp33_ASAP7_75t_L g1680 ( 
.A(n_1454),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1510),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1355),
.B(n_1149),
.Y(n_1682)
);

INVx4_ASAP7_75t_SL g1683 ( 
.A(n_1455),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1559),
.B(n_1311),
.Y(n_1684)
);

INVx8_ASAP7_75t_L g1685 ( 
.A(n_1455),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_L g1686 ( 
.A(n_1445),
.B(n_1133),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1452),
.B(n_1457),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1412),
.Y(n_1688)
);

AND2x2_ASAP7_75t_SL g1689 ( 
.A(n_1335),
.B(n_1368),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1412),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1401),
.B(n_1312),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1413),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1510),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1452),
.B(n_1149),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1331),
.B(n_1151),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1413),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1419),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1419),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1457),
.B(n_1151),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1476),
.B(n_556),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1384),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1510),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1541),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1476),
.B(n_556),
.Y(n_1704)
);

NAND2x1p5_ASAP7_75t_L g1705 ( 
.A(n_1445),
.B(n_1164),
.Y(n_1705)
);

AO22x2_ASAP7_75t_L g1706 ( 
.A1(n_1327),
.A2(n_584),
.B1(n_589),
.B2(n_583),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1463),
.B(n_729),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1423),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1401),
.B(n_1559),
.Y(n_1709)
);

BUFx4f_ASAP7_75t_L g1710 ( 
.A(n_1341),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1423),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1509),
.B(n_1160),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_R g1713 ( 
.A(n_1400),
.B(n_1152),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1426),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1426),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1472),
.B(n_729),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1439),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1509),
.A2(n_1252),
.B1(n_1253),
.B2(n_1250),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1439),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1446),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1565),
.B(n_1317),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1386),
.Y(n_1722)
);

AND2x6_ASAP7_75t_L g1723 ( 
.A(n_1337),
.B(n_1347),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1565),
.B(n_1160),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1438),
.B(n_1164),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1446),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1331),
.B(n_1165),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1386),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1448),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1390),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1541),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1448),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1472),
.B(n_809),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1390),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1442),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1332),
.B(n_1165),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1445),
.B(n_1166),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1539),
.B(n_1473),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1342),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1473),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_L g1741 ( 
.A(n_1354),
.B(n_1166),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1453),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1442),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1394),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1453),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1456),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1507),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1342),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1445),
.B(n_1250),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1456),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1495),
.B(n_809),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1394),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1350),
.A2(n_1253),
.B1(n_1255),
.B2(n_1252),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1510),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1445),
.B(n_1255),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1354),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1491),
.B(n_809),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1458),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1393),
.B(n_1258),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1389),
.B(n_1258),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1539),
.B(n_1315),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1342),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1458),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1527),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1325),
.B(n_1354),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1325),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1542),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1354),
.B(n_1315),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1527),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1415),
.B(n_1259),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1397),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1397),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1445),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1536),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1399),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1332),
.B(n_1259),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1403),
.B(n_817),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1399),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1536),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1537),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1537),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1403),
.B(n_817),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1542),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1544),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1336),
.B(n_1260),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1429),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1544),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1421),
.B(n_1433),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1450),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1545),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1341),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1542),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1545),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1354),
.B(n_1317),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1470),
.Y(n_1795)
);

AND2x6_ASAP7_75t_L g1796 ( 
.A(n_1337),
.B(n_1260),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1560),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1336),
.B(n_817),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1554),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1348),
.Y(n_1800)
);

INVx5_ASAP7_75t_L g1801 ( 
.A(n_1504),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1560),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1348),
.B(n_1320),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1339),
.B(n_1320),
.Y(n_1804)
);

INVx4_ASAP7_75t_SL g1805 ( 
.A(n_1455),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1562),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1470),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1455),
.A2(n_589),
.B1(n_592),
.B2(n_584),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1562),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1482),
.B(n_1164),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1474),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1474),
.Y(n_1812)
);

NAND2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1460),
.B(n_1164),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1339),
.B(n_817),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1477),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1596),
.B(n_1349),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1568),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1585),
.Y(n_1818)
);

AND2x6_ASAP7_75t_L g1819 ( 
.A(n_1573),
.B(n_1409),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1609),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1569),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1596),
.B(n_1349),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1649),
.A2(n_1351),
.B1(n_1469),
.B2(n_1356),
.Y(n_1823)
);

NAND3xp33_ASAP7_75t_L g1824 ( 
.A(n_1751),
.B(n_1615),
.C(n_1610),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1577),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1634),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1577),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1590),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1581),
.B(n_1460),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1571),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1640),
.B(n_1447),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1583),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1586),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1581),
.B(n_1460),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1590),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1648),
.B(n_1665),
.Y(n_1836)
);

NAND2x1_ASAP7_75t_L g1837 ( 
.A(n_1585),
.B(n_1488),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1648),
.B(n_1351),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1788),
.A2(n_1343),
.B1(n_1330),
.B2(n_1328),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1651),
.B(n_1666),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1663),
.A2(n_1558),
.B1(n_1391),
.B2(n_1395),
.C(n_1502),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1649),
.A2(n_1356),
.B1(n_1469),
.B2(n_1408),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1689),
.B(n_1460),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1615),
.A2(n_1518),
.B1(n_1475),
.B2(n_1519),
.Y(n_1844)
);

BUFx12f_ASAP7_75t_L g1845 ( 
.A(n_1620),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1665),
.B(n_1407),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1680),
.B(n_1407),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1680),
.B(n_1408),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1682),
.A2(n_1689),
.B1(n_1759),
.B2(n_1611),
.Y(n_1849)
);

NOR2x1p5_ASAP7_75t_L g1850 ( 
.A(n_1620),
.B(n_1283),
.Y(n_1850)
);

BUFx8_ASAP7_75t_L g1851 ( 
.A(n_1791),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1593),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_L g1853 ( 
.A(n_1573),
.B(n_1460),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_R g1854 ( 
.A(n_1671),
.B(n_1283),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1670),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1593),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1591),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1601),
.A2(n_1518),
.B1(n_1475),
.B2(n_1500),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1682),
.A2(n_1402),
.B1(n_1357),
.B2(n_1350),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1759),
.B(n_1411),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1647),
.A2(n_1411),
.B(n_1418),
.C(n_1417),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1709),
.B(n_1691),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1650),
.A2(n_1417),
.B1(n_1422),
.B2(n_1418),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1570),
.B(n_1422),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1592),
.Y(n_1865)
);

AND2x6_ASAP7_75t_SL g1866 ( 
.A(n_1651),
.B(n_1391),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1709),
.B(n_1430),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1687),
.B(n_1460),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1578),
.B(n_1430),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1687),
.B(n_1357),
.Y(n_1870)
);

AND3x1_ASAP7_75t_L g1871 ( 
.A(n_1655),
.B(n_1635),
.C(n_1664),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1588),
.B(n_1432),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1687),
.B(n_1357),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1597),
.B(n_1432),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1738),
.B(n_1434),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1651),
.B(n_1391),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1667),
.B(n_1391),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1740),
.B(n_1434),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1738),
.B(n_1437),
.Y(n_1879)
);

BUFx5_ASAP7_75t_L g1880 ( 
.A(n_1723),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1773),
.A2(n_1402),
.B(n_1357),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1645),
.B(n_1437),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1707),
.A2(n_1442),
.B1(n_1395),
.B2(n_1391),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1601),
.B(n_1440),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1670),
.B(n_1440),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1765),
.B(n_1402),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1599),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1602),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1595),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1606),
.B(n_1444),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1608),
.B(n_1444),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1612),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_SL g1893 ( 
.A(n_1594),
.B(n_1283),
.Y(n_1893)
);

NOR2x1p5_ASAP7_75t_L g1894 ( 
.A(n_1671),
.B(n_1459),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1773),
.A2(n_1402),
.B(n_1409),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1765),
.B(n_1459),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1786),
.A2(n_1466),
.B1(n_1424),
.B2(n_1462),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1725),
.B(n_1703),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1636),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1618),
.B(n_1462),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1626),
.A2(n_1414),
.B(n_1409),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1619),
.B(n_1471),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1576),
.Y(n_1903)
);

AND2x2_ASAP7_75t_SL g1904 ( 
.A(n_1598),
.B(n_1501),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1604),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1622),
.B(n_1623),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1595),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_1575),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1765),
.B(n_1471),
.Y(n_1909)
);

OAI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1627),
.A2(n_1383),
.B1(n_1395),
.B2(n_1528),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1631),
.B(n_1365),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1684),
.B(n_1414),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1614),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1632),
.B(n_1374),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1614),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1637),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1638),
.B(n_1477),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1684),
.B(n_1414),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1621),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1641),
.B(n_1478),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1700),
.B(n_1395),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1642),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1762),
.Y(n_1923)
);

NAND3xp33_ASAP7_75t_SL g1924 ( 
.A(n_1777),
.B(n_566),
.C(n_563),
.Y(n_1924)
);

INVx4_ASAP7_75t_L g1925 ( 
.A(n_1585),
.Y(n_1925)
);

INVx8_ASAP7_75t_L g1926 ( 
.A(n_1580),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1617),
.A2(n_1464),
.B1(n_1465),
.B2(n_1443),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1617),
.A2(n_1678),
.B1(n_1688),
.B2(n_1659),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1757),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1575),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1690),
.B(n_1478),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1789),
.A2(n_1549),
.B1(n_1443),
.B2(n_1465),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1692),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1650),
.A2(n_1548),
.B1(n_1483),
.B2(n_1486),
.Y(n_1934)
);

OAI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1696),
.A2(n_1395),
.B1(n_1528),
.B2(n_1484),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1580),
.A2(n_1584),
.B1(n_1770),
.B2(n_1760),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1604),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1672),
.B(n_1425),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1697),
.B(n_1483),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1703),
.B(n_1484),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1698),
.B(n_1486),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1739),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1576),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1708),
.B(n_1487),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1580),
.B(n_1443),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1731),
.B(n_1487),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1711),
.B(n_1490),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1714),
.B(n_1490),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1795),
.B(n_1464),
.Y(n_1949)
);

AND2x2_ASAP7_75t_SL g1950 ( 
.A(n_1598),
.B(n_1461),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1715),
.A2(n_1465),
.B1(n_1467),
.B2(n_1464),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1760),
.A2(n_1467),
.B(n_1517),
.C(n_1505),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_R g1953 ( 
.A(n_1735),
.B(n_1467),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1584),
.A2(n_1468),
.B1(n_1529),
.B2(n_1524),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1654),
.A2(n_1526),
.B1(n_1517),
.B2(n_1505),
.C(n_1564),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1717),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1719),
.A2(n_1427),
.B1(n_1436),
.B2(n_1431),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1621),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1720),
.B(n_1526),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1704),
.B(n_1528),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1808),
.A2(n_1782),
.B1(n_1706),
.B2(n_1729),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1726),
.B(n_1563),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1625),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1732),
.B(n_1551),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1742),
.B(n_1746),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1745),
.B(n_1551),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1589),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1589),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1750),
.B(n_1552),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1758),
.B(n_1552),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1763),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1625),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1731),
.B(n_1470),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1716),
.B(n_1557),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1733),
.B(n_1557),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1770),
.B(n_1561),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1795),
.B(n_1504),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1633),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1724),
.B(n_1561),
.Y(n_1979)
);

INVx4_ASAP7_75t_L g1980 ( 
.A(n_1573),
.Y(n_1980)
);

AND3x1_ASAP7_75t_L g1981 ( 
.A(n_1747),
.B(n_1069),
.C(n_597),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1764),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1808),
.A2(n_1528),
.B1(n_1499),
.B2(n_597),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1706),
.A2(n_1528),
.B1(n_598),
.B2(n_599),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1706),
.A2(n_598),
.B1(n_599),
.B2(n_592),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1799),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1798),
.B(n_1347),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1633),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1639),
.A2(n_605),
.B1(n_608),
.B2(n_604),
.Y(n_1989)
);

INVxp67_ASAP7_75t_SL g1990 ( 
.A(n_1799),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1639),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1769),
.B(n_1774),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1724),
.B(n_1497),
.Y(n_1993)
);

BUFx12f_ASAP7_75t_SL g1994 ( 
.A(n_1803),
.Y(n_1994)
);

OR2x6_ASAP7_75t_L g1995 ( 
.A(n_1603),
.B(n_1353),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1814),
.B(n_1353),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1779),
.B(n_1511),
.Y(n_1997)
);

NOR2x2_ASAP7_75t_L g1998 ( 
.A(n_1657),
.B(n_1069),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1780),
.B(n_1497),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1781),
.B(n_1497),
.Y(n_2000)
);

AND2x6_ASAP7_75t_SL g2001 ( 
.A(n_1652),
.B(n_604),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1667),
.B(n_1511),
.Y(n_2002)
);

A2O1A1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_1776),
.A2(n_1398),
.B(n_1513),
.C(n_1511),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1643),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1784),
.B(n_1513),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1787),
.B(n_1513),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1584),
.A2(n_1420),
.B1(n_1416),
.B2(n_1451),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1790),
.B(n_1793),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1807),
.B(n_1508),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1657),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1797),
.B(n_1521),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1723),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1802),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1806),
.B(n_1521),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1809),
.B(n_1521),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1658),
.A2(n_608),
.B1(n_614),
.B2(n_605),
.Y(n_2016)
);

AND2x6_ASAP7_75t_SL g2017 ( 
.A(n_1803),
.B(n_614),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1762),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1811),
.B(n_1480),
.Y(n_2019)
);

BUFx12f_ASAP7_75t_L g2020 ( 
.A(n_1735),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1675),
.A2(n_1582),
.B1(n_1616),
.B2(n_1600),
.Y(n_2021)
);

NAND2xp33_ASAP7_75t_L g2022 ( 
.A(n_1573),
.B(n_1554),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1812),
.B(n_1480),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1658),
.A2(n_631),
.B1(n_632),
.B2(n_630),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1739),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1815),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1626),
.A2(n_1496),
.B(n_1488),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1579),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1825),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1877),
.B(n_1643),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1821),
.Y(n_2031)
);

BUFx5_ASAP7_75t_L g2032 ( 
.A(n_1819),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1818),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_2012),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1827),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1836),
.B(n_1849),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1905),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_1820),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_2012),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_2012),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1828),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1942),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1817),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1862),
.B(n_1675),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1859),
.B(n_1600),
.Y(n_2045)
);

INVx5_ASAP7_75t_L g2046 ( 
.A(n_1819),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1830),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_SL g2048 ( 
.A(n_1893),
.B(n_1743),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1862),
.B(n_1582),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1835),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1852),
.Y(n_2051)
);

BUFx3_ASAP7_75t_L g2052 ( 
.A(n_1826),
.Y(n_2052)
);

AO22x1_ASAP7_75t_L g2053 ( 
.A1(n_1831),
.A2(n_1743),
.B1(n_1800),
.B2(n_1721),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1832),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1845),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1847),
.B(n_1582),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1816),
.B(n_1721),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1824),
.A2(n_1661),
.B1(n_1701),
.B2(n_1660),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_1818),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1822),
.B(n_1734),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1833),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1924),
.A2(n_1710),
.B1(n_1616),
.B2(n_1761),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1857),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_1899),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1854),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1865),
.Y(n_2066)
);

CKINVDCx6p67_ASAP7_75t_R g2067 ( 
.A(n_2020),
.Y(n_2067)
);

INVx5_ASAP7_75t_L g2068 ( 
.A(n_1819),
.Y(n_2068)
);

CKINVDCx20_ASAP7_75t_R g2069 ( 
.A(n_1854),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1887),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1925),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1877),
.B(n_1783),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_1943),
.B(n_1783),
.Y(n_2073)
);

NOR2xp67_ASAP7_75t_L g2074 ( 
.A(n_1929),
.B(n_1810),
.Y(n_2074)
);

AOI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1871),
.A2(n_1921),
.B1(n_1938),
.B2(n_1960),
.Y(n_2075)
);

INVx2_ASAP7_75t_SL g2076 ( 
.A(n_1968),
.Y(n_2076)
);

INVx5_ASAP7_75t_L g2077 ( 
.A(n_1819),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1888),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1847),
.B(n_1660),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1841),
.A2(n_1710),
.B1(n_1616),
.B2(n_1761),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1856),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1892),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_2012),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1942),
.Y(n_2084)
);

BUFx12f_ASAP7_75t_L g2085 ( 
.A(n_1866),
.Y(n_2085)
);

AND3x1_ASAP7_75t_SL g2086 ( 
.A(n_1894),
.B(n_1850),
.C(n_631),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_1908),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_SL g2088 ( 
.A1(n_1950),
.A2(n_1713),
.B1(n_1603),
.B2(n_1685),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1848),
.B(n_1661),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1930),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1916),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1926),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1851),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1889),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1907),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1925),
.Y(n_2096)
);

CKINVDCx20_ASAP7_75t_R g2097 ( 
.A(n_1937),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1922),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1933),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_1882),
.B(n_1701),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1848),
.B(n_1722),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1838),
.B(n_1722),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1980),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1936),
.B(n_1730),
.Y(n_2104)
);

INVxp67_ASAP7_75t_SL g2105 ( 
.A(n_2022),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_1844),
.A2(n_1761),
.B1(n_1694),
.B2(n_1712),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2002),
.B(n_1768),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1851),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1884),
.B(n_1771),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1913),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1884),
.B(n_1730),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_1855),
.B(n_1807),
.Y(n_2112)
);

INVx4_ASAP7_75t_L g2113 ( 
.A(n_1926),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1915),
.Y(n_2114)
);

INVx3_ASAP7_75t_L g2115 ( 
.A(n_1980),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1903),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1919),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_1898),
.B(n_1572),
.Y(n_2118)
);

HB1xp67_ASAP7_75t_L g2119 ( 
.A(n_2025),
.Y(n_2119)
);

AND3x1_ASAP7_75t_L g2120 ( 
.A(n_1967),
.B(n_632),
.C(n_630),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1958),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1867),
.B(n_1778),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2025),
.Y(n_2123)
);

INVx3_ASAP7_75t_L g2124 ( 
.A(n_2002),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1956),
.Y(n_2125)
);

NOR2xp67_ASAP7_75t_L g2126 ( 
.A(n_2004),
.B(n_1574),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_1994),
.Y(n_2127)
);

AOI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_1981),
.A2(n_1694),
.B1(n_1712),
.B2(n_1699),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1971),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1982),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_1840),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1840),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_L g2133 ( 
.A1(n_1985),
.A2(n_1734),
.B1(n_1744),
.B2(n_1728),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_1998),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1963),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1858),
.A2(n_1694),
.B1(n_1712),
.B2(n_1699),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1972),
.Y(n_2137)
);

INVx5_ASAP7_75t_L g2138 ( 
.A(n_1819),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1885),
.B(n_1804),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1978),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1898),
.B(n_1572),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2013),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1867),
.B(n_1728),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2026),
.Y(n_2144)
);

OR2x4_ASAP7_75t_L g2145 ( 
.A(n_1940),
.B(n_1579),
.Y(n_2145)
);

BUFx2_ASAP7_75t_L g2146 ( 
.A(n_1840),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_2017),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1988),
.Y(n_2148)
);

HB1xp67_ASAP7_75t_SL g2149 ( 
.A(n_1885),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1926),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1991),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_1940),
.B(n_1946),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_1946),
.B(n_1878),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1995),
.Y(n_2154)
);

AND2x4_ASAP7_75t_SL g2155 ( 
.A(n_1995),
.B(n_1579),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_1876),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1878),
.B(n_1699),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2010),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1906),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1995),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1923),
.Y(n_2161)
);

AND2x6_ASAP7_75t_L g2162 ( 
.A(n_1987),
.B(n_1579),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_1883),
.A2(n_1741),
.B1(n_1628),
.B2(n_1574),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_1875),
.B(n_1744),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_1985),
.A2(n_1771),
.B1(n_1772),
.B2(n_1752),
.Y(n_2165)
);

INVx2_ASAP7_75t_SL g2166 ( 
.A(n_1876),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1879),
.B(n_1804),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1880),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1965),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2008),
.Y(n_2170)
);

AOI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_1853),
.A2(n_1656),
.B(n_1626),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_2028),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1961),
.B(n_1804),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_1876),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_1953),
.Y(n_2175)
);

CKINVDCx20_ASAP7_75t_R g2176 ( 
.A(n_2021),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1872),
.B(n_1752),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_1953),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1874),
.B(n_1772),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1923),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1839),
.A2(n_1741),
.B1(n_1748),
.B2(n_1628),
.Y(n_2181)
);

AND2x4_ASAP7_75t_SL g2182 ( 
.A(n_2018),
.B(n_1607),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_2001),
.Y(n_2183)
);

BUFx4f_ASAP7_75t_L g2184 ( 
.A(n_1904),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1964),
.Y(n_2185)
);

INVxp67_ASAP7_75t_SL g2186 ( 
.A(n_1986),
.Y(n_2186)
);

INVx2_ASAP7_75t_SL g2187 ( 
.A(n_1973),
.Y(n_2187)
);

INVx3_ASAP7_75t_L g2188 ( 
.A(n_2018),
.Y(n_2188)
);

BUFx4f_ASAP7_75t_L g2189 ( 
.A(n_1904),
.Y(n_2189)
);

BUFx4f_ASAP7_75t_L g2190 ( 
.A(n_1950),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1966),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1969),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1846),
.B(n_1775),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1970),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_2028),
.Y(n_2195)
);

NAND2x1p5_ASAP7_75t_L g2196 ( 
.A(n_1837),
.B(n_1767),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1973),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1880),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2019),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_1868),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1974),
.B(n_1775),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1860),
.B(n_1778),
.Y(n_2202)
);

NOR2x1_ASAP7_75t_L g2203 ( 
.A(n_1992),
.B(n_1748),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_1975),
.B(n_1676),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1961),
.B(n_1713),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1864),
.B(n_1776),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1897),
.B(n_1767),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1868),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2023),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1843),
.A2(n_1992),
.B1(n_1869),
.B2(n_1935),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1880),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1996),
.B(n_1723),
.Y(n_2212)
);

AOI211xp5_ASAP7_75t_L g2213 ( 
.A1(n_1935),
.A2(n_642),
.B(n_651),
.C(n_641),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1880),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1886),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1880),
.Y(n_2216)
);

CKINVDCx20_ASAP7_75t_R g2217 ( 
.A(n_1843),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1890),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_1945),
.B(n_1768),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_1984),
.A2(n_1983),
.B1(n_2016),
.B2(n_1989),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_1917),
.B(n_1766),
.Y(n_2221)
);

NAND3xp33_ASAP7_75t_SL g2222 ( 
.A(n_1984),
.B(n_572),
.C(n_570),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1891),
.Y(n_2223)
);

INVxp67_ASAP7_75t_L g2224 ( 
.A(n_1896),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1900),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1911),
.B(n_1723),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1886),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_1986),
.Y(n_2228)
);

OR2x4_ASAP7_75t_L g2229 ( 
.A(n_1920),
.B(n_1607),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_1880),
.Y(n_2230)
);

AND3x1_ASAP7_75t_L g2231 ( 
.A(n_1989),
.B(n_642),
.C(n_641),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1997),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1902),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_1990),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1931),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_1990),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_1896),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_1939),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1999),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1914),
.B(n_1962),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_1909),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1823),
.B(n_1723),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1941),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2016),
.B(n_1768),
.Y(n_2244)
);

AOI22xp33_ASAP7_75t_L g2245 ( 
.A1(n_1983),
.A2(n_768),
.B1(n_786),
.B2(n_759),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_1909),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2007),
.B(n_1792),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_L g2248 ( 
.A(n_1944),
.B(n_1766),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2000),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1823),
.B(n_1677),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_1912),
.B(n_1794),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1947),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1910),
.B(n_1954),
.Y(n_2253)
);

BUFx3_ASAP7_75t_L g2254 ( 
.A(n_1948),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1912),
.B(n_1794),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_1932),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2005),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_1870),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2006),
.Y(n_2259)
);

CKINVDCx11_ASAP7_75t_R g2260 ( 
.A(n_1928),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2149),
.B(n_1918),
.Y(n_2261)
);

A2O1A1Ixp33_ASAP7_75t_L g2262 ( 
.A1(n_2190),
.A2(n_1861),
.B(n_1834),
.C(n_1829),
.Y(n_2262)
);

AOI221xp5_ASAP7_75t_L g2263 ( 
.A1(n_2036),
.A2(n_2220),
.B1(n_2231),
.B2(n_2222),
.C(n_2253),
.Y(n_2263)
);

O2A1O1Ixp33_ASAP7_75t_L g2264 ( 
.A1(n_2036),
.A2(n_1910),
.B(n_1952),
.C(n_652),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2029),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_2152),
.B(n_1918),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2152),
.B(n_1959),
.Y(n_2267)
);

AOI21xp5_ASAP7_75t_L g2268 ( 
.A1(n_2105),
.A2(n_2240),
.B(n_2171),
.Y(n_2268)
);

INVx2_ASAP7_75t_SL g2269 ( 
.A(n_2043),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2043),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2075),
.A2(n_1870),
.B1(n_1873),
.B2(n_1955),
.Y(n_2271)
);

O2A1O1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_2253),
.A2(n_652),
.B(n_655),
.C(n_651),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2118),
.B(n_1976),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2153),
.B(n_1842),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2105),
.A2(n_1834),
.B(n_1829),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_2052),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2118),
.B(n_1979),
.Y(n_2277)
);

AO21x2_ASAP7_75t_L g2278 ( 
.A1(n_2247),
.A2(n_2003),
.B(n_1977),
.Y(n_2278)
);

BUFx2_ASAP7_75t_L g2279 ( 
.A(n_2052),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2141),
.B(n_1842),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2045),
.A2(n_1873),
.B(n_2027),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_L g2282 ( 
.A(n_2038),
.B(n_2153),
.Y(n_2282)
);

INVx3_ASAP7_75t_SL g2283 ( 
.A(n_2067),
.Y(n_2283)
);

AO21x2_ASAP7_75t_L g2284 ( 
.A1(n_2247),
.A2(n_2009),
.B(n_1977),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2141),
.B(n_1993),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2206),
.B(n_2011),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_2064),
.B(n_2134),
.Y(n_2287)
);

NAND2xp33_ASAP7_75t_SL g2288 ( 
.A(n_2069),
.B(n_1607),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2031),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2092),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2056),
.B(n_2024),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_2045),
.A2(n_1656),
.B(n_1626),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2190),
.B(n_2014),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2159),
.B(n_2024),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2139),
.B(n_1794),
.Y(n_2295)
);

OR2x6_ASAP7_75t_L g2296 ( 
.A(n_2156),
.B(n_2009),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2047),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_2092),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2169),
.B(n_672),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2186),
.A2(n_1801),
.B(n_1656),
.Y(n_2300)
);

A2O1A1Ixp33_ASAP7_75t_L g2301 ( 
.A1(n_2220),
.A2(n_1934),
.B(n_1603),
.C(n_1685),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2054),
.Y(n_2302)
);

OR2x6_ASAP7_75t_SL g2303 ( 
.A(n_2065),
.B(n_574),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2029),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2035),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2061),
.Y(n_2306)
);

A2O1A1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2213),
.A2(n_1934),
.B(n_1685),
.C(n_1863),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2042),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2260),
.A2(n_1957),
.B1(n_1753),
.B2(n_1653),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2238),
.B(n_655),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2035),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2170),
.B(n_2235),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2063),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2243),
.B(n_1863),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_SL g2315 ( 
.A(n_2037),
.B(n_1607),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2186),
.A2(n_1801),
.B(n_1656),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_L g2317 ( 
.A(n_2037),
.B(n_676),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2252),
.B(n_2015),
.Y(n_2318)
);

AOI21x1_ASAP7_75t_L g2319 ( 
.A1(n_2207),
.A2(n_1785),
.B(n_1520),
.Y(n_2319)
);

O2A1O1Ixp33_ASAP7_75t_L g2320 ( 
.A1(n_2049),
.A2(n_661),
.B(n_665),
.C(n_658),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2122),
.B(n_1695),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2044),
.B(n_1481),
.Y(n_2322)
);

A2O1A1Ixp33_ASAP7_75t_L g2323 ( 
.A1(n_2080),
.A2(n_1718),
.B(n_1792),
.C(n_1881),
.Y(n_2323)
);

AOI21x1_ASAP7_75t_L g2324 ( 
.A1(n_2207),
.A2(n_2060),
.B(n_2104),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2066),
.Y(n_2325)
);

INVxp67_ASAP7_75t_L g2326 ( 
.A(n_2076),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2034),
.Y(n_2327)
);

AO22x1_ASAP7_75t_L g2328 ( 
.A1(n_2205),
.A2(n_580),
.B1(n_586),
.B2(n_578),
.Y(n_2328)
);

A2O1A1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2184),
.A2(n_1901),
.B(n_1727),
.C(n_1736),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2097),
.B(n_677),
.Y(n_2330)
);

A2O1A1Ixp33_ASAP7_75t_L g2331 ( 
.A1(n_2184),
.A2(n_1895),
.B(n_1949),
.C(n_1587),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_2087),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_2092),
.Y(n_2333)
);

OAI33xp33_ASAP7_75t_L g2334 ( 
.A1(n_2070),
.A2(n_593),
.A3(n_590),
.B1(n_601),
.B2(n_591),
.B3(n_588),
.Y(n_2334)
);

INVx1_ASAP7_75t_SL g2335 ( 
.A(n_2097),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_2250),
.A2(n_1801),
.B(n_1587),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2143),
.B(n_1796),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2102),
.A2(n_1801),
.B(n_1496),
.Y(n_2338)
);

OAI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2145),
.A2(n_1624),
.B1(n_1629),
.B2(n_1613),
.Y(n_2339)
);

BUFx4f_ASAP7_75t_L g2340 ( 
.A(n_2092),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2145),
.A2(n_1624),
.B1(n_1629),
.B2(n_1613),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2189),
.B(n_1799),
.Y(n_2342)
);

NAND2x1p5_ASAP7_75t_L g2343 ( 
.A(n_2046),
.B(n_1799),
.Y(n_2343)
);

INVx1_ASAP7_75t_SL g2344 ( 
.A(n_2234),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2042),
.B(n_1949),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2078),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_2055),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_SL g2348 ( 
.A(n_2048),
.B(n_2069),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2189),
.B(n_1613),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2111),
.A2(n_1496),
.B(n_1488),
.Y(n_2350)
);

O2A1O1Ixp5_ASAP7_75t_L g2351 ( 
.A1(n_2053),
.A2(n_1927),
.B(n_1951),
.C(n_1668),
.Y(n_2351)
);

AOI221xp5_ASAP7_75t_L g2352 ( 
.A1(n_2120),
.A2(n_610),
.B1(n_612),
.B2(n_609),
.C(n_606),
.Y(n_2352)
);

OAI21x1_ASAP7_75t_L g2353 ( 
.A1(n_2198),
.A2(n_1392),
.B(n_1381),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_L g2354 ( 
.A(n_2147),
.B(n_661),
.C(n_658),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2082),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_2087),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2091),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2254),
.B(n_1613),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2084),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2030),
.Y(n_2360)
);

OAI22x1_ASAP7_75t_L g2361 ( 
.A1(n_2166),
.A2(n_667),
.B1(n_669),
.B2(n_665),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2057),
.B(n_1796),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2109),
.B(n_1796),
.Y(n_2363)
);

NOR3xp33_ASAP7_75t_SL g2364 ( 
.A(n_2183),
.B(n_615),
.C(n_613),
.Y(n_2364)
);

CKINVDCx14_ASAP7_75t_R g2365 ( 
.A(n_2108),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2218),
.B(n_1481),
.Y(n_2366)
);

O2A1O1Ixp5_ASAP7_75t_L g2367 ( 
.A1(n_2104),
.A2(n_1668),
.B(n_1669),
.C(n_1662),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2030),
.B(n_667),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2254),
.B(n_2157),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_2111),
.A2(n_1496),
.B(n_1488),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2223),
.B(n_2225),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2098),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_R g2373 ( 
.A(n_2090),
.B(n_2256),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2157),
.B(n_1624),
.Y(n_2374)
);

OAI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2210),
.A2(n_2136),
.B1(n_2176),
.B2(n_2217),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2034),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2060),
.A2(n_1392),
.B(n_1381),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2127),
.Y(n_2378)
);

CKINVDCx20_ASAP7_75t_R g2379 ( 
.A(n_2086),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2187),
.B(n_1624),
.Y(n_2380)
);

OAI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2176),
.A2(n_1630),
.B1(n_1644),
.B2(n_1629),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_2124),
.B(n_680),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2233),
.B(n_1796),
.Y(n_2383)
);

INVx3_ASAP7_75t_SL g2384 ( 
.A(n_2093),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2185),
.B(n_1796),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2099),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_L g2387 ( 
.A(n_2260),
.B(n_673),
.C(n_669),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2062),
.A2(n_2174),
.B1(n_2132),
.B2(n_2086),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2193),
.A2(n_1392),
.B(n_1381),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_2202),
.A2(n_1566),
.B(n_1550),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_2034),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2191),
.B(n_1361),
.Y(n_2392)
);

OAI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_2217),
.A2(n_1630),
.B1(n_1644),
.B2(n_1629),
.Y(n_2393)
);

NOR3xp33_ASAP7_75t_SL g2394 ( 
.A(n_2112),
.B(n_622),
.C(n_620),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2125),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2041),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_2084),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_SL g2398 ( 
.A1(n_2085),
.A2(n_624),
.B1(n_625),
.B2(n_623),
.Y(n_2398)
);

HB1xp67_ASAP7_75t_L g2399 ( 
.A(n_2119),
.Y(n_2399)
);

NAND3xp33_ASAP7_75t_SL g2400 ( 
.A(n_2128),
.B(n_635),
.C(n_628),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_2124),
.B(n_693),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2226),
.A2(n_1644),
.B(n_1630),
.Y(n_2402)
);

AOI21xp33_ASAP7_75t_L g2403 ( 
.A1(n_2204),
.A2(n_1492),
.B(n_1489),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2107),
.B(n_696),
.Y(n_2404)
);

AOI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_2046),
.A2(n_1644),
.B(n_1630),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2215),
.B(n_1646),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_2034),
.Y(n_2407)
);

A2O1A1Ixp33_ASAP7_75t_SL g2408 ( 
.A1(n_2201),
.A2(n_1553),
.B(n_1531),
.C(n_1489),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2197),
.B(n_673),
.Y(n_2409)
);

INVx4_ASAP7_75t_L g2410 ( 
.A(n_2039),
.Y(n_2410)
);

AO22x1_ASAP7_75t_L g2411 ( 
.A1(n_2090),
.A2(n_636),
.B1(n_638),
.B2(n_629),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2129),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2107),
.B(n_697),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2072),
.B(n_1646),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2041),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2046),
.A2(n_2077),
.B(n_2068),
.Y(n_2416)
);

AO32x2_ASAP7_75t_L g2417 ( 
.A1(n_2237),
.A2(n_1520),
.A3(n_706),
.B1(n_707),
.B2(n_694),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2192),
.B(n_1361),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2175),
.B(n_710),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_2072),
.B(n_1646),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2215),
.B(n_1646),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2050),
.Y(n_2422)
);

O2A1O1Ixp33_ASAP7_75t_L g2423 ( 
.A1(n_2197),
.A2(n_694),
.B(n_706),
.C(n_681),
.Y(n_2423)
);

OA22x2_ASAP7_75t_L g2424 ( 
.A1(n_2119),
.A2(n_707),
.B1(n_713),
.B2(n_681),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2050),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2123),
.B(n_713),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2194),
.B(n_1492),
.Y(n_2427)
);

INVx1_ASAP7_75t_SL g2428 ( 
.A(n_2116),
.Y(n_2428)
);

OAI21x1_ASAP7_75t_L g2429 ( 
.A1(n_2198),
.A2(n_1813),
.B(n_1705),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2123),
.B(n_716),
.Y(n_2430)
);

OR2x2_ASAP7_75t_L g2431 ( 
.A(n_2100),
.B(n_1493),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_SL g2432 ( 
.A(n_2215),
.B(n_1674),
.Y(n_2432)
);

NAND2xp33_ASAP7_75t_R g2433 ( 
.A(n_2131),
.B(n_736),
.Y(n_2433)
);

AO21x1_ASAP7_75t_L g2434 ( 
.A1(n_2221),
.A2(n_1813),
.B(n_1705),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2112),
.B(n_740),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2106),
.A2(n_1679),
.B1(n_1681),
.B2(n_1674),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2199),
.B(n_1493),
.Y(n_2437)
);

AOI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2046),
.A2(n_2077),
.B(n_2068),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2228),
.Y(n_2439)
);

AOI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_2068),
.A2(n_1679),
.B(n_1674),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_R g2441 ( 
.A(n_2178),
.B(n_1674),
.Y(n_2441)
);

O2A1O1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_2146),
.A2(n_718),
.B(n_720),
.C(n_716),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2068),
.A2(n_1681),
.B(n_1679),
.Y(n_2443)
);

AO21x1_ASAP7_75t_L g2444 ( 
.A1(n_2221),
.A2(n_1669),
.B(n_1662),
.Y(n_2444)
);

O2A1O1Ixp33_ASAP7_75t_L g2445 ( 
.A1(n_2224),
.A2(n_720),
.B(n_723),
.C(n_718),
.Y(n_2445)
);

O2A1O1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2209),
.A2(n_2142),
.B(n_2144),
.C(n_2130),
.Y(n_2446)
);

O2A1O1Ixp33_ASAP7_75t_L g2447 ( 
.A1(n_2241),
.A2(n_726),
.B(n_727),
.C(n_723),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2079),
.B(n_1494),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2077),
.A2(n_1681),
.B(n_1679),
.Y(n_2449)
);

HB1xp67_ASAP7_75t_L g2450 ( 
.A(n_2236),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2051),
.Y(n_2451)
);

BUFx2_ASAP7_75t_L g2452 ( 
.A(n_2073),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2077),
.A2(n_1693),
.B(n_1681),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2215),
.B(n_1693),
.Y(n_2454)
);

AOI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2085),
.A2(n_778),
.B1(n_779),
.B2(n_761),
.Y(n_2455)
);

O2A1O1Ixp33_ASAP7_75t_L g2456 ( 
.A1(n_2246),
.A2(n_727),
.B(n_735),
.C(n_726),
.Y(n_2456)
);

O2A1O1Ixp33_ASAP7_75t_SL g2457 ( 
.A1(n_2089),
.A2(n_1737),
.B(n_1673),
.C(n_1749),
.Y(n_2457)
);

INVx2_ASAP7_75t_SL g2458 ( 
.A(n_2108),
.Y(n_2458)
);

INVx1_ASAP7_75t_SL g2459 ( 
.A(n_2073),
.Y(n_2459)
);

O2A1O1Ixp33_ASAP7_75t_L g2460 ( 
.A1(n_2101),
.A2(n_747),
.B(n_753),
.C(n_735),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2167),
.B(n_747),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2173),
.B(n_753),
.Y(n_2462)
);

O2A1O1Ixp33_ASAP7_75t_SL g2463 ( 
.A1(n_2242),
.A2(n_1737),
.B(n_1673),
.C(n_1749),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2201),
.B(n_1494),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_L g2465 ( 
.A(n_2200),
.B(n_780),
.Y(n_2465)
);

BUFx2_ASAP7_75t_L g2466 ( 
.A(n_2229),
.Y(n_2466)
);

NAND2x1p5_ASAP7_75t_L g2467 ( 
.A(n_2138),
.B(n_2154),
.Y(n_2467)
);

INVx3_ASAP7_75t_SL g2468 ( 
.A(n_2113),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2177),
.B(n_1503),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2051),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2150),
.B(n_1693),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2150),
.B(n_1693),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_SL g2473 ( 
.A(n_2245),
.B(n_646),
.C(n_639),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2081),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2138),
.A2(n_1754),
.B(n_1702),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2081),
.Y(n_2476)
);

OR2x6_ASAP7_75t_L g2477 ( 
.A(n_2258),
.B(n_1702),
.Y(n_2477)
);

A2O1A1Ixp33_ASAP7_75t_L g2478 ( 
.A1(n_2074),
.A2(n_1754),
.B(n_1756),
.C(n_1702),
.Y(n_2478)
);

OAI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2245),
.A2(n_1754),
.B1(n_1756),
.B2(n_1702),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2232),
.B(n_1503),
.Y(n_2480)
);

INVx4_ASAP7_75t_L g2481 ( 
.A(n_2039),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2244),
.B(n_2219),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2219),
.B(n_760),
.Y(n_2483)
);

AOI21xp5_ASAP7_75t_L g2484 ( 
.A1(n_2138),
.A2(n_1756),
.B(n_1754),
.Y(n_2484)
);

HB1xp67_ASAP7_75t_L g2485 ( 
.A(n_2229),
.Y(n_2485)
);

OAI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2133),
.A2(n_1756),
.B1(n_765),
.B2(n_774),
.Y(n_2486)
);

O2A1O1Ixp33_ASAP7_75t_L g2487 ( 
.A1(n_2248),
.A2(n_765),
.B(n_774),
.C(n_760),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2094),
.Y(n_2488)
);

A2O1A1Ixp33_ASAP7_75t_L g2489 ( 
.A1(n_2177),
.A2(n_776),
.B(n_799),
.C(n_794),
.Y(n_2489)
);

AOI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2088),
.A2(n_797),
.B1(n_800),
.B2(n_781),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2094),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2200),
.B(n_801),
.Y(n_2492)
);

OAI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2133),
.A2(n_2165),
.B1(n_2138),
.B2(n_2179),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2095),
.Y(n_2494)
);

AOI22x1_ASAP7_75t_L g2495 ( 
.A1(n_2232),
.A2(n_1514),
.B1(n_1516),
.B2(n_1512),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2200),
.B(n_805),
.Y(n_2496)
);

AOI21xp5_ASAP7_75t_L g2497 ( 
.A1(n_2248),
.A2(n_1755),
.B(n_1686),
.Y(n_2497)
);

O2A1O1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_2179),
.A2(n_776),
.B(n_799),
.C(n_794),
.Y(n_2498)
);

OAI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2165),
.A2(n_819),
.B1(n_820),
.B2(n_812),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2239),
.A2(n_2249),
.B1(n_2259),
.B2(n_2257),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2095),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2110),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2239),
.B(n_1512),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2172),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2110),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2249),
.B(n_1514),
.Y(n_2506)
);

BUFx2_ASAP7_75t_L g2507 ( 
.A(n_2195),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2114),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2257),
.B(n_1516),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2114),
.Y(n_2510)
);

AND2x4_ASAP7_75t_L g2511 ( 
.A(n_2113),
.B(n_1683),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2259),
.B(n_1522),
.Y(n_2512)
);

NOR3xp33_ASAP7_75t_L g2513 ( 
.A(n_2154),
.B(n_819),
.C(n_812),
.Y(n_2513)
);

BUFx2_ASAP7_75t_L g2514 ( 
.A(n_2195),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2200),
.B(n_644),
.Y(n_2515)
);

A2O1A1Ixp33_ASAP7_75t_SL g2516 ( 
.A1(n_2160),
.A2(n_1553),
.B(n_1531),
.C(n_1522),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2251),
.B(n_958),
.Y(n_2517)
);

AOI21xp5_ASAP7_75t_L g2518 ( 
.A1(n_2212),
.A2(n_1755),
.B(n_1686),
.Y(n_2518)
);

INVxp67_ASAP7_75t_SL g2519 ( 
.A(n_2164),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2227),
.B(n_1683),
.Y(n_2520)
);

OAI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_2181),
.A2(n_1533),
.B(n_1525),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2117),
.Y(n_2522)
);

BUFx3_ASAP7_75t_L g2523 ( 
.A(n_2172),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2039),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_2208),
.B(n_647),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2276),
.Y(n_2526)
);

INVx2_ASAP7_75t_SL g2527 ( 
.A(n_2356),
.Y(n_2527)
);

INVx3_ASAP7_75t_L g2528 ( 
.A(n_2504),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2265),
.Y(n_2529)
);

OAI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2274),
.A2(n_2058),
.B1(n_2163),
.B2(n_2227),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2482),
.B(n_2251),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2373),
.Y(n_2532)
);

OR2x6_ASAP7_75t_L g2533 ( 
.A(n_2268),
.B(n_2258),
.Y(n_2533)
);

OAI22xp5_ASAP7_75t_L g2534 ( 
.A1(n_2307),
.A2(n_2058),
.B1(n_2227),
.B2(n_2258),
.Y(n_2534)
);

BUFx8_ASAP7_75t_L g2535 ( 
.A(n_2279),
.Y(n_2535)
);

OAI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2348),
.A2(n_2375),
.B1(n_2263),
.B2(n_2388),
.Y(n_2536)
);

AND2x4_ASAP7_75t_L g2537 ( 
.A(n_2466),
.B(n_2485),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2273),
.B(n_2208),
.Y(n_2538)
);

AOI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2300),
.A2(n_2214),
.B(n_2230),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2289),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2347),
.Y(n_2541)
);

INVx4_ASAP7_75t_L g2542 ( 
.A(n_2356),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2387),
.A2(n_2208),
.B1(n_2227),
.B2(n_2258),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_2356),
.Y(n_2544)
);

INVx1_ASAP7_75t_SL g2545 ( 
.A(n_2439),
.Y(n_2545)
);

OAI22xp5_ASAP7_75t_L g2546 ( 
.A1(n_2309),
.A2(n_2280),
.B1(n_2301),
.B2(n_2375),
.Y(n_2546)
);

O2A1O1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2267),
.A2(n_786),
.B(n_787),
.C(n_768),
.Y(n_2547)
);

XOR2xp5_ASAP7_75t_L g2548 ( 
.A(n_2365),
.B(n_2208),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2312),
.B(n_2203),
.Y(n_2549)
);

BUFx2_ASAP7_75t_L g2550 ( 
.A(n_2452),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2273),
.B(n_2117),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2507),
.B(n_2160),
.Y(n_2552)
);

AOI221x1_ASAP7_75t_L g2553 ( 
.A1(n_2513),
.A2(n_2255),
.B1(n_821),
.B2(n_808),
.C(n_787),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2304),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_2270),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_L g2556 ( 
.A(n_2335),
.B(n_2172),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2297),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2285),
.B(n_2277),
.Y(n_2558)
);

AO32x1_ASAP7_75t_L g2559 ( 
.A1(n_2493),
.A2(n_2216),
.A3(n_2211),
.B1(n_2168),
.B2(n_2121),
.Y(n_2559)
);

CKINVDCx20_ASAP7_75t_R g2560 ( 
.A(n_2283),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2462),
.B(n_2517),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2308),
.B(n_2121),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2316),
.A2(n_2214),
.B(n_2230),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2483),
.B(n_2255),
.Y(n_2564)
);

INVx6_ASAP7_75t_SL g2565 ( 
.A(n_2477),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2292),
.A2(n_2211),
.B(n_2168),
.Y(n_2566)
);

CKINVDCx20_ASAP7_75t_R g2567 ( 
.A(n_2360),
.Y(n_2567)
);

A2O1A1Ixp33_ASAP7_75t_L g2568 ( 
.A1(n_2320),
.A2(n_2126),
.B(n_2155),
.C(n_2059),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2305),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2461),
.B(n_2135),
.Y(n_2570)
);

BUFx12f_ASAP7_75t_L g2571 ( 
.A(n_2270),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2317),
.A2(n_2330),
.B1(n_2379),
.B2(n_2400),
.Y(n_2572)
);

INVx3_ASAP7_75t_SL g2573 ( 
.A(n_2384),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2302),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2281),
.A2(n_2216),
.B(n_2196),
.Y(n_2575)
);

BUFx6f_ASAP7_75t_L g2576 ( 
.A(n_2270),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2306),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2285),
.B(n_2135),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2324),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2277),
.B(n_2137),
.Y(n_2580)
);

BUFx6f_ASAP7_75t_L g2581 ( 
.A(n_2332),
.Y(n_2581)
);

AOI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2261),
.A2(n_2266),
.B1(n_2525),
.B2(n_2515),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2313),
.Y(n_2583)
);

CKINVDCx5p33_ASAP7_75t_R g2584 ( 
.A(n_2344),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2325),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2340),
.Y(n_2586)
);

INVx4_ASAP7_75t_L g2587 ( 
.A(n_2340),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2295),
.B(n_2137),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2282),
.B(n_2172),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2287),
.B(n_2378),
.Y(n_2590)
);

OAI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2280),
.A2(n_2155),
.B1(n_2148),
.B2(n_2151),
.Y(n_2591)
);

OR2x6_ASAP7_75t_L g2592 ( 
.A(n_2275),
.B(n_2196),
.Y(n_2592)
);

AOI222xp33_ASAP7_75t_L g2593 ( 
.A1(n_2473),
.A2(n_821),
.B1(n_808),
.B2(n_674),
.C1(n_668),
.C2(n_675),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2303),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2311),
.Y(n_2595)
);

O2A1O1Ixp33_ASAP7_75t_L g2596 ( 
.A1(n_2498),
.A2(n_962),
.B(n_963),
.C(n_961),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2519),
.B(n_2140),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2346),
.Y(n_2598)
);

INVxp67_ASAP7_75t_L g2599 ( 
.A(n_2359),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2355),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2504),
.Y(n_2601)
);

NOR2x1_ASAP7_75t_L g2602 ( 
.A(n_2371),
.B(n_2033),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2409),
.B(n_2140),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2493),
.A2(n_2182),
.B(n_1605),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2357),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2269),
.Y(n_2606)
);

INVx2_ASAP7_75t_SL g2607 ( 
.A(n_2428),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2372),
.Y(n_2608)
);

INVx4_ASAP7_75t_L g2609 ( 
.A(n_2290),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2450),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2459),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2399),
.Y(n_2612)
);

BUFx3_ASAP7_75t_L g2613 ( 
.A(n_2458),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2504),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2407),
.Y(n_2615)
);

AOI21x1_ASAP7_75t_SL g2616 ( 
.A1(n_2314),
.A2(n_2032),
.B(n_1346),
.Y(n_2616)
);

OR2x2_ASAP7_75t_L g2617 ( 
.A(n_2369),
.B(n_2148),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2514),
.B(n_2397),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2414),
.B(n_2033),
.Y(n_2619)
);

CKINVDCx16_ASAP7_75t_R g2620 ( 
.A(n_2315),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2396),
.Y(n_2621)
);

OAI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2371),
.A2(n_2158),
.B1(n_2151),
.B2(n_2040),
.Y(n_2622)
);

OAI22xp5_ASAP7_75t_L g2623 ( 
.A1(n_2294),
.A2(n_2158),
.B1(n_2040),
.B2(n_2083),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2415),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2422),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2523),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2425),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2474),
.Y(n_2628)
);

INVx3_ASAP7_75t_L g2629 ( 
.A(n_2407),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2293),
.B(n_2059),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2386),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2488),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2291),
.B(n_2161),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2491),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2395),
.Y(n_2635)
);

BUFx2_ASAP7_75t_L g2636 ( 
.A(n_2441),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2414),
.B(n_2071),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2412),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2494),
.Y(n_2639)
);

INVx3_ASAP7_75t_L g2640 ( 
.A(n_2410),
.Y(n_2640)
);

AND2x6_ASAP7_75t_L g2641 ( 
.A(n_2271),
.B(n_2039),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2290),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2410),
.Y(n_2643)
);

INVx2_ASAP7_75t_SL g2644 ( 
.A(n_2368),
.Y(n_2644)
);

AOI221x1_ASAP7_75t_L g2645 ( 
.A1(n_2361),
.A2(n_2180),
.B1(n_2161),
.B2(n_2188),
.C(n_2083),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2426),
.B(n_2180),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2481),
.Y(n_2647)
);

AOI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2334),
.A2(n_2162),
.B1(n_670),
.B2(n_679),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2446),
.Y(n_2649)
);

OAI21xp5_ASAP7_75t_L g2650 ( 
.A1(n_2264),
.A2(n_2162),
.B(n_2188),
.Y(n_2650)
);

INVx3_ASAP7_75t_L g2651 ( 
.A(n_2481),
.Y(n_2651)
);

INVx2_ASAP7_75t_SL g2652 ( 
.A(n_2290),
.Y(n_2652)
);

HB1xp67_ASAP7_75t_L g2653 ( 
.A(n_2500),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2451),
.Y(n_2654)
);

HB1xp67_ASAP7_75t_L g2655 ( 
.A(n_2345),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2470),
.Y(n_2656)
);

CKINVDCx6p67_ASAP7_75t_R g2657 ( 
.A(n_2468),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2502),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_2298),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2435),
.B(n_2071),
.Y(n_2660)
);

OR2x6_ASAP7_75t_L g2661 ( 
.A(n_2416),
.B(n_2438),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2430),
.B(n_2096),
.Y(n_2662)
);

BUFx2_ASAP7_75t_L g2663 ( 
.A(n_2298),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2505),
.Y(n_2664)
);

INVx5_ASAP7_75t_L g2665 ( 
.A(n_2477),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2299),
.A2(n_2162),
.B1(n_683),
.B2(n_685),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2420),
.B(n_2096),
.Y(n_2667)
);

BUFx4_ASAP7_75t_SL g2668 ( 
.A(n_2477),
.Y(n_2668)
);

INVx2_ASAP7_75t_SL g2669 ( 
.A(n_2298),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2333),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2394),
.A2(n_2162),
.B1(n_687),
.B2(n_688),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2500),
.B(n_2162),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2420),
.B(n_2103),
.Y(n_2673)
);

AOI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_2424),
.A2(n_581),
.B1(n_540),
.B2(n_649),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2336),
.A2(n_2182),
.B(n_1605),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2310),
.B(n_2103),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2476),
.Y(n_2677)
);

CKINVDCx6p67_ASAP7_75t_R g2678 ( 
.A(n_2333),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2424),
.B(n_2115),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2501),
.Y(n_2680)
);

BUFx12f_ASAP7_75t_L g2681 ( 
.A(n_2333),
.Y(n_2681)
);

A2O1A1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_2487),
.A2(n_2115),
.B(n_2083),
.C(n_2040),
.Y(n_2682)
);

BUFx2_ASAP7_75t_L g2683 ( 
.A(n_2327),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2508),
.Y(n_2684)
);

INVxp33_ASAP7_75t_L g2685 ( 
.A(n_2419),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2286),
.B(n_2040),
.Y(n_2686)
);

BUFx2_ASAP7_75t_L g2687 ( 
.A(n_2327),
.Y(n_2687)
);

INVx5_ASAP7_75t_L g2688 ( 
.A(n_2296),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2510),
.Y(n_2689)
);

BUFx6f_ASAP7_75t_L g2690 ( 
.A(n_2471),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2286),
.B(n_2321),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2522),
.Y(n_2692)
);

AOI22xp33_ASAP7_75t_L g2693 ( 
.A1(n_2465),
.A2(n_2492),
.B1(n_2496),
.B2(n_2354),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_SL g2694 ( 
.A(n_2471),
.Y(n_2694)
);

INVx5_ASAP7_75t_L g2695 ( 
.A(n_2296),
.Y(n_2695)
);

AOI21xp5_ASAP7_75t_L g2696 ( 
.A1(n_2478),
.A2(n_2083),
.B(n_1338),
.Y(n_2696)
);

BUFx6f_ASAP7_75t_L g2697 ( 
.A(n_2472),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2480),
.Y(n_2698)
);

INVx4_ASAP7_75t_L g2699 ( 
.A(n_2472),
.Y(n_2699)
);

AOI22xp33_ASAP7_75t_SL g2700 ( 
.A1(n_2486),
.A2(n_698),
.B1(n_699),
.B2(n_692),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2376),
.Y(n_2701)
);

INVx4_ASAP7_75t_L g2702 ( 
.A(n_2376),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2391),
.B(n_2524),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_2337),
.B(n_962),
.Y(n_2704)
);

OAI21x1_ASAP7_75t_SL g2705 ( 
.A1(n_2444),
.A2(n_1533),
.B(n_1525),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2480),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_SL g2707 ( 
.A1(n_2398),
.A2(n_702),
.B1(n_705),
.B2(n_700),
.Y(n_2707)
);

CKINVDCx5p33_ASAP7_75t_R g2708 ( 
.A(n_2433),
.Y(n_2708)
);

INVx8_ASAP7_75t_L g2709 ( 
.A(n_2511),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2431),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2489),
.B(n_540),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2321),
.B(n_2032),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2374),
.A2(n_581),
.B1(n_711),
.B2(n_709),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2404),
.A2(n_2413),
.B1(n_2455),
.B2(n_2328),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2382),
.A2(n_712),
.B1(n_717),
.B2(n_715),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_SL g2716 ( 
.A(n_2381),
.B(n_2393),
.Y(n_2716)
);

OAI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2486),
.A2(n_721),
.B1(n_724),
.B2(n_719),
.Y(n_2717)
);

AOI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2401),
.A2(n_725),
.B1(n_732),
.B2(n_728),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_2391),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2503),
.Y(n_2720)
);

BUFx2_ASAP7_75t_L g2721 ( 
.A(n_2524),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2296),
.B(n_581),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_SL g2723 ( 
.A(n_2318),
.B(n_2032),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2342),
.B(n_1683),
.Y(n_2724)
);

BUFx3_ASAP7_75t_L g2725 ( 
.A(n_2467),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2464),
.B(n_2469),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2284),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2503),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2520),
.B(n_1805),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2392),
.B(n_2032),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2511),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2506),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2506),
.Y(n_2733)
);

BUFx3_ASAP7_75t_L g2734 ( 
.A(n_2467),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2499),
.A2(n_581),
.B1(n_739),
.B2(n_738),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2509),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2392),
.B(n_2032),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2329),
.A2(n_1555),
.B(n_1554),
.Y(n_2738)
);

AOI21xp33_ASAP7_75t_L g2739 ( 
.A1(n_2460),
.A2(n_1535),
.B(n_1534),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2343),
.Y(n_2740)
);

OAI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2262),
.A2(n_742),
.B1(n_743),
.B2(n_741),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2509),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2343),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2418),
.B(n_2032),
.Y(n_2744)
);

CKINVDCx20_ASAP7_75t_R g2745 ( 
.A(n_2364),
.Y(n_2745)
);

INVx6_ASAP7_75t_L g2746 ( 
.A(n_2326),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2512),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_SL g2748 ( 
.A(n_2411),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2512),
.Y(n_2749)
);

INVx4_ASAP7_75t_L g2750 ( 
.A(n_2284),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2429),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_SL g2752 ( 
.A(n_2381),
.B(n_581),
.Y(n_2752)
);

INVx3_ASAP7_75t_L g2753 ( 
.A(n_2278),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_2383),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2358),
.B(n_2322),
.Y(n_2755)
);

NAND2x1p5_ASAP7_75t_L g2756 ( 
.A(n_2380),
.B(n_1554),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2427),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_2383),
.Y(n_2758)
);

INVx3_ASAP7_75t_L g2759 ( 
.A(n_2278),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2323),
.A2(n_2338),
.B(n_2479),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2385),
.B(n_963),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_2499),
.A2(n_2352),
.B1(n_2288),
.B2(n_2362),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2427),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_2349),
.Y(n_2764)
);

CKINVDCx20_ASAP7_75t_R g2765 ( 
.A(n_2490),
.Y(n_2765)
);

O2A1O1Ixp33_ASAP7_75t_L g2766 ( 
.A1(n_2423),
.A2(n_965),
.B(n_966),
.C(n_964),
.Y(n_2766)
);

BUFx12f_ASAP7_75t_L g2767 ( 
.A(n_2442),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2385),
.Y(n_2768)
);

BUFx6f_ASAP7_75t_L g2769 ( 
.A(n_2406),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2418),
.B(n_1534),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2337),
.B(n_1535),
.Y(n_2771)
);

CKINVDCx14_ASAP7_75t_R g2772 ( 
.A(n_2393),
.Y(n_2772)
);

BUFx12f_ASAP7_75t_L g2773 ( 
.A(n_2272),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2436),
.A2(n_746),
.B1(n_749),
.B2(n_744),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2363),
.Y(n_2775)
);

INVx4_ASAP7_75t_L g2776 ( 
.A(n_2339),
.Y(n_2776)
);

BUFx6f_ASAP7_75t_L g2777 ( 
.A(n_2421),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2363),
.Y(n_2778)
);

NAND2xp33_ASAP7_75t_L g2779 ( 
.A(n_2331),
.B(n_752),
.Y(n_2779)
);

INVxp67_ASAP7_75t_L g2780 ( 
.A(n_2362),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2366),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2497),
.B(n_1805),
.Y(n_2782)
);

BUFx3_ASAP7_75t_L g2783 ( 
.A(n_2437),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2436),
.A2(n_755),
.B1(n_756),
.B2(n_754),
.Y(n_2784)
);

BUFx4f_ASAP7_75t_SL g2785 ( 
.A(n_2432),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2417),
.Y(n_2786)
);

NAND2x1p5_ASAP7_75t_L g2787 ( 
.A(n_2602),
.B(n_2454),
.Y(n_2787)
);

AOI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2779),
.A2(n_2479),
.B(n_2370),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2540),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_L g2790 ( 
.A(n_2581),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_2581),
.Y(n_2791)
);

AND2x4_ASAP7_75t_L g2792 ( 
.A(n_2655),
.B(n_2402),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2557),
.Y(n_2793)
);

OAI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2582),
.A2(n_2448),
.B1(n_2341),
.B2(n_2339),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2552),
.Y(n_2795)
);

OAI21x1_ASAP7_75t_L g2796 ( 
.A1(n_2738),
.A2(n_2389),
.B(n_2353),
.Y(n_2796)
);

INVxp67_ASAP7_75t_L g2797 ( 
.A(n_2610),
.Y(n_2797)
);

A2O1A1Ixp33_ASAP7_75t_L g2798 ( 
.A1(n_2693),
.A2(n_2445),
.B(n_2456),
.C(n_2447),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2558),
.B(n_2434),
.Y(n_2799)
);

INVx1_ASAP7_75t_SL g2800 ( 
.A(n_2611),
.Y(n_2800)
);

OAI21x1_ASAP7_75t_L g2801 ( 
.A1(n_2738),
.A2(n_2319),
.B(n_2377),
.Y(n_2801)
);

O2A1O1Ixp33_ASAP7_75t_SL g2802 ( 
.A1(n_2536),
.A2(n_2341),
.B(n_2408),
.C(n_2516),
.Y(n_2802)
);

AO32x2_ASAP7_75t_L g2803 ( 
.A1(n_2591),
.A2(n_2417),
.A3(n_2463),
.B1(n_2457),
.B2(n_2403),
.Y(n_2803)
);

OAI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_2765),
.A2(n_2518),
.B1(n_2453),
.B2(n_2475),
.Y(n_2804)
);

OAI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2593),
.A2(n_2741),
.B(n_2714),
.Y(n_2805)
);

NAND2xp33_ASAP7_75t_SL g2806 ( 
.A(n_2748),
.B(n_2532),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2572),
.A2(n_2484),
.B1(n_2449),
.B2(n_2440),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2616),
.A2(n_2521),
.B(n_2350),
.Y(n_2808)
);

NOR2x1_ASAP7_75t_SL g2809 ( 
.A(n_2533),
.B(n_2417),
.Y(n_2809)
);

AOI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2760),
.A2(n_2390),
.B(n_2405),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2581),
.Y(n_2811)
);

AOI221xp5_ASAP7_75t_L g2812 ( 
.A1(n_2741),
.A2(n_764),
.B1(n_766),
.B2(n_763),
.C(n_762),
.Y(n_2812)
);

HB1xp67_ASAP7_75t_L g2813 ( 
.A(n_2612),
.Y(n_2813)
);

A2O1A1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2774),
.A2(n_2351),
.B(n_2367),
.C(n_2443),
.Y(n_2814)
);

OAI21x1_ASAP7_75t_L g2815 ( 
.A1(n_2616),
.A2(n_2521),
.B(n_2495),
.Y(n_2815)
);

O2A1O1Ixp33_ASAP7_75t_L g2816 ( 
.A1(n_2593),
.A2(n_2403),
.B(n_965),
.C(n_966),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2760),
.A2(n_1555),
.B(n_1554),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2531),
.B(n_964),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2633),
.B(n_967),
.Y(n_2819)
);

OAI21x1_ASAP7_75t_L g2820 ( 
.A1(n_2575),
.A2(n_1553),
.B(n_1531),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2574),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2561),
.B(n_967),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2660),
.B(n_968),
.Y(n_2823)
);

OAI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2575),
.A2(n_1540),
.B(n_1538),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2773),
.A2(n_772),
.B1(n_773),
.B2(n_771),
.Y(n_2825)
);

AO31x2_ASAP7_75t_L g2826 ( 
.A1(n_2750),
.A2(n_1538),
.A3(n_1543),
.B(n_1540),
.Y(n_2826)
);

O2A1O1Ixp33_ASAP7_75t_L g2827 ( 
.A1(n_2568),
.A2(n_970),
.B(n_971),
.C(n_968),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2577),
.Y(n_2828)
);

OAI21x1_ASAP7_75t_L g2829 ( 
.A1(n_2539),
.A2(n_1546),
.B(n_1543),
.Y(n_2829)
);

OAI22xp33_ASAP7_75t_L g2830 ( 
.A1(n_2767),
.A2(n_777),
.B1(n_783),
.B2(n_775),
.Y(n_2830)
);

OAI222xp33_ASAP7_75t_L g2831 ( 
.A1(n_2546),
.A2(n_796),
.B1(n_791),
.B2(n_798),
.C1(n_792),
.C2(n_790),
.Y(n_2831)
);

OR2x2_ASAP7_75t_L g2832 ( 
.A(n_2612),
.B(n_970),
.Y(n_2832)
);

INVxp67_ASAP7_75t_SL g2833 ( 
.A(n_2579),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2533),
.A2(n_1555),
.B(n_1805),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2535),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2583),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2533),
.A2(n_1555),
.B(n_1546),
.Y(n_2837)
);

AO31x2_ASAP7_75t_L g2838 ( 
.A1(n_2750),
.A2(n_1322),
.A3(n_1262),
.B(n_1267),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2564),
.B(n_971),
.Y(n_2839)
);

AO32x2_ASAP7_75t_L g2840 ( 
.A1(n_2591),
.A2(n_2546),
.A3(n_2622),
.B1(n_2623),
.B2(n_2530),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2780),
.B(n_2),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2748),
.A2(n_806),
.B1(n_807),
.B2(n_802),
.Y(n_2842)
);

INVx3_ASAP7_75t_SL g2843 ( 
.A(n_2573),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2555),
.Y(n_2844)
);

OA21x2_ASAP7_75t_L g2845 ( 
.A1(n_2645),
.A2(n_1246),
.B(n_1245),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2685),
.B(n_810),
.Y(n_2846)
);

INVx5_ASAP7_75t_L g2847 ( 
.A(n_2661),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2585),
.Y(n_2848)
);

O2A1O1Ixp33_ASAP7_75t_L g2849 ( 
.A1(n_2717),
.A2(n_1254),
.B(n_813),
.C(n_815),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2541),
.Y(n_2850)
);

OAI222xp33_ASAP7_75t_L g2851 ( 
.A1(n_2700),
.A2(n_816),
.B1(n_818),
.B2(n_811),
.C1(n_6),
.C2(n_8),
.Y(n_2851)
);

AOI21x1_ASAP7_75t_L g2852 ( 
.A1(n_2579),
.A2(n_1155),
.B(n_1143),
.Y(n_2852)
);

NAND2xp33_ASAP7_75t_L g2853 ( 
.A(n_2708),
.B(n_835),
.Y(n_2853)
);

INVxp67_ASAP7_75t_L g2854 ( 
.A(n_2607),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2675),
.A2(n_1555),
.B(n_1265),
.Y(n_2855)
);

INVx4_ASAP7_75t_L g2856 ( 
.A(n_2555),
.Y(n_2856)
);

O2A1O1Ixp33_ASAP7_75t_L g2857 ( 
.A1(n_2717),
.A2(n_1156),
.B(n_1158),
.C(n_1155),
.Y(n_2857)
);

O2A1O1Ixp33_ASAP7_75t_SL g2858 ( 
.A1(n_2682),
.A2(n_6),
.B(n_3),
.C(n_5),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2590),
.B(n_7),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2539),
.A2(n_1322),
.B(n_1265),
.Y(n_2860)
);

OR2x6_ASAP7_75t_L g2861 ( 
.A(n_2709),
.B(n_1156),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2598),
.Y(n_2862)
);

AOI221xp5_ASAP7_75t_L g2863 ( 
.A1(n_2707),
.A2(n_1178),
.B1(n_1192),
.B2(n_1162),
.C(n_1158),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2600),
.Y(n_2864)
);

AO31x2_ASAP7_75t_L g2865 ( 
.A1(n_2786),
.A2(n_1267),
.A3(n_1262),
.B(n_1178),
.Y(n_2865)
);

OAI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2666),
.A2(n_1192),
.B(n_1162),
.Y(n_2866)
);

CKINVDCx9p33_ASAP7_75t_R g2867 ( 
.A(n_2636),
.Y(n_2867)
);

A2O1A1Ixp33_ASAP7_75t_L g2868 ( 
.A1(n_2700),
.A2(n_2671),
.B(n_2547),
.C(n_2772),
.Y(n_2868)
);

CKINVDCx6p67_ASAP7_75t_R g2869 ( 
.A(n_2560),
.Y(n_2869)
);

INVxp67_ASAP7_75t_SL g2870 ( 
.A(n_2649),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2675),
.A2(n_1305),
.B(n_1288),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2558),
.B(n_7),
.Y(n_2872)
);

AOI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2641),
.A2(n_1209),
.B1(n_1221),
.B2(n_1197),
.Y(n_2873)
);

OAI22xp33_ASAP7_75t_L g2874 ( 
.A1(n_2716),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2745),
.A2(n_1209),
.B1(n_1221),
.B2(n_1197),
.Y(n_2875)
);

NOR2xp67_ASAP7_75t_L g2876 ( 
.A(n_2542),
.B(n_10),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2605),
.Y(n_2877)
);

OR2x2_ASAP7_75t_L g2878 ( 
.A(n_2780),
.B(n_12),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2604),
.A2(n_2592),
.B(n_2782),
.Y(n_2879)
);

OAI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2547),
.A2(n_1227),
.B(n_1226),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2604),
.A2(n_1508),
.B(n_1227),
.Y(n_2881)
);

OAI21x1_ASAP7_75t_L g2882 ( 
.A1(n_2563),
.A2(n_1234),
.B(n_1226),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2691),
.B(n_13),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2589),
.B(n_13),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2584),
.B(n_14),
.Y(n_2885)
);

O2A1O1Ixp33_ASAP7_75t_SL g2886 ( 
.A1(n_2630),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_2886)
);

O2A1O1Ixp33_ASAP7_75t_SL g2887 ( 
.A1(n_2549),
.A2(n_20),
.B(n_15),
.C(n_19),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2608),
.Y(n_2888)
);

O2A1O1Ixp33_ASAP7_75t_L g2889 ( 
.A1(n_2530),
.A2(n_1235),
.B(n_1234),
.C(n_1123),
.Y(n_2889)
);

NOR2xp67_ASAP7_75t_L g2890 ( 
.A(n_2542),
.B(n_2599),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2592),
.A2(n_1508),
.B(n_1235),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2631),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2688),
.B(n_366),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2592),
.A2(n_1508),
.B(n_1169),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2752),
.A2(n_1169),
.B(n_1168),
.Y(n_2895)
);

CKINVDCx11_ASAP7_75t_R g2896 ( 
.A(n_2567),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2752),
.A2(n_1169),
.B(n_1168),
.Y(n_2897)
);

AO31x2_ASAP7_75t_L g2898 ( 
.A1(n_2623),
.A2(n_1251),
.A3(n_1257),
.B(n_1247),
.Y(n_2898)
);

OAI22x1_ASAP7_75t_L g2899 ( 
.A1(n_2599),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_2899)
);

O2A1O1Ixp33_ASAP7_75t_SL g2900 ( 
.A1(n_2691),
.A2(n_26),
.B(n_23),
.C(n_24),
.Y(n_2900)
);

O2A1O1Ixp33_ASAP7_75t_SL g2901 ( 
.A1(n_2686),
.A2(n_27),
.B(n_23),
.C(n_26),
.Y(n_2901)
);

BUFx3_ASAP7_75t_L g2902 ( 
.A(n_2535),
.Y(n_2902)
);

O2A1O1Ixp33_ASAP7_75t_SL g2903 ( 
.A1(n_2686),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2903)
);

BUFx3_ASAP7_75t_L g2904 ( 
.A(n_2571),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2566),
.A2(n_1169),
.B(n_1168),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2635),
.Y(n_2906)
);

O2A1O1Ixp33_ASAP7_75t_L g2907 ( 
.A1(n_2534),
.A2(n_1123),
.B(n_1138),
.C(n_1105),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2710),
.B(n_29),
.Y(n_2908)
);

O2A1O1Ixp33_ASAP7_75t_SL g2909 ( 
.A1(n_2545),
.A2(n_33),
.B(n_30),
.C(n_32),
.Y(n_2909)
);

INVx5_ASAP7_75t_L g2910 ( 
.A(n_2661),
.Y(n_2910)
);

O2A1O1Ixp33_ASAP7_75t_L g2911 ( 
.A1(n_2534),
.A2(n_1123),
.B(n_1138),
.C(n_1105),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2566),
.A2(n_1194),
.B(n_1169),
.Y(n_2912)
);

O2A1O1Ixp33_ASAP7_75t_SL g2913 ( 
.A1(n_2545),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_2913)
);

AO31x2_ASAP7_75t_L g2914 ( 
.A1(n_2622),
.A2(n_1251),
.A3(n_1257),
.B(n_1247),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2638),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2552),
.Y(n_2916)
);

BUFx3_ASAP7_75t_L g2917 ( 
.A(n_2544),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2654),
.Y(n_2918)
);

INVx1_ASAP7_75t_SL g2919 ( 
.A(n_2746),
.Y(n_2919)
);

OAI21x1_ASAP7_75t_L g2920 ( 
.A1(n_2563),
.A2(n_1138),
.B(n_1105),
.Y(n_2920)
);

OR2x2_ASAP7_75t_L g2921 ( 
.A(n_2775),
.B(n_2778),
.Y(n_2921)
);

OAI21x1_ASAP7_75t_L g2922 ( 
.A1(n_2705),
.A2(n_1150),
.B(n_1146),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2537),
.B(n_34),
.Y(n_2923)
);

OAI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2711),
.A2(n_1269),
.B(n_1264),
.Y(n_2924)
);

AOI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2716),
.A2(n_1449),
.B1(n_1150),
.B2(n_1195),
.Y(n_2925)
);

OAI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2715),
.A2(n_2718),
.B(n_2553),
.Y(n_2926)
);

O2A1O1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_2644),
.A2(n_1150),
.B(n_1195),
.C(n_1146),
.Y(n_2927)
);

A2O1A1Ixp33_ASAP7_75t_L g2928 ( 
.A1(n_2648),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2688),
.B(n_367),
.Y(n_2929)
);

OAI211xp5_ASAP7_75t_L g2930 ( 
.A1(n_2784),
.A2(n_43),
.B(n_39),
.C(n_41),
.Y(n_2930)
);

O2A1O1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2650),
.A2(n_1195),
.B(n_1225),
.C(n_1146),
.Y(n_2931)
);

BUFx12f_ASAP7_75t_L g2932 ( 
.A(n_2594),
.Y(n_2932)
);

OA21x2_ASAP7_75t_L g2933 ( 
.A1(n_2727),
.A2(n_1269),
.B(n_1264),
.Y(n_2933)
);

OAI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2735),
.A2(n_1282),
.B(n_1270),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2555),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2538),
.B(n_43),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2562),
.Y(n_2937)
);

O2A1O1Ixp33_ASAP7_75t_SL g2938 ( 
.A1(n_2726),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2543),
.A2(n_1449),
.B1(n_1232),
.B2(n_1268),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2650),
.A2(n_1202),
.B(n_1194),
.Y(n_2940)
);

AOI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2641),
.A2(n_1449),
.B1(n_1232),
.B2(n_1268),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2692),
.Y(n_2942)
);

OAI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2762),
.A2(n_1282),
.B(n_1270),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2641),
.A2(n_1449),
.B1(n_1232),
.B2(n_1268),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2656),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2713),
.A2(n_1289),
.B(n_1280),
.Y(n_2946)
);

OR2x6_ASAP7_75t_L g2947 ( 
.A(n_2709),
.B(n_1010),
.Y(n_2947)
);

OAI21x1_ASAP7_75t_SL g2948 ( 
.A1(n_2776),
.A2(n_44),
.B(n_45),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_2746),
.B(n_46),
.Y(n_2949)
);

OA21x2_ASAP7_75t_L g2950 ( 
.A1(n_2727),
.A2(n_1289),
.B(n_47),
.Y(n_2950)
);

A2O1A1Ixp33_ASAP7_75t_L g2951 ( 
.A1(n_2674),
.A2(n_52),
.B(n_49),
.C(n_51),
.Y(n_2951)
);

OAI21x1_ASAP7_75t_L g2952 ( 
.A1(n_2753),
.A2(n_1280),
.B(n_1225),
.Y(n_2952)
);

AO32x2_ASAP7_75t_L g2953 ( 
.A1(n_2776),
.A2(n_55),
.A3(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2764),
.A2(n_1280),
.B1(n_1293),
.B2(n_1225),
.Y(n_2954)
);

CKINVDCx5p33_ASAP7_75t_R g2955 ( 
.A(n_2657),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2538),
.B(n_55),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2696),
.A2(n_1202),
.B(n_1194),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2722),
.A2(n_1316),
.B(n_1293),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2641),
.A2(n_1316),
.B1(n_1293),
.B2(n_1010),
.Y(n_2959)
);

AND2x4_ASAP7_75t_L g2960 ( 
.A(n_2688),
.B(n_370),
.Y(n_2960)
);

AND2x6_ASAP7_75t_L g2961 ( 
.A(n_2672),
.B(n_2724),
.Y(n_2961)
);

OAI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2620),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2783),
.B(n_60),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2677),
.Y(n_2964)
);

OAI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2746),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2576),
.Y(n_2966)
);

A2O1A1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2596),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2556),
.A2(n_1316),
.B1(n_1010),
.B2(n_1014),
.Y(n_2968)
);

O2A1O1Ixp33_ASAP7_75t_SL g2969 ( 
.A1(n_2726),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2680),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_SL g2971 ( 
.A1(n_2672),
.A2(n_67),
.B(n_68),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2769),
.Y(n_2972)
);

AOI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2679),
.A2(n_1010),
.B1(n_1014),
.B2(n_1011),
.Y(n_2973)
);

OAI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2696),
.A2(n_372),
.B(n_371),
.Y(n_2974)
);

BUFx2_ASAP7_75t_L g2975 ( 
.A(n_2526),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_L g2976 ( 
.A1(n_2761),
.A2(n_1011),
.B1(n_1014),
.B2(n_1010),
.Y(n_2976)
);

AOI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_2723),
.A2(n_1202),
.B(n_1194),
.Y(n_2977)
);

A2O1A1Ixp33_ASAP7_75t_L g2978 ( 
.A1(n_2596),
.A2(n_2766),
.B(n_2606),
.C(n_2695),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2597),
.B(n_67),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2684),
.Y(n_2980)
);

OAI21xp5_ASAP7_75t_L g2981 ( 
.A1(n_2704),
.A2(n_374),
.B(n_373),
.Y(n_2981)
);

NOR2xp67_ASAP7_75t_L g2982 ( 
.A(n_2527),
.B(n_2688),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2529),
.Y(n_2983)
);

OAI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2766),
.A2(n_378),
.B(n_377),
.Y(n_2984)
);

OAI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2570),
.A2(n_2676),
.B(n_2597),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2578),
.B(n_69),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2554),
.Y(n_2987)
);

OAI21x1_ASAP7_75t_L g2988 ( 
.A1(n_2753),
.A2(n_380),
.B(n_379),
.Y(n_2988)
);

OAI21x1_ASAP7_75t_L g2989 ( 
.A1(n_2759),
.A2(n_383),
.B(n_382),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2653),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2569),
.Y(n_2991)
);

OAI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2785),
.A2(n_1202),
.B1(n_1206),
.B2(n_1194),
.Y(n_2992)
);

AOI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2537),
.A2(n_1011),
.B1(n_1022),
.B2(n_1014),
.Y(n_2993)
);

AO31x2_ASAP7_75t_L g2994 ( 
.A1(n_2712),
.A2(n_1053),
.A3(n_1016),
.B(n_71),
.Y(n_2994)
);

A2O1A1Ixp33_ASAP7_75t_L g2995 ( 
.A1(n_2695),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2578),
.B(n_2755),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2653),
.Y(n_2997)
);

AOI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_2661),
.A2(n_1206),
.B(n_1202),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2595),
.Y(n_2999)
);

AOI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2662),
.A2(n_1011),
.B1(n_1022),
.B2(n_1014),
.Y(n_3000)
);

O2A1O1Ixp33_ASAP7_75t_L g3001 ( 
.A1(n_2712),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2559),
.A2(n_1230),
.B(n_1206),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2551),
.B(n_74),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2621),
.Y(n_3004)
);

O2A1O1Ixp33_ASAP7_75t_L g3005 ( 
.A1(n_2781),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_3005)
);

O2A1O1Ixp33_ASAP7_75t_SL g3006 ( 
.A1(n_2551),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2624),
.Y(n_3007)
);

OAI21x1_ASAP7_75t_L g3008 ( 
.A1(n_2759),
.A2(n_2751),
.B(n_2771),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2559),
.A2(n_1230),
.B(n_1206),
.Y(n_3009)
);

INVx5_ASAP7_75t_L g3010 ( 
.A(n_2576),
.Y(n_3010)
);

O2A1O1Ixp33_ASAP7_75t_SL g3011 ( 
.A1(n_2831),
.A2(n_2652),
.B(n_2669),
.C(n_2617),
.Y(n_3011)
);

CKINVDCx6p67_ASAP7_75t_R g3012 ( 
.A(n_2843),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2896),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2821),
.Y(n_3014)
);

INVx6_ASAP7_75t_L g3015 ( 
.A(n_2790),
.Y(n_3015)
);

BUFx2_ASAP7_75t_L g3016 ( 
.A(n_2795),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2805),
.A2(n_2548),
.B1(n_2665),
.B2(n_2695),
.Y(n_3017)
);

INVx4_ASAP7_75t_L g3018 ( 
.A(n_3010),
.Y(n_3018)
);

AOI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2926),
.A2(n_2758),
.B1(n_2768),
.B2(n_2754),
.Y(n_3019)
);

OAI21xp5_ASAP7_75t_L g3020 ( 
.A1(n_2974),
.A2(n_2771),
.B(n_2580),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2789),
.Y(n_3021)
);

INVx2_ASAP7_75t_SL g3022 ( 
.A(n_2790),
.Y(n_3022)
);

INVx3_ASAP7_75t_L g3023 ( 
.A(n_2795),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2828),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2848),
.Y(n_3025)
);

AOI221xp5_ASAP7_75t_L g3026 ( 
.A1(n_2851),
.A2(n_2603),
.B1(n_2646),
.B2(n_2618),
.C(n_2550),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2984),
.A2(n_2734),
.B1(n_2725),
.B2(n_2695),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_2850),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2800),
.B(n_2576),
.Y(n_3029)
);

BUFx4_ASAP7_75t_R g3030 ( 
.A(n_2835),
.Y(n_3030)
);

AOI22xp33_ASAP7_75t_L g3031 ( 
.A1(n_2859),
.A2(n_2618),
.B1(n_2588),
.B2(n_2694),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2868),
.A2(n_2665),
.B1(n_2580),
.B2(n_2757),
.Y(n_3032)
);

OR2x6_ASAP7_75t_L g3033 ( 
.A(n_2879),
.B(n_2730),
.Y(n_3033)
);

AO21x2_ASAP7_75t_L g3034 ( 
.A1(n_2998),
.A2(n_2737),
.B(n_2730),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2793),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_2874),
.A2(n_2665),
.B1(n_2763),
.B2(n_2565),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2804),
.A2(n_2694),
.B1(n_2777),
.B2(n_2769),
.Y(n_3037)
);

NAND3x1_ASAP7_75t_L g3038 ( 
.A(n_2885),
.B(n_2601),
.C(n_2528),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_L g3039 ( 
.A(n_2790),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2862),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2836),
.Y(n_3041)
);

AOI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_2962),
.A2(n_2777),
.B1(n_2769),
.B2(n_2724),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2847),
.B(n_2777),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2892),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2864),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2830),
.A2(n_2613),
.B1(n_2729),
.B2(n_2637),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2877),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_L g3048 ( 
.A1(n_2825),
.A2(n_2729),
.B1(n_2619),
.B2(n_2667),
.Y(n_3048)
);

O2A1O1Ixp33_ASAP7_75t_L g3049 ( 
.A1(n_2995),
.A2(n_2701),
.B(n_2740),
.C(n_2756),
.Y(n_3049)
);

O2A1O1Ixp5_ASAP7_75t_L g3050 ( 
.A1(n_2930),
.A2(n_2615),
.B(n_2640),
.C(n_2629),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2971),
.A2(n_2619),
.B1(n_2667),
.B2(n_2637),
.Y(n_3051)
);

OR2x2_ASAP7_75t_L g3052 ( 
.A(n_2813),
.B(n_2737),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2996),
.B(n_2744),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_2869),
.Y(n_3054)
);

XNOR2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2955),
.B(n_2975),
.Y(n_3055)
);

BUFx10_ASAP7_75t_L g3056 ( 
.A(n_2846),
.Y(n_3056)
);

O2A1O1Ixp33_ASAP7_75t_SL g3057 ( 
.A1(n_2965),
.A2(n_2967),
.B(n_2798),
.C(n_2951),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2888),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_SL g3059 ( 
.A1(n_2981),
.A2(n_2665),
.B1(n_2587),
.B2(n_2709),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2906),
.Y(n_3060)
);

AOI221xp5_ASAP7_75t_L g3061 ( 
.A1(n_3001),
.A2(n_2720),
.B1(n_2728),
.B2(n_2706),
.C(n_2698),
.Y(n_3061)
);

OAI22xp5_ASAP7_75t_L g3062 ( 
.A1(n_2928),
.A2(n_2565),
.B1(n_2744),
.B2(n_2736),
.Y(n_3062)
);

O2A1O1Ixp33_ASAP7_75t_L g3063 ( 
.A1(n_2858),
.A2(n_2701),
.B(n_2740),
.C(n_2756),
.Y(n_3063)
);

NAND3xp33_ASAP7_75t_L g3064 ( 
.A(n_3005),
.B(n_2627),
.C(n_2625),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2937),
.B(n_2751),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2895),
.A2(n_2559),
.B(n_2739),
.Y(n_3066)
);

AOI221xp5_ASAP7_75t_L g3067 ( 
.A1(n_2909),
.A2(n_2747),
.B1(n_2742),
.B2(n_2733),
.C(n_2632),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2915),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2918),
.Y(n_3069)
);

AOI221xp5_ASAP7_75t_L g3070 ( 
.A1(n_2913),
.A2(n_2634),
.B1(n_2658),
.B2(n_2639),
.C(n_2628),
.Y(n_3070)
);

O2A1O1Ixp33_ASAP7_75t_SL g3071 ( 
.A1(n_2963),
.A2(n_2668),
.B(n_2601),
.C(n_2614),
.Y(n_3071)
);

AND2x4_ASAP7_75t_L g3072 ( 
.A(n_2916),
.B(n_2683),
.Y(n_3072)
);

OAI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_2919),
.A2(n_2587),
.B1(n_2699),
.B2(n_2626),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2797),
.B(n_2732),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2807),
.A2(n_2697),
.B1(n_2690),
.B2(n_2699),
.Y(n_3075)
);

INVx2_ASAP7_75t_SL g3076 ( 
.A(n_2791),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2964),
.Y(n_3077)
);

OAI221xp5_ASAP7_75t_L g3078 ( 
.A1(n_2812),
.A2(n_2629),
.B1(n_2643),
.B2(n_2640),
.C(n_2615),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2985),
.B(n_2749),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2970),
.Y(n_3080)
);

INVx2_ASAP7_75t_SL g3081 ( 
.A(n_2791),
.Y(n_3081)
);

AND2x6_ASAP7_75t_L g3082 ( 
.A(n_2893),
.B(n_2743),
.Y(n_3082)
);

AOI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_2806),
.A2(n_2673),
.B1(n_2703),
.B2(n_2731),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_2818),
.B(n_2731),
.Y(n_3084)
);

OAI22xp33_ASAP7_75t_L g3085 ( 
.A1(n_2959),
.A2(n_2731),
.B1(n_2697),
.B2(n_2690),
.Y(n_3085)
);

CKINVDCx20_ASAP7_75t_R g3086 ( 
.A(n_2867),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2980),
.Y(n_3087)
);

AOI22xp33_ASAP7_75t_SL g3088 ( 
.A1(n_2948),
.A2(n_2809),
.B1(n_2961),
.B2(n_2910),
.Y(n_3088)
);

CKINVDCx20_ASAP7_75t_R g3089 ( 
.A(n_2902),
.Y(n_3089)
);

INVx3_ASAP7_75t_L g3090 ( 
.A(n_2916),
.Y(n_3090)
);

OAI221xp5_ASAP7_75t_L g3091 ( 
.A1(n_2842),
.A2(n_2647),
.B1(n_2651),
.B2(n_2643),
.C(n_2687),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2870),
.B(n_2799),
.Y(n_3092)
);

NOR4xp25_ASAP7_75t_L g3093 ( 
.A(n_2900),
.B(n_2689),
.C(n_2664),
.D(n_2651),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2792),
.B(n_2721),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2945),
.Y(n_3095)
);

O2A1O1Ixp33_ASAP7_75t_SL g3096 ( 
.A1(n_2872),
.A2(n_2668),
.B(n_2614),
.C(n_2528),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2942),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_SL g3098 ( 
.A1(n_2961),
.A2(n_2743),
.B1(n_2586),
.B2(n_2697),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2917),
.B(n_2854),
.Y(n_3099)
);

AOI22xp33_ASAP7_75t_SL g3100 ( 
.A1(n_2961),
.A2(n_2743),
.B1(n_2586),
.B2(n_2690),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_SL g3101 ( 
.A1(n_2961),
.A2(n_2847),
.B1(n_2910),
.B2(n_2940),
.Y(n_3101)
);

OAI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_2899),
.A2(n_2586),
.B1(n_2702),
.B2(n_2719),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_3004),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2990),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_2817),
.A2(n_2770),
.B(n_2647),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2839),
.B(n_2703),
.Y(n_3106)
);

AOI22xp33_ASAP7_75t_L g3107 ( 
.A1(n_2792),
.A2(n_2673),
.B1(n_2719),
.B2(n_2702),
.Y(n_3107)
);

INVx4_ASAP7_75t_L g3108 ( 
.A(n_3010),
.Y(n_3108)
);

BUFx3_ASAP7_75t_L g3109 ( 
.A(n_2791),
.Y(n_3109)
);

OR2x6_ASAP7_75t_L g3110 ( 
.A(n_2810),
.B(n_2681),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3007),
.B(n_2663),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_2832),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2997),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_SL g3114 ( 
.A1(n_2847),
.A2(n_2719),
.B1(n_2642),
.B2(n_2670),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2983),
.Y(n_3115)
);

OAI21xp5_ASAP7_75t_SL g3116 ( 
.A1(n_2849),
.A2(n_2670),
.B(n_2642),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2833),
.Y(n_3117)
);

AOI22xp33_ASAP7_75t_SL g3118 ( 
.A1(n_2910),
.A2(n_2642),
.B1(n_2670),
.B2(n_2609),
.Y(n_3118)
);

OAI22xp5_ASAP7_75t_SL g3119 ( 
.A1(n_2949),
.A2(n_2609),
.B1(n_2659),
.B2(n_2770),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2921),
.Y(n_3120)
);

OAI22xp5_ASAP7_75t_SL g3121 ( 
.A1(n_2932),
.A2(n_83),
.B1(n_79),
.B2(n_82),
.Y(n_3121)
);

OAI221xp5_ASAP7_75t_L g3122 ( 
.A1(n_2853),
.A2(n_2739),
.B1(n_86),
.B2(n_84),
.C(n_85),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_2822),
.A2(n_2678),
.B1(n_1022),
.B2(n_1033),
.Y(n_3123)
);

INVx3_ASAP7_75t_SL g3124 ( 
.A(n_2811),
.Y(n_3124)
);

AND2x4_ASAP7_75t_L g3125 ( 
.A(n_2890),
.B(n_84),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2819),
.B(n_86),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2987),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_2811),
.Y(n_3128)
);

BUFx3_ASAP7_75t_L g3129 ( 
.A(n_2811),
.Y(n_3129)
);

AOI22xp33_ASAP7_75t_L g3130 ( 
.A1(n_2958),
.A2(n_1022),
.B1(n_1033),
.B2(n_1011),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2844),
.Y(n_3131)
);

OAI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_2925),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2972),
.B(n_87),
.Y(n_3133)
);

OR2x6_ASAP7_75t_L g3134 ( 
.A(n_2982),
.B(n_2881),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_2884),
.A2(n_1033),
.B1(n_1035),
.B2(n_1022),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2991),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_2904),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_2788),
.A2(n_1035),
.B1(n_1062),
.B2(n_1033),
.Y(n_3138)
);

O2A1O1Ixp33_ASAP7_75t_L g3139 ( 
.A1(n_2938),
.A2(n_92),
.B(n_88),
.C(n_91),
.Y(n_3139)
);

OAI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2883),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_3140)
);

CKINVDCx5p33_ASAP7_75t_R g3141 ( 
.A(n_2844),
.Y(n_3141)
);

BUFx10_ASAP7_75t_L g3142 ( 
.A(n_2893),
.Y(n_3142)
);

OR2x2_ASAP7_75t_L g3143 ( 
.A(n_3008),
.B(n_93),
.Y(n_3143)
);

NAND2xp33_ASAP7_75t_L g3144 ( 
.A(n_2978),
.B(n_1033),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2999),
.Y(n_3145)
);

AOI22xp33_ASAP7_75t_SL g3146 ( 
.A1(n_2929),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_2876),
.A2(n_1062),
.B1(n_1063),
.B2(n_1035),
.Y(n_3147)
);

OR2x6_ASAP7_75t_L g3148 ( 
.A(n_2834),
.B(n_2894),
.Y(n_3148)
);

AOI221xp5_ASAP7_75t_L g3149 ( 
.A1(n_2969),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.C(n_99),
.Y(n_3149)
);

AOI222xp33_ASAP7_75t_L g3150 ( 
.A1(n_2979),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.C1(n_103),
.C2(n_104),
.Y(n_3150)
);

AOI221xp5_ASAP7_75t_L g3151 ( 
.A1(n_2901),
.A2(n_106),
.B1(n_101),
.B2(n_105),
.C(n_107),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_2923),
.A2(n_1062),
.B1(n_1063),
.B2(n_1035),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2972),
.Y(n_3153)
);

BUFx2_ASAP7_75t_L g3154 ( 
.A(n_2856),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2865),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_2794),
.A2(n_1062),
.B1(n_1063),
.B2(n_1035),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2856),
.B(n_105),
.Y(n_3157)
);

AOI22xp33_ASAP7_75t_L g3158 ( 
.A1(n_2929),
.A2(n_1063),
.B1(n_1065),
.B2(n_1062),
.Y(n_3158)
);

CKINVDCx11_ASAP7_75t_R g3159 ( 
.A(n_2844),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2865),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2936),
.B(n_106),
.Y(n_3161)
);

BUFx2_ASAP7_75t_L g3162 ( 
.A(n_2935),
.Y(n_3162)
);

OAI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2941),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3163)
);

AOI222xp33_ASAP7_75t_L g3164 ( 
.A1(n_2986),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.C1(n_114),
.C2(n_115),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2787),
.Y(n_3165)
);

AND2x4_ASAP7_75t_L g3166 ( 
.A(n_3010),
.B(n_112),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2935),
.B(n_113),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2935),
.B(n_114),
.Y(n_3168)
);

OR2x6_ASAP7_75t_L g3169 ( 
.A(n_2957),
.B(n_1063),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2841),
.Y(n_3170)
);

A2O1A1Ixp33_ASAP7_75t_L g3171 ( 
.A1(n_2814),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_3171)
);

AOI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_2960),
.A2(n_1070),
.B1(n_1077),
.B2(n_1065),
.Y(n_3172)
);

OAI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_2944),
.A2(n_119),
.B1(n_116),
.B2(n_117),
.Y(n_3173)
);

OA21x2_ASAP7_75t_L g3174 ( 
.A1(n_2905),
.A2(n_120),
.B(n_123),
.Y(n_3174)
);

OAI22xp5_ASAP7_75t_L g3175 ( 
.A1(n_2897),
.A2(n_124),
.B1(n_120),
.B2(n_123),
.Y(n_3175)
);

CKINVDCx5p33_ASAP7_75t_R g3176 ( 
.A(n_2966),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2878),
.Y(n_3177)
);

BUFx3_ASAP7_75t_L g3178 ( 
.A(n_2966),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2956),
.B(n_125),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2966),
.B(n_125),
.Y(n_3180)
);

INVx3_ASAP7_75t_L g3181 ( 
.A(n_2960),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_2861),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2861),
.Y(n_3183)
);

AND2x2_ASAP7_75t_SL g3184 ( 
.A(n_2950),
.B(n_126),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2994),
.Y(n_3185)
);

AOI221xp5_ASAP7_75t_L g3186 ( 
.A1(n_2903),
.A2(n_3006),
.B1(n_2887),
.B2(n_2886),
.C(n_2823),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_3003),
.A2(n_1070),
.B1(n_1077),
.B2(n_1065),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_2924),
.A2(n_1070),
.B1(n_1077),
.B2(n_1065),
.Y(n_3188)
);

BUFx4f_ASAP7_75t_SL g3189 ( 
.A(n_2908),
.Y(n_3189)
);

OAI21x1_ASAP7_75t_L g3190 ( 
.A1(n_2801),
.A2(n_387),
.B(n_385),
.Y(n_3190)
);

AOI221xp5_ASAP7_75t_L g3191 ( 
.A1(n_2827),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.C(n_130),
.Y(n_3191)
);

AOI22xp33_ASAP7_75t_L g3192 ( 
.A1(n_2866),
.A2(n_1070),
.B1(n_1077),
.B2(n_1065),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2840),
.B(n_129),
.Y(n_3193)
);

NAND3x1_ASAP7_75t_L g3194 ( 
.A(n_2953),
.B(n_130),
.C(n_131),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2865),
.Y(n_3195)
);

OAI222xp33_ASAP7_75t_L g3196 ( 
.A1(n_2973),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.C1(n_136),
.C2(n_137),
.Y(n_3196)
);

OAI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2993),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_3197)
);

OR2x6_ASAP7_75t_L g3198 ( 
.A(n_2855),
.B(n_1070),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2994),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2953),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_3200)
);

INVx8_ASAP7_75t_L g3201 ( 
.A(n_2947),
.Y(n_3201)
);

AOI22xp5_ASAP7_75t_L g3202 ( 
.A1(n_2875),
.A2(n_1079),
.B1(n_1082),
.B2(n_1077),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_2873),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_3203)
);

AOI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_2976),
.A2(n_1082),
.B1(n_1079),
.B2(n_1206),
.Y(n_3204)
);

OR2x2_ASAP7_75t_SL g3205 ( 
.A(n_3170),
.B(n_2950),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3113),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3014),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_3060),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_3068),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_3024),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3104),
.Y(n_3211)
);

BUFx2_ASAP7_75t_SL g3212 ( 
.A(n_3086),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3025),
.Y(n_3213)
);

OAI21x1_ASAP7_75t_L g3214 ( 
.A1(n_3155),
.A2(n_2912),
.B(n_2952),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_3040),
.Y(n_3215)
);

BUFx3_ASAP7_75t_L g3216 ( 
.A(n_3012),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3016),
.B(n_2840),
.Y(n_3217)
);

BUFx3_ASAP7_75t_L g3218 ( 
.A(n_3089),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3045),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_3165),
.B(n_2838),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_3047),
.Y(n_3221)
);

INVx1_ASAP7_75t_SL g3222 ( 
.A(n_3030),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3058),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3092),
.B(n_2994),
.Y(n_3224)
);

OAI21x1_ASAP7_75t_L g3225 ( 
.A1(n_3160),
.A2(n_3195),
.B(n_3185),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3069),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3077),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3080),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3087),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3117),
.Y(n_3230)
);

OAI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_3171),
.A2(n_2816),
.B(n_2988),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3095),
.Y(n_3232)
);

CKINVDCx6p67_ASAP7_75t_R g3233 ( 
.A(n_3166),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_3103),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3021),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3035),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3041),
.Y(n_3237)
);

AO21x2_ASAP7_75t_L g3238 ( 
.A1(n_3199),
.A2(n_3009),
.B(n_3002),
.Y(n_3238)
);

HB1xp67_ASAP7_75t_L g3239 ( 
.A(n_3112),
.Y(n_3239)
);

OAI21x1_ASAP7_75t_L g3240 ( 
.A1(n_3105),
.A2(n_2796),
.B(n_3066),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3056),
.B(n_2947),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3044),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3097),
.Y(n_3243)
);

OAI21x1_ASAP7_75t_L g3244 ( 
.A1(n_3190),
.A2(n_2920),
.B(n_2808),
.Y(n_3244)
);

AOI21x1_ASAP7_75t_L g3245 ( 
.A1(n_3200),
.A2(n_2852),
.B(n_2977),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3120),
.B(n_3177),
.Y(n_3246)
);

OAI21x1_ASAP7_75t_L g3247 ( 
.A1(n_3043),
.A2(n_2922),
.B(n_2815),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_3065),
.Y(n_3248)
);

BUFx3_ASAP7_75t_L g3249 ( 
.A(n_3154),
.Y(n_3249)
);

OAI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_3032),
.A2(n_2989),
.B(n_2911),
.Y(n_3250)
);

AOI21x1_ASAP7_75t_L g3251 ( 
.A1(n_3200),
.A2(n_3193),
.B(n_3032),
.Y(n_3251)
);

INVx3_ASAP7_75t_SL g3252 ( 
.A(n_3013),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3127),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3145),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_3115),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3136),
.Y(n_3256)
);

HB1xp67_ASAP7_75t_L g3257 ( 
.A(n_3112),
.Y(n_3257)
);

BUFx2_ASAP7_75t_L g3258 ( 
.A(n_3094),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3052),
.Y(n_3259)
);

HB1xp67_ASAP7_75t_L g3260 ( 
.A(n_3033),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3074),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_3023),
.B(n_2840),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3143),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_3023),
.B(n_2803),
.Y(n_3264)
);

OR2x2_ASAP7_75t_L g3265 ( 
.A(n_3053),
.B(n_2838),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3111),
.Y(n_3266)
);

OA21x2_ASAP7_75t_L g3267 ( 
.A1(n_3019),
.A2(n_2837),
.B(n_2891),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3153),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3033),
.Y(n_3269)
);

INVxp67_ASAP7_75t_L g3270 ( 
.A(n_3161),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3144),
.A2(n_3000),
.B1(n_2968),
.B2(n_2954),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3079),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3090),
.B(n_2803),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3090),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3033),
.Y(n_3275)
);

BUFx2_ASAP7_75t_L g3276 ( 
.A(n_3094),
.Y(n_3276)
);

OAI21x1_ASAP7_75t_L g3277 ( 
.A1(n_3017),
.A2(n_2933),
.B(n_2820),
.Y(n_3277)
);

OR2x2_ASAP7_75t_L g3278 ( 
.A(n_3034),
.B(n_2838),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3034),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3072),
.Y(n_3280)
);

BUFx3_ASAP7_75t_L g3281 ( 
.A(n_3159),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3072),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3057),
.A2(n_2802),
.B(n_2889),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3162),
.Y(n_3284)
);

OAI21x1_ASAP7_75t_L g3285 ( 
.A1(n_3017),
.A2(n_2933),
.B(n_2860),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3174),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3174),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3184),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3134),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_3015),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3134),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3099),
.B(n_2803),
.Y(n_3292)
);

BUFx3_ASAP7_75t_L g3293 ( 
.A(n_3015),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3148),
.Y(n_3294)
);

CKINVDCx5p33_ASAP7_75t_R g3295 ( 
.A(n_3028),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3101),
.B(n_2953),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3062),
.A2(n_2907),
.B(n_2931),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3134),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3109),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3129),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3022),
.Y(n_3301)
);

AND2x4_ASAP7_75t_L g3302 ( 
.A(n_3110),
.B(n_2898),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3148),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3148),
.Y(n_3304)
);

OAI21xp33_ASAP7_75t_L g3305 ( 
.A1(n_3164),
.A2(n_2943),
.B(n_2927),
.Y(n_3305)
);

CKINVDCx6p67_ASAP7_75t_R g3306 ( 
.A(n_3166),
.Y(n_3306)
);

INVx2_ASAP7_75t_SL g3307 ( 
.A(n_3039),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3110),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3076),
.Y(n_3309)
);

OAI21x1_ASAP7_75t_L g3310 ( 
.A1(n_3020),
.A2(n_2882),
.B(n_2824),
.Y(n_3310)
);

OR2x2_ASAP7_75t_L g3311 ( 
.A(n_3110),
.B(n_2914),
.Y(n_3311)
);

INVx3_ASAP7_75t_L g3312 ( 
.A(n_3018),
.Y(n_3312)
);

OAI21x1_ASAP7_75t_L g3313 ( 
.A1(n_3020),
.A2(n_2829),
.B(n_2845),
.Y(n_3313)
);

AOI21x1_ASAP7_75t_L g3314 ( 
.A1(n_3073),
.A2(n_2845),
.B(n_2871),
.Y(n_3314)
);

BUFx3_ASAP7_75t_L g3315 ( 
.A(n_3054),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3081),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3178),
.Y(n_3317)
);

INVx3_ASAP7_75t_L g3318 ( 
.A(n_3018),
.Y(n_3318)
);

INVx2_ASAP7_75t_SL g3319 ( 
.A(n_3039),
.Y(n_3319)
);

BUFx6f_ASAP7_75t_L g3320 ( 
.A(n_3108),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3039),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3108),
.Y(n_3322)
);

INVx3_ASAP7_75t_L g3323 ( 
.A(n_3131),
.Y(n_3323)
);

AO21x2_ASAP7_75t_L g3324 ( 
.A1(n_3093),
.A2(n_2992),
.B(n_2880),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3061),
.B(n_2914),
.Y(n_3325)
);

BUFx2_ASAP7_75t_L g3326 ( 
.A(n_3181),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_3088),
.B(n_2898),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3131),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3131),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3181),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3133),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3169),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3194),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3169),
.Y(n_3334)
);

OAI21x1_ASAP7_75t_L g3335 ( 
.A1(n_3049),
.A2(n_2939),
.B(n_2857),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3169),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_3125),
.B(n_2898),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3124),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3167),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3106),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3125),
.Y(n_3341)
);

HB1xp67_ASAP7_75t_L g3342 ( 
.A(n_3128),
.Y(n_3342)
);

BUFx12f_ASAP7_75t_L g3343 ( 
.A(n_3056),
.Y(n_3343)
);

BUFx2_ASAP7_75t_L g3344 ( 
.A(n_3055),
.Y(n_3344)
);

INVx2_ASAP7_75t_SL g3345 ( 
.A(n_3141),
.Y(n_3345)
);

OR2x6_ASAP7_75t_L g3346 ( 
.A(n_3201),
.B(n_2946),
.Y(n_3346)
);

CKINVDCx5p33_ASAP7_75t_R g3347 ( 
.A(n_3176),
.Y(n_3347)
);

INVx3_ASAP7_75t_L g3348 ( 
.A(n_3038),
.Y(n_3348)
);

INVx2_ASAP7_75t_SL g3349 ( 
.A(n_3201),
.Y(n_3349)
);

BUFx3_ASAP7_75t_L g3350 ( 
.A(n_3137),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3168),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3064),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3098),
.B(n_2914),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3064),
.Y(n_3354)
);

INVxp67_ASAP7_75t_L g3355 ( 
.A(n_3179),
.Y(n_3355)
);

BUFx2_ASAP7_75t_SL g3356 ( 
.A(n_3082),
.Y(n_3356)
);

INVx3_ASAP7_75t_L g3357 ( 
.A(n_3142),
.Y(n_3357)
);

OAI21x1_ASAP7_75t_L g3358 ( 
.A1(n_3063),
.A2(n_2826),
.B(n_2934),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3107),
.B(n_2826),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3100),
.B(n_2826),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3126),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3029),
.B(n_144),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3119),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3114),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3198),
.Y(n_3365)
);

NOR2xp33_ASAP7_75t_L g3366 ( 
.A(n_3252),
.B(n_3189),
.Y(n_3366)
);

AOI222xp33_ASAP7_75t_L g3367 ( 
.A1(n_3333),
.A2(n_3121),
.B1(n_3140),
.B2(n_3151),
.C1(n_3149),
.C2(n_3026),
.Y(n_3367)
);

AOI22xp5_ASAP7_75t_L g3368 ( 
.A1(n_3305),
.A2(n_3062),
.B1(n_3164),
.B2(n_3150),
.Y(n_3368)
);

AOI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3283),
.A2(n_3150),
.B1(n_3121),
.B2(n_3119),
.Y(n_3369)
);

AOI221xp5_ASAP7_75t_L g3370 ( 
.A1(n_3352),
.A2(n_3354),
.B1(n_3333),
.B2(n_3140),
.C(n_3288),
.Y(n_3370)
);

BUFx2_ASAP7_75t_R g3371 ( 
.A(n_3281),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_3231),
.A2(n_3059),
.B1(n_3027),
.B2(n_3191),
.Y(n_3372)
);

CKINVDCx5p33_ASAP7_75t_R g3373 ( 
.A(n_3295),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3363),
.A2(n_3036),
.B1(n_3037),
.B2(n_3075),
.Y(n_3374)
);

OR2x2_ASAP7_75t_L g3375 ( 
.A(n_3239),
.B(n_3257),
.Y(n_3375)
);

AOI221xp5_ASAP7_75t_L g3376 ( 
.A1(n_3352),
.A2(n_3139),
.B1(n_3011),
.B2(n_3175),
.C(n_3197),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3258),
.B(n_3084),
.Y(n_3377)
);

AOI21xp33_ASAP7_75t_L g3378 ( 
.A1(n_3354),
.A2(n_3091),
.B(n_3102),
.Y(n_3378)
);

AOI222xp33_ASAP7_75t_L g3379 ( 
.A1(n_3288),
.A2(n_3175),
.B1(n_3196),
.B2(n_3186),
.C1(n_3132),
.C2(n_3122),
.Y(n_3379)
);

AOI21xp33_ASAP7_75t_L g3380 ( 
.A1(n_3303),
.A2(n_3036),
.B(n_3078),
.Y(n_3380)
);

OA21x2_ASAP7_75t_L g3381 ( 
.A1(n_3279),
.A2(n_3298),
.B(n_3291),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3330),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3296),
.A2(n_3297),
.B1(n_3344),
.B2(n_3146),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3296),
.A2(n_3156),
.B1(n_3031),
.B2(n_3163),
.Y(n_3384)
);

AOI21xp33_ASAP7_75t_L g3385 ( 
.A1(n_3303),
.A2(n_3116),
.B(n_3050),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3210),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_3258),
.B(n_3083),
.Y(n_3387)
);

AOI222xp33_ASAP7_75t_L g3388 ( 
.A1(n_3344),
.A2(n_3270),
.B1(n_3355),
.B2(n_3361),
.C1(n_3250),
.C2(n_3173),
.Y(n_3388)
);

AOI22xp33_ASAP7_75t_L g3389 ( 
.A1(n_3364),
.A2(n_3042),
.B1(n_3046),
.B2(n_3082),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_3324),
.A2(n_3093),
.B(n_3116),
.Y(n_3390)
);

AND2x2_ASAP7_75t_L g3391 ( 
.A(n_3276),
.B(n_3118),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3210),
.Y(n_3392)
);

OAI22xp5_ASAP7_75t_L g3393 ( 
.A1(n_3222),
.A2(n_3051),
.B1(n_3123),
.B2(n_3182),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_SL g3394 ( 
.A1(n_3348),
.A2(n_3180),
.B1(n_3157),
.B2(n_3082),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3330),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3215),
.Y(n_3396)
);

INVx3_ASAP7_75t_L g3397 ( 
.A(n_3320),
.Y(n_3397)
);

OAI211xp5_ASAP7_75t_L g3398 ( 
.A1(n_3251),
.A2(n_3286),
.B(n_3287),
.C(n_3070),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3276),
.B(n_3142),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_3364),
.A2(n_3082),
.B1(n_3048),
.B2(n_3203),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_3218),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_L g3402 ( 
.A(n_3252),
.B(n_3343),
.Y(n_3402)
);

OAI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_3233),
.A2(n_3306),
.B1(n_3271),
.B2(n_3251),
.Y(n_3403)
);

OAI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3233),
.A2(n_3067),
.B1(n_3183),
.B2(n_3202),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3282),
.B(n_3157),
.Y(n_3405)
);

OAI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3306),
.A2(n_3201),
.B1(n_3172),
.B2(n_3085),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3215),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3221),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3346),
.A2(n_3135),
.B1(n_3152),
.B2(n_3187),
.Y(n_3409)
);

OAI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_3346),
.A2(n_3348),
.B1(n_3341),
.B2(n_3338),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_R g3411 ( 
.A(n_3295),
.B(n_3347),
.Y(n_3411)
);

AOI33xp33_ASAP7_75t_L g3412 ( 
.A1(n_3286),
.A2(n_3180),
.A3(n_3071),
.B1(n_3096),
.B2(n_3138),
.B3(n_3147),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3272),
.B(n_3198),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3221),
.Y(n_3414)
);

AOI22xp33_ASAP7_75t_L g3415 ( 
.A1(n_3308),
.A2(n_3198),
.B1(n_3158),
.B2(n_3130),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3346),
.A2(n_3192),
.B1(n_3188),
.B2(n_3204),
.Y(n_3416)
);

AOI221xp5_ASAP7_75t_L g3417 ( 
.A1(n_3287),
.A2(n_3263),
.B1(n_3224),
.B2(n_3261),
.C(n_3275),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3280),
.B(n_145),
.Y(n_3418)
);

AOI221xp5_ASAP7_75t_L g3419 ( 
.A1(n_3263),
.A2(n_2863),
.B1(n_150),
.B2(n_146),
.C(n_148),
.Y(n_3419)
);

OR2x2_ASAP7_75t_L g3420 ( 
.A(n_3248),
.B(n_148),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3227),
.Y(n_3421)
);

INVx3_ASAP7_75t_L g3422 ( 
.A(n_3320),
.Y(n_3422)
);

AOI221xp5_ASAP7_75t_L g3423 ( 
.A1(n_3261),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_3423)
);

AOI221xp5_ASAP7_75t_L g3424 ( 
.A1(n_3266),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_3424)
);

OAI211xp5_ASAP7_75t_SL g3425 ( 
.A1(n_3304),
.A2(n_159),
.B(n_156),
.C(n_157),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3227),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3308),
.A2(n_1082),
.B1(n_1079),
.B2(n_1108),
.Y(n_3427)
);

CKINVDCx5p33_ASAP7_75t_R g3428 ( 
.A(n_3212),
.Y(n_3428)
);

AOI221xp5_ASAP7_75t_L g3429 ( 
.A1(n_3304),
.A2(n_159),
.B1(n_156),
.B2(n_157),
.C(n_160),
.Y(n_3429)
);

OAI22xp5_ASAP7_75t_L g3430 ( 
.A1(n_3346),
.A2(n_163),
.B1(n_160),
.B2(n_161),
.Y(n_3430)
);

OAI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_3348),
.A2(n_165),
.B1(n_161),
.B2(n_163),
.Y(n_3431)
);

BUFx2_ASAP7_75t_L g3432 ( 
.A(n_3343),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3320),
.Y(n_3433)
);

AOI22xp33_ASAP7_75t_L g3434 ( 
.A1(n_3338),
.A2(n_1082),
.B1(n_1079),
.B2(n_1108),
.Y(n_3434)
);

BUFx2_ASAP7_75t_L g3435 ( 
.A(n_3249),
.Y(n_3435)
);

AND2x4_ASAP7_75t_L g3436 ( 
.A(n_3289),
.B(n_3291),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3289),
.B(n_165),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3229),
.Y(n_3438)
);

CKINVDCx5p33_ASAP7_75t_R g3439 ( 
.A(n_3212),
.Y(n_3439)
);

OAI221xp5_ASAP7_75t_L g3440 ( 
.A1(n_3298),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.C(n_169),
.Y(n_3440)
);

INVx4_ASAP7_75t_L g3441 ( 
.A(n_3216),
.Y(n_3441)
);

OAI221xp5_ASAP7_75t_L g3442 ( 
.A1(n_3294),
.A2(n_166),
.B1(n_167),
.B2(n_170),
.C(n_171),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3324),
.A2(n_1082),
.B1(n_1079),
.B2(n_1108),
.Y(n_3443)
);

OAI221xp5_ASAP7_75t_L g3444 ( 
.A1(n_3260),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.C(n_174),
.Y(n_3444)
);

AOI22xp33_ASAP7_75t_SL g3445 ( 
.A1(n_3324),
.A2(n_177),
.B1(n_172),
.B2(n_175),
.Y(n_3445)
);

AOI222xp33_ASAP7_75t_L g3446 ( 
.A1(n_3325),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.C1(n_179),
.C2(n_180),
.Y(n_3446)
);

AND2x4_ASAP7_75t_L g3447 ( 
.A(n_3336),
.B(n_178),
.Y(n_3447)
);

CKINVDCx20_ASAP7_75t_R g3448 ( 
.A(n_3218),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_SL g3449 ( 
.A1(n_3217),
.A2(n_184),
.B1(n_179),
.B2(n_182),
.Y(n_3449)
);

AO21x2_ASAP7_75t_L g3450 ( 
.A1(n_3279),
.A2(n_182),
.B(n_184),
.Y(n_3450)
);

INVx4_ASAP7_75t_L g3451 ( 
.A(n_3216),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3269),
.A2(n_3341),
.B1(n_3340),
.B2(n_3339),
.Y(n_3452)
);

AOI221xp5_ASAP7_75t_L g3453 ( 
.A1(n_3211),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.C(n_188),
.Y(n_3453)
);

OAI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3281),
.A2(n_3350),
.B1(n_3351),
.B2(n_3339),
.Y(n_3454)
);

INVx4_ASAP7_75t_L g3455 ( 
.A(n_3315),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3229),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3269),
.A2(n_1109),
.B1(n_1147),
.B2(n_1108),
.Y(n_3457)
);

CKINVDCx5p33_ASAP7_75t_R g3458 ( 
.A(n_3347),
.Y(n_3458)
);

CKINVDCx5p33_ASAP7_75t_R g3459 ( 
.A(n_3315),
.Y(n_3459)
);

AOI222xp33_ASAP7_75t_L g3460 ( 
.A1(n_3217),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.C1(n_190),
.C2(n_191),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3336),
.B(n_190),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3326),
.Y(n_3462)
);

BUFx2_ASAP7_75t_L g3463 ( 
.A(n_3249),
.Y(n_3463)
);

OAI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3350),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_3351),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_3465)
);

AOI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3340),
.A2(n_1109),
.B1(n_1147),
.B2(n_1108),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_L g3467 ( 
.A1(n_3331),
.A2(n_1147),
.B1(n_1148),
.B2(n_1109),
.Y(n_3467)
);

INVx8_ASAP7_75t_L g3468 ( 
.A(n_3320),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3207),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3248),
.B(n_194),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_SL g3471 ( 
.A1(n_3267),
.A2(n_201),
.B1(n_198),
.B2(n_200),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3326),
.Y(n_3472)
);

BUFx6f_ASAP7_75t_L g3473 ( 
.A(n_3320),
.Y(n_3473)
);

NAND3xp33_ASAP7_75t_L g3474 ( 
.A(n_3359),
.B(n_198),
.C(n_201),
.Y(n_3474)
);

CKINVDCx11_ASAP7_75t_R g3475 ( 
.A(n_3293),
.Y(n_3475)
);

AOI22xp33_ASAP7_75t_L g3476 ( 
.A1(n_3331),
.A2(n_1147),
.B1(n_1148),
.B2(n_1109),
.Y(n_3476)
);

AOI22xp33_ASAP7_75t_SL g3477 ( 
.A1(n_3267),
.A2(n_205),
.B1(n_202),
.B2(n_203),
.Y(n_3477)
);

HB1xp67_ASAP7_75t_L g3478 ( 
.A(n_3264),
.Y(n_3478)
);

OAI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3349),
.A2(n_206),
.B1(n_203),
.B2(n_205),
.Y(n_3479)
);

AOI22xp33_ASAP7_75t_L g3480 ( 
.A1(n_3337),
.A2(n_3365),
.B1(n_3267),
.B2(n_3327),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3207),
.Y(n_3481)
);

OAI211xp5_ASAP7_75t_SL g3482 ( 
.A1(n_3241),
.A2(n_209),
.B(n_206),
.C(n_207),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3337),
.A2(n_1147),
.B1(n_1148),
.B2(n_1109),
.Y(n_3483)
);

CKINVDCx14_ASAP7_75t_R g3484 ( 
.A(n_3342),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3322),
.Y(n_3485)
);

AOI22xp33_ASAP7_75t_L g3486 ( 
.A1(n_3337),
.A2(n_1159),
.B1(n_1148),
.B2(n_1230),
.Y(n_3486)
);

AOI221xp5_ASAP7_75t_L g3487 ( 
.A1(n_3230),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.C(n_212),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3322),
.Y(n_3488)
);

OAI221xp5_ASAP7_75t_SL g3489 ( 
.A1(n_3327),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.C(n_214),
.Y(n_3489)
);

AOI221xp5_ASAP7_75t_L g3490 ( 
.A1(n_3230),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.C(n_218),
.Y(n_3490)
);

AOI33xp33_ASAP7_75t_L g3491 ( 
.A1(n_3262),
.A2(n_3292),
.A3(n_3273),
.B1(n_3264),
.B2(n_3259),
.B3(n_3219),
.Y(n_3491)
);

OAI22xp5_ASAP7_75t_L g3492 ( 
.A1(n_3349),
.A2(n_3356),
.B1(n_3345),
.B2(n_3293),
.Y(n_3492)
);

AOI221xp5_ASAP7_75t_L g3493 ( 
.A1(n_3259),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_SL g3494 ( 
.A1(n_3267),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3292),
.B(n_3262),
.Y(n_3495)
);

AOI21x1_ASAP7_75t_L g3496 ( 
.A1(n_3328),
.A2(n_222),
.B(n_225),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_L g3497 ( 
.A1(n_3365),
.A2(n_1159),
.B1(n_1148),
.B2(n_1230),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3381),
.Y(n_3498)
);

NOR2xp33_ASAP7_75t_L g3499 ( 
.A(n_3371),
.B(n_3345),
.Y(n_3499)
);

AOI21x1_ASAP7_75t_L g3500 ( 
.A1(n_3432),
.A2(n_3362),
.B(n_3328),
.Y(n_3500)
);

INVxp67_ASAP7_75t_L g3501 ( 
.A(n_3435),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3478),
.B(n_3312),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3478),
.B(n_3312),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3391),
.B(n_3312),
.Y(n_3504)
);

BUFx2_ASAP7_75t_L g3505 ( 
.A(n_3441),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3370),
.B(n_3246),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3469),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3436),
.B(n_3318),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3397),
.B(n_3422),
.Y(n_3509)
);

INVx2_ASAP7_75t_SL g3510 ( 
.A(n_3468),
.Y(n_3510)
);

BUFx3_ASAP7_75t_L g3511 ( 
.A(n_3475),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3495),
.B(n_3205),
.Y(n_3512)
);

INVx2_ASAP7_75t_SL g3513 ( 
.A(n_3468),
.Y(n_3513)
);

AND2x4_ASAP7_75t_L g3514 ( 
.A(n_3397),
.B(n_3332),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3381),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3481),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3386),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3436),
.B(n_3318),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3422),
.B(n_3318),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3433),
.B(n_3273),
.Y(n_3520)
);

AND2x4_ASAP7_75t_L g3521 ( 
.A(n_3433),
.B(n_3473),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3392),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3368),
.A2(n_3302),
.B1(n_3334),
.B2(n_3332),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3382),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3395),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3462),
.B(n_3472),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3407),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3399),
.B(n_3357),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3387),
.B(n_3357),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3421),
.Y(n_3530)
);

INVx2_ASAP7_75t_SL g3531 ( 
.A(n_3468),
.Y(n_3531)
);

AOI222xp33_ASAP7_75t_L g3532 ( 
.A1(n_3376),
.A2(n_3362),
.B1(n_3353),
.B2(n_3360),
.C1(n_3246),
.C2(n_3302),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3426),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3438),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3396),
.Y(n_3535)
);

INVx3_ASAP7_75t_L g3536 ( 
.A(n_3473),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3408),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3463),
.B(n_3357),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3414),
.Y(n_3539)
);

BUFx3_ASAP7_75t_L g3540 ( 
.A(n_3428),
.Y(n_3540)
);

OA21x2_ASAP7_75t_L g3541 ( 
.A1(n_3390),
.A2(n_3240),
.B(n_3225),
.Y(n_3541)
);

INVx3_ASAP7_75t_L g3542 ( 
.A(n_3473),
.Y(n_3542)
);

AND2x4_ASAP7_75t_SL g3543 ( 
.A(n_3441),
.B(n_3302),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3485),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3491),
.B(n_3290),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3488),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3456),
.Y(n_3547)
);

INVx3_ASAP7_75t_L g3548 ( 
.A(n_3451),
.Y(n_3548)
);

HB1xp67_ASAP7_75t_L g3549 ( 
.A(n_3375),
.Y(n_3549)
);

AOI222xp33_ASAP7_75t_L g3550 ( 
.A1(n_3429),
.A2(n_3353),
.B1(n_3360),
.B2(n_3213),
.C1(n_3206),
.C2(n_3226),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3450),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3410),
.B(n_3290),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3450),
.Y(n_3553)
);

OR2x2_ASAP7_75t_L g3554 ( 
.A(n_3398),
.B(n_3205),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3420),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3480),
.B(n_3321),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3398),
.Y(n_3557)
);

AND2x4_ASAP7_75t_L g3558 ( 
.A(n_3390),
.B(n_3334),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3470),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3413),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3447),
.Y(n_3561)
);

AND2x2_ASAP7_75t_L g3562 ( 
.A(n_3377),
.B(n_3403),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3437),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3447),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3405),
.B(n_3452),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3492),
.Y(n_3566)
);

HB1xp67_ASAP7_75t_L g3567 ( 
.A(n_3484),
.Y(n_3567)
);

AO22x1_ASAP7_75t_L g3568 ( 
.A1(n_3451),
.A2(n_3323),
.B1(n_3329),
.B2(n_3321),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3454),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3454),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3496),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3461),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3418),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3417),
.B(n_3329),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3455),
.B(n_3284),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3388),
.B(n_3223),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3378),
.B(n_3223),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3461),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3474),
.Y(n_3579)
);

AND2x4_ASAP7_75t_L g3580 ( 
.A(n_3455),
.B(n_3220),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3385),
.B(n_3299),
.Y(n_3581)
);

HB1xp67_ASAP7_75t_L g3582 ( 
.A(n_3401),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3445),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3439),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3445),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3394),
.B(n_3299),
.Y(n_3586)
);

OAI322xp33_ASAP7_75t_L g3587 ( 
.A1(n_3369),
.A2(n_3464),
.A3(n_3440),
.B1(n_3444),
.B2(n_3442),
.C1(n_3404),
.C2(n_3431),
.Y(n_3587)
);

OR2x2_ASAP7_75t_L g3588 ( 
.A(n_3380),
.B(n_3265),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3394),
.B(n_3300),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3471),
.B(n_3300),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3471),
.B(n_3317),
.Y(n_3591)
);

NOR2x1_ASAP7_75t_L g3592 ( 
.A(n_3402),
.B(n_3356),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3477),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_3477),
.B(n_3317),
.Y(n_3594)
);

BUFx6f_ASAP7_75t_L g3595 ( 
.A(n_3459),
.Y(n_3595)
);

INVxp67_ASAP7_75t_L g3596 ( 
.A(n_3430),
.Y(n_3596)
);

AND2x4_ASAP7_75t_L g3597 ( 
.A(n_3448),
.B(n_3220),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3383),
.B(n_3226),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3494),
.B(n_3274),
.Y(n_3599)
);

INVxp67_ASAP7_75t_L g3600 ( 
.A(n_3366),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3458),
.Y(n_3601)
);

INVxp67_ASAP7_75t_L g3602 ( 
.A(n_3379),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3494),
.Y(n_3603)
);

AO21x2_ASAP7_75t_L g3604 ( 
.A1(n_3404),
.A2(n_3225),
.B(n_3314),
.Y(n_3604)
);

OR2x2_ASAP7_75t_L g3605 ( 
.A(n_3443),
.B(n_3265),
.Y(n_3605)
);

AND2x4_ASAP7_75t_L g3606 ( 
.A(n_3389),
.B(n_3220),
.Y(n_3606)
);

HB1xp67_ASAP7_75t_L g3607 ( 
.A(n_3393),
.Y(n_3607)
);

AO21x2_ASAP7_75t_L g3608 ( 
.A1(n_3464),
.A2(n_3425),
.B(n_3482),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3449),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3374),
.B(n_3323),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3383),
.B(n_3323),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3449),
.Y(n_3612)
);

HB1xp67_ASAP7_75t_L g3613 ( 
.A(n_3411),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3412),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3406),
.Y(n_3615)
);

OR2x2_ASAP7_75t_L g3616 ( 
.A(n_3486),
.B(n_3208),
.Y(n_3616)
);

INVxp67_ASAP7_75t_L g3617 ( 
.A(n_3367),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3483),
.B(n_3307),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3415),
.B(n_3307),
.Y(n_3619)
);

BUFx2_ASAP7_75t_L g3620 ( 
.A(n_3373),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3400),
.B(n_3319),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3372),
.B(n_3319),
.Y(n_3622)
);

OAI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_3384),
.A2(n_3311),
.B1(n_3301),
.B2(n_3309),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3406),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3479),
.Y(n_3625)
);

AOI221xp5_ASAP7_75t_L g3626 ( 
.A1(n_3557),
.A2(n_3617),
.B1(n_3602),
.B2(n_3587),
.C(n_3614),
.Y(n_3626)
);

AOI22xp5_ASAP7_75t_L g3627 ( 
.A1(n_3557),
.A2(n_3446),
.B1(n_3460),
.B2(n_3493),
.Y(n_3627)
);

AOI22xp33_ASAP7_75t_SL g3628 ( 
.A1(n_3607),
.A2(n_3593),
.B1(n_3603),
.B2(n_3583),
.Y(n_3628)
);

NOR2x1_ASAP7_75t_L g3629 ( 
.A(n_3548),
.B(n_3425),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3507),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3507),
.Y(n_3631)
);

BUFx2_ASAP7_75t_L g3632 ( 
.A(n_3567),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_L g3633 ( 
.A1(n_3614),
.A2(n_3419),
.B1(n_3453),
.B2(n_3482),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_L g3634 ( 
.A(n_3511),
.B(n_3489),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3516),
.Y(n_3635)
);

AOI22xp33_ASAP7_75t_L g3636 ( 
.A1(n_3593),
.A2(n_3487),
.B1(n_3490),
.B2(n_3423),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_SL g3637 ( 
.A1(n_3585),
.A2(n_3409),
.B1(n_3416),
.B2(n_3489),
.Y(n_3637)
);

AOI22xp33_ASAP7_75t_SL g3638 ( 
.A1(n_3609),
.A2(n_3335),
.B1(n_3240),
.B2(n_3311),
.Y(n_3638)
);

AOI22xp33_ASAP7_75t_L g3639 ( 
.A1(n_3608),
.A2(n_3424),
.B1(n_3465),
.B2(n_3335),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_3576),
.A2(n_3465),
.B(n_3206),
.Y(n_3640)
);

OR2x2_ASAP7_75t_L g3641 ( 
.A(n_3549),
.B(n_3228),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3555),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_L g3643 ( 
.A1(n_3608),
.A2(n_3609),
.B1(n_3612),
.B2(n_3615),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3555),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3522),
.Y(n_3645)
);

AOI222xp33_ASAP7_75t_L g3646 ( 
.A1(n_3612),
.A2(n_3358),
.B1(n_3427),
.B2(n_3253),
.C1(n_3254),
.C2(n_3434),
.Y(n_3646)
);

AOI22xp33_ASAP7_75t_L g3647 ( 
.A1(n_3608),
.A2(n_3358),
.B1(n_3466),
.B2(n_3457),
.Y(n_3647)
);

AOI221xp5_ASAP7_75t_L g3648 ( 
.A1(n_3579),
.A2(n_3554),
.B1(n_3598),
.B2(n_3596),
.C(n_3623),
.Y(n_3648)
);

OAI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_3554),
.A2(n_3506),
.B1(n_3624),
.B2(n_3523),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3571),
.B(n_3228),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3550),
.A2(n_3238),
.B1(n_3497),
.B2(n_3316),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3504),
.B(n_3232),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3548),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3548),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3505),
.Y(n_3655)
);

OR2x2_ASAP7_75t_L g3656 ( 
.A(n_3512),
.B(n_3253),
.Y(n_3656)
);

AOI33xp33_ASAP7_75t_L g3657 ( 
.A1(n_3569),
.A2(n_3232),
.A3(n_3254),
.B1(n_3476),
.B2(n_3467),
.B3(n_3242),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3522),
.Y(n_3658)
);

OAI221xp5_ASAP7_75t_L g3659 ( 
.A1(n_3532),
.A2(n_3242),
.B1(n_3235),
.B2(n_3236),
.C(n_3237),
.Y(n_3659)
);

OAI221xp5_ASAP7_75t_L g3660 ( 
.A1(n_3592),
.A2(n_3243),
.B1(n_3235),
.B2(n_3236),
.C(n_3237),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3551),
.B(n_3208),
.Y(n_3661)
);

AOI221xp5_ASAP7_75t_L g3662 ( 
.A1(n_3577),
.A2(n_3243),
.B1(n_3209),
.B2(n_3255),
.C(n_3256),
.Y(n_3662)
);

OAI222xp33_ASAP7_75t_L g3663 ( 
.A1(n_3570),
.A2(n_3314),
.B1(n_3245),
.B2(n_3278),
.C1(n_3209),
.C2(n_3255),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3606),
.A2(n_3238),
.B1(n_3278),
.B2(n_3313),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3505),
.Y(n_3665)
);

BUFx3_ASAP7_75t_L g3666 ( 
.A(n_3511),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3551),
.B(n_3234),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3504),
.B(n_3268),
.Y(n_3668)
);

OAI211xp5_ASAP7_75t_L g3669 ( 
.A1(n_3611),
.A2(n_3245),
.B(n_3256),
.C(n_3313),
.Y(n_3669)
);

OA21x2_ASAP7_75t_L g3670 ( 
.A1(n_3498),
.A2(n_3247),
.B(n_3277),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3512),
.B(n_3234),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3529),
.B(n_3552),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3553),
.B(n_3611),
.Y(n_3673)
);

INVxp67_ASAP7_75t_L g3674 ( 
.A(n_3582),
.Y(n_3674)
);

AOI31xp33_ASAP7_75t_L g3675 ( 
.A1(n_3613),
.A2(n_3268),
.A3(n_3247),
.B(n_3285),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3509),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3527),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3553),
.B(n_3238),
.Y(n_3678)
);

OA222x2_ASAP7_75t_L g3679 ( 
.A1(n_3588),
.A2(n_3285),
.B1(n_3277),
.B2(n_3310),
.C1(n_3244),
.C2(n_3214),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_SL g3680 ( 
.A1(n_3562),
.A2(n_3244),
.B1(n_3310),
.B2(n_3214),
.Y(n_3680)
);

NAND4xp25_ASAP7_75t_L g3681 ( 
.A(n_3622),
.B(n_228),
.C(n_226),
.D(n_227),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3529),
.B(n_226),
.Y(n_3682)
);

OAI221xp5_ASAP7_75t_L g3683 ( 
.A1(n_3600),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.C(n_230),
.Y(n_3683)
);

HB1xp67_ASAP7_75t_L g3684 ( 
.A(n_3501),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3527),
.Y(n_3685)
);

OAI211xp5_ASAP7_75t_L g3686 ( 
.A1(n_3588),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_3686)
);

OAI211xp5_ASAP7_75t_SL g3687 ( 
.A1(n_3560),
.A2(n_3566),
.B(n_3625),
.C(n_3563),
.Y(n_3687)
);

OAI211xp5_ASAP7_75t_L g3688 ( 
.A1(n_3622),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3530),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_SL g3690 ( 
.A1(n_3562),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3509),
.Y(n_3691)
);

OAI22xp5_ASAP7_75t_L g3692 ( 
.A1(n_3625),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_3692)
);

BUFx2_ASAP7_75t_L g3693 ( 
.A(n_3620),
.Y(n_3693)
);

OAI221xp5_ASAP7_75t_L g3694 ( 
.A1(n_3560),
.A2(n_3499),
.B1(n_3545),
.B2(n_3531),
.C(n_3510),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3530),
.Y(n_3695)
);

OAI31xp33_ASAP7_75t_L g3696 ( 
.A1(n_3545),
.A2(n_235),
.A3(n_236),
.B(n_238),
.Y(n_3696)
);

OAI31xp33_ASAP7_75t_L g3697 ( 
.A1(n_3574),
.A2(n_238),
.A3(n_239),
.B(n_240),
.Y(n_3697)
);

AOI33xp33_ASAP7_75t_L g3698 ( 
.A1(n_3574),
.A2(n_3599),
.A3(n_3594),
.B1(n_3590),
.B2(n_3591),
.B3(n_3558),
.Y(n_3698)
);

NAND3xp33_ASAP7_75t_L g3699 ( 
.A(n_3581),
.B(n_3605),
.C(n_3610),
.Y(n_3699)
);

OAI22xp5_ASAP7_75t_L g3700 ( 
.A1(n_3561),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_3700)
);

OAI221xp5_ASAP7_75t_SL g3701 ( 
.A1(n_3590),
.A2(n_241),
.B1(n_243),
.B2(n_245),
.C(n_246),
.Y(n_3701)
);

AOI22xp33_ASAP7_75t_SL g3702 ( 
.A1(n_3606),
.A2(n_243),
.B1(n_245),
.B2(n_247),
.Y(n_3702)
);

NAND3xp33_ASAP7_75t_L g3703 ( 
.A(n_3581),
.B(n_247),
.C(n_248),
.Y(n_3703)
);

AOI211xp5_ASAP7_75t_L g3704 ( 
.A1(n_3591),
.A2(n_248),
.B(n_249),
.C(n_251),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3533),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3533),
.Y(n_3706)
);

INVx1_ASAP7_75t_SL g3707 ( 
.A(n_3620),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3534),
.Y(n_3708)
);

INVx2_ASAP7_75t_SL g3709 ( 
.A(n_3595),
.Y(n_3709)
);

NOR2xp67_ASAP7_75t_L g3710 ( 
.A(n_3500),
.B(n_251),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3534),
.Y(n_3711)
);

NOR2xp67_ASAP7_75t_L g3712 ( 
.A(n_3500),
.B(n_252),
.Y(n_3712)
);

OAI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3561),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_3713)
);

INVxp67_ASAP7_75t_SL g3714 ( 
.A(n_3584),
.Y(n_3714)
);

OAI221xp5_ASAP7_75t_L g3715 ( 
.A1(n_3510),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.C(n_260),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3509),
.Y(n_3716)
);

INVx1_ASAP7_75t_SL g3717 ( 
.A(n_3595),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3536),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3564),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_3719)
);

OAI211xp5_ASAP7_75t_L g3720 ( 
.A1(n_3594),
.A2(n_261),
.B(n_262),
.C(n_264),
.Y(n_3720)
);

AOI22xp5_ASAP7_75t_L g3721 ( 
.A1(n_3586),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_3721)
);

NAND3xp33_ASAP7_75t_L g3722 ( 
.A(n_3605),
.B(n_265),
.C(n_267),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3536),
.Y(n_3723)
);

OAI22xp5_ASAP7_75t_L g3724 ( 
.A1(n_3564),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_3724)
);

OA21x2_ASAP7_75t_L g3725 ( 
.A1(n_3498),
.A2(n_270),
.B(n_271),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3547),
.Y(n_3726)
);

AOI22xp33_ASAP7_75t_SL g3727 ( 
.A1(n_3606),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3547),
.Y(n_3728)
);

NAND2xp33_ASAP7_75t_R g3729 ( 
.A(n_3601),
.B(n_272),
.Y(n_3729)
);

AOI22xp33_ASAP7_75t_L g3730 ( 
.A1(n_3565),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3599),
.B(n_274),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3559),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3559),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3517),
.Y(n_3734)
);

AOI221xp5_ASAP7_75t_L g3735 ( 
.A1(n_3558),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.C(n_279),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_3595),
.Y(n_3736)
);

OAI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3572),
.A2(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_3737)
);

OAI211xp5_ASAP7_75t_L g3738 ( 
.A1(n_3586),
.A2(n_280),
.B(n_281),
.C(n_282),
.Y(n_3738)
);

INVx4_ASAP7_75t_L g3739 ( 
.A(n_3595),
.Y(n_3739)
);

INVxp67_ASAP7_75t_L g3740 ( 
.A(n_3621),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3632),
.B(n_3552),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3693),
.Y(n_3742)
);

BUFx2_ASAP7_75t_L g3743 ( 
.A(n_3739),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3630),
.Y(n_3744)
);

OR2x2_ASAP7_75t_L g3745 ( 
.A(n_3673),
.B(n_3684),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3631),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3645),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3658),
.Y(n_3748)
);

OR2x2_ASAP7_75t_L g3749 ( 
.A(n_3673),
.B(n_3535),
.Y(n_3749)
);

BUFx2_ASAP7_75t_L g3750 ( 
.A(n_3739),
.Y(n_3750)
);

AND2x4_ASAP7_75t_L g3751 ( 
.A(n_3707),
.B(n_3589),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3672),
.B(n_3508),
.Y(n_3752)
);

OR2x2_ASAP7_75t_L g3753 ( 
.A(n_3740),
.B(n_3674),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3677),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3709),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3714),
.B(n_3508),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3736),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3676),
.B(n_3518),
.Y(n_3758)
);

HB1xp67_ASAP7_75t_L g3759 ( 
.A(n_3710),
.Y(n_3759)
);

AND2x4_ASAP7_75t_L g3760 ( 
.A(n_3691),
.B(n_3589),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3634),
.B(n_3610),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3716),
.B(n_3518),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3666),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3685),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3696),
.B(n_3572),
.Y(n_3765)
);

BUFx2_ASAP7_75t_L g3766 ( 
.A(n_3629),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3655),
.B(n_3665),
.Y(n_3767)
);

OR2x2_ASAP7_75t_L g3768 ( 
.A(n_3656),
.B(n_3535),
.Y(n_3768)
);

NAND2xp33_ASAP7_75t_R g3769 ( 
.A(n_3725),
.B(n_3601),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3652),
.B(n_3502),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3689),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3637),
.B(n_3578),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3695),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3705),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3668),
.B(n_3502),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3706),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3628),
.A2(n_3604),
.B1(n_3558),
.B2(n_3565),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3708),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3717),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3711),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3718),
.B(n_3503),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3723),
.B(n_3503),
.Y(n_3782)
);

OR2x2_ASAP7_75t_L g3783 ( 
.A(n_3641),
.B(n_3537),
.Y(n_3783)
);

INVxp67_ASAP7_75t_SL g3784 ( 
.A(n_3712),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3731),
.B(n_3595),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3726),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3653),
.B(n_3521),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_SL g3788 ( 
.A(n_3639),
.B(n_3597),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3698),
.B(n_3578),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3728),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_L g3791 ( 
.A(n_3731),
.B(n_3540),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3725),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3654),
.B(n_3521),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3732),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3638),
.B(n_3521),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3670),
.Y(n_3796)
);

AND2x4_ASAP7_75t_L g3797 ( 
.A(n_3642),
.B(n_3543),
.Y(n_3797)
);

OAI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3643),
.A2(n_3556),
.B(n_3621),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3733),
.B(n_3543),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3648),
.B(n_3619),
.Y(n_3800)
);

INVxp67_ASAP7_75t_SL g3801 ( 
.A(n_3729),
.Y(n_3801)
);

OR2x2_ASAP7_75t_L g3802 ( 
.A(n_3644),
.B(n_3537),
.Y(n_3802)
);

AND2x4_ASAP7_75t_L g3803 ( 
.A(n_3635),
.B(n_3513),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3682),
.B(n_3538),
.Y(n_3804)
);

NAND2x1_ASAP7_75t_L g3805 ( 
.A(n_3675),
.B(n_3580),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3671),
.B(n_3538),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3679),
.B(n_3519),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3670),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3680),
.B(n_3519),
.Y(n_3809)
);

INVx5_ASAP7_75t_L g3810 ( 
.A(n_3686),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3662),
.B(n_3536),
.Y(n_3811)
);

HB1xp67_ASAP7_75t_L g3812 ( 
.A(n_3650),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3640),
.B(n_3619),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3734),
.B(n_3542),
.Y(n_3814)
);

OR2x2_ASAP7_75t_L g3815 ( 
.A(n_3699),
.B(n_3539),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3650),
.Y(n_3816)
);

BUFx2_ASAP7_75t_L g3817 ( 
.A(n_3703),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3651),
.B(n_3542),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3649),
.B(n_3542),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3627),
.B(n_3573),
.Y(n_3820)
);

NOR2xp33_ASAP7_75t_L g3821 ( 
.A(n_3694),
.B(n_3540),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3649),
.B(n_3580),
.Y(n_3822)
);

OR2x2_ASAP7_75t_L g3823 ( 
.A(n_3661),
.B(n_3539),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3657),
.B(n_3580),
.Y(n_3824)
);

CKINVDCx5p33_ASAP7_75t_R g3825 ( 
.A(n_3690),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3697),
.B(n_3633),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3678),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3636),
.B(n_3556),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3626),
.B(n_3575),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3647),
.B(n_3528),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3661),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3721),
.B(n_3575),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3667),
.B(n_3528),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3743),
.B(n_3513),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3741),
.B(n_3531),
.Y(n_3835)
);

BUFx6f_ASAP7_75t_L g3836 ( 
.A(n_3743),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3741),
.B(n_3597),
.Y(n_3837)
);

NOR2x1p5_ASAP7_75t_L g3838 ( 
.A(n_3801),
.B(n_3763),
.Y(n_3838)
);

NAND3xp33_ASAP7_75t_L g3839 ( 
.A(n_3810),
.B(n_3704),
.C(n_3735),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3753),
.Y(n_3840)
);

NOR3xp33_ASAP7_75t_L g3841 ( 
.A(n_3766),
.B(n_3800),
.C(n_3828),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3810),
.B(n_3722),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3750),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3756),
.B(n_3597),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3810),
.A2(n_3720),
.B1(n_3738),
.B2(n_3681),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3756),
.B(n_3520),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3772),
.B(n_3659),
.Y(n_3847)
);

NAND3xp33_ASAP7_75t_L g3848 ( 
.A(n_3810),
.B(n_3701),
.C(n_3702),
.Y(n_3848)
);

BUFx2_ASAP7_75t_L g3849 ( 
.A(n_3750),
.Y(n_3849)
);

INVx1_ASAP7_75t_SL g3850 ( 
.A(n_3766),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3763),
.Y(n_3851)
);

INVx5_ASAP7_75t_L g3852 ( 
.A(n_3810),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3753),
.Y(n_3853)
);

NOR2xp33_ASAP7_75t_L g3854 ( 
.A(n_3825),
.B(n_3687),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3817),
.B(n_3692),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3817),
.B(n_3692),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3742),
.Y(n_3857)
);

INVx3_ASAP7_75t_L g3858 ( 
.A(n_3797),
.Y(n_3858)
);

BUFx2_ASAP7_75t_L g3859 ( 
.A(n_3751),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3804),
.B(n_3520),
.Y(n_3860)
);

AND2x4_ASAP7_75t_L g3861 ( 
.A(n_3742),
.B(n_3526),
.Y(n_3861)
);

AOI221xp5_ASAP7_75t_L g3862 ( 
.A1(n_3826),
.A2(n_3798),
.B1(n_3829),
.B2(n_3777),
.C(n_3761),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3804),
.B(n_3526),
.Y(n_3863)
);

OR2x2_ASAP7_75t_L g3864 ( 
.A(n_3745),
.B(n_3667),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3751),
.B(n_3514),
.Y(n_3865)
);

OAI33xp33_ASAP7_75t_L g3866 ( 
.A1(n_3813),
.A2(n_3737),
.A3(n_3700),
.B1(n_3724),
.B2(n_3719),
.B3(n_3713),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3751),
.B(n_3514),
.Y(n_3867)
);

OAI31xp33_ASAP7_75t_L g3868 ( 
.A1(n_3788),
.A2(n_3688),
.A3(n_3669),
.B(n_3663),
.Y(n_3868)
);

OR2x2_ASAP7_75t_L g3869 ( 
.A(n_3745),
.B(n_3700),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_L g3870 ( 
.A(n_3825),
.B(n_3683),
.Y(n_3870)
);

INVx2_ASAP7_75t_SL g3871 ( 
.A(n_3797),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3752),
.B(n_3514),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3802),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3802),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3752),
.Y(n_3875)
);

INVxp67_ASAP7_75t_L g3876 ( 
.A(n_3769),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3747),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3747),
.Y(n_3878)
);

INVx1_ASAP7_75t_SL g3879 ( 
.A(n_3819),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3822),
.B(n_3758),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3748),
.Y(n_3881)
);

AO21x2_ASAP7_75t_L g3882 ( 
.A1(n_3792),
.A2(n_3515),
.B(n_3713),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3748),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3773),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3789),
.B(n_3779),
.Y(n_3885)
);

NAND3xp33_ASAP7_75t_L g3886 ( 
.A(n_3759),
.B(n_3727),
.C(n_3646),
.Y(n_3886)
);

HB1xp67_ASAP7_75t_L g3887 ( 
.A(n_3792),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3773),
.Y(n_3888)
);

OR2x2_ASAP7_75t_L g3889 ( 
.A(n_3779),
.B(n_3765),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3774),
.Y(n_3890)
);

NAND4xp25_ASAP7_75t_L g3891 ( 
.A(n_3821),
.B(n_3730),
.C(n_3646),
.D(n_3715),
.Y(n_3891)
);

AND2x4_ASAP7_75t_L g3892 ( 
.A(n_3760),
.B(n_3544),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3784),
.B(n_3544),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3767),
.B(n_3546),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3797),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3774),
.Y(n_3896)
);

AND2x4_ASAP7_75t_L g3897 ( 
.A(n_3760),
.B(n_3755),
.Y(n_3897)
);

OAI31xp33_ASAP7_75t_L g3898 ( 
.A1(n_3807),
.A2(n_3830),
.A3(n_3795),
.B(n_3824),
.Y(n_3898)
);

BUFx2_ASAP7_75t_L g3899 ( 
.A(n_3760),
.Y(n_3899)
);

AOI211xp5_ASAP7_75t_SL g3900 ( 
.A1(n_3819),
.A2(n_3724),
.B(n_3719),
.C(n_3737),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3822),
.B(n_3758),
.Y(n_3901)
);

AOI211xp5_ASAP7_75t_SL g3902 ( 
.A1(n_3820),
.A2(n_3660),
.B(n_3515),
.C(n_3678),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3787),
.Y(n_3903)
);

NAND4xp25_ASAP7_75t_L g3904 ( 
.A(n_3785),
.B(n_3664),
.C(n_3618),
.D(n_3616),
.Y(n_3904)
);

OAI211xp5_ASAP7_75t_SL g3905 ( 
.A1(n_3832),
.A2(n_3616),
.B(n_3546),
.C(n_3525),
.Y(n_3905)
);

OR2x2_ASAP7_75t_L g3906 ( 
.A(n_3815),
.B(n_3524),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3787),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3830),
.A2(n_3604),
.B1(n_3541),
.B2(n_3618),
.Y(n_3908)
);

OAI31xp33_ASAP7_75t_L g3909 ( 
.A1(n_3807),
.A2(n_3604),
.A3(n_3525),
.B(n_3524),
.Y(n_3909)
);

OR2x2_ASAP7_75t_L g3910 ( 
.A(n_3815),
.B(n_3568),
.Y(n_3910)
);

HB1xp67_ASAP7_75t_L g3911 ( 
.A(n_3806),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3762),
.B(n_3806),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3793),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3762),
.B(n_3568),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_SL g3915 ( 
.A1(n_3824),
.A2(n_3541),
.B1(n_283),
.B2(n_284),
.Y(n_3915)
);

INVxp67_ASAP7_75t_L g3916 ( 
.A(n_3791),
.Y(n_3916)
);

AOI221xp5_ASAP7_75t_SL g3917 ( 
.A1(n_3795),
.A2(n_3541),
.B1(n_283),
.B2(n_285),
.C(n_286),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3744),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3755),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3746),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_3757),
.Y(n_3921)
);

AOI221x1_ASAP7_75t_L g3922 ( 
.A1(n_3757),
.A2(n_3541),
.B1(n_285),
.B2(n_286),
.C(n_287),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3793),
.B(n_282),
.Y(n_3923)
);

NOR3xp33_ASAP7_75t_L g3924 ( 
.A(n_3818),
.B(n_288),
.C(n_290),
.Y(n_3924)
);

OAI33xp33_ASAP7_75t_L g3925 ( 
.A1(n_3754),
.A2(n_3776),
.A3(n_3764),
.B1(n_3790),
.B2(n_3786),
.B3(n_3771),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3803),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3887),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3887),
.Y(n_3928)
);

HB1xp67_ASAP7_75t_L g3929 ( 
.A(n_3852),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3852),
.B(n_3767),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_L g3931 ( 
.A(n_3852),
.B(n_3803),
.Y(n_3931)
);

OR2x2_ASAP7_75t_L g3932 ( 
.A(n_3889),
.B(n_3859),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3839),
.A2(n_3805),
.B1(n_3809),
.B2(n_3818),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_3880),
.B(n_3799),
.Y(n_3934)
);

OR2x2_ASAP7_75t_L g3935 ( 
.A(n_3885),
.B(n_3749),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3911),
.Y(n_3936)
);

NAND2x1p5_ASAP7_75t_L g3937 ( 
.A(n_3852),
.B(n_3803),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3849),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3899),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3836),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3836),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3836),
.Y(n_3942)
);

OR2x2_ASAP7_75t_L g3943 ( 
.A(n_3869),
.B(n_3749),
.Y(n_3943)
);

OR2x2_ASAP7_75t_L g3944 ( 
.A(n_3842),
.B(n_3783),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3901),
.B(n_3814),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3926),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3924),
.B(n_3794),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3924),
.B(n_3778),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3919),
.Y(n_3949)
);

OR2x2_ASAP7_75t_L g3950 ( 
.A(n_3842),
.B(n_3783),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3876),
.B(n_3814),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3921),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3876),
.B(n_3780),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3840),
.Y(n_3954)
);

OR2x2_ASAP7_75t_L g3955 ( 
.A(n_3879),
.B(n_3768),
.Y(n_3955)
);

OR2x2_ASAP7_75t_L g3956 ( 
.A(n_3879),
.B(n_3768),
.Y(n_3956)
);

OAI221xp5_ASAP7_75t_L g3957 ( 
.A1(n_3868),
.A2(n_3805),
.B1(n_3811),
.B2(n_3809),
.C(n_3812),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3837),
.B(n_3799),
.Y(n_3958)
);

INVxp67_ASAP7_75t_L g3959 ( 
.A(n_3865),
.Y(n_3959)
);

HB1xp67_ASAP7_75t_L g3960 ( 
.A(n_3838),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3858),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3858),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3844),
.B(n_3775),
.Y(n_3963)
);

BUFx3_ASAP7_75t_L g3964 ( 
.A(n_3871),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3853),
.Y(n_3965)
);

INVx1_ASAP7_75t_SL g3966 ( 
.A(n_3850),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3897),
.Y(n_3967)
);

OAI21xp33_ASAP7_75t_L g3968 ( 
.A1(n_3862),
.A2(n_3811),
.B(n_3816),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3897),
.Y(n_3969)
);

AND2x4_ASAP7_75t_L g3970 ( 
.A(n_3895),
.B(n_3781),
.Y(n_3970)
);

OR2x2_ASAP7_75t_L g3971 ( 
.A(n_3855),
.B(n_3833),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3841),
.B(n_3833),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3893),
.Y(n_3973)
);

INVx2_ASAP7_75t_SL g3974 ( 
.A(n_3867),
.Y(n_3974)
);

INVxp67_ASAP7_75t_L g3975 ( 
.A(n_3835),
.Y(n_3975)
);

OR2x2_ASAP7_75t_L g3976 ( 
.A(n_3855),
.B(n_3775),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3912),
.B(n_3846),
.Y(n_3977)
);

AND2x4_ASAP7_75t_L g3978 ( 
.A(n_3843),
.B(n_3781),
.Y(n_3978)
);

OR2x2_ASAP7_75t_L g3979 ( 
.A(n_3856),
.B(n_3831),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3845),
.B(n_3782),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3863),
.B(n_3782),
.Y(n_3981)
);

NOR2xp67_ASAP7_75t_L g3982 ( 
.A(n_3848),
.B(n_3796),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3872),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3875),
.B(n_3770),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3903),
.B(n_3770),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3900),
.B(n_3823),
.Y(n_3986)
);

OR2x2_ASAP7_75t_L g3987 ( 
.A(n_3856),
.B(n_3823),
.Y(n_3987)
);

OR2x2_ASAP7_75t_L g3988 ( 
.A(n_3851),
.B(n_3827),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3862),
.A2(n_3808),
.B(n_3796),
.Y(n_3989)
);

OR2x2_ASAP7_75t_L g3990 ( 
.A(n_3857),
.B(n_3827),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3893),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3907),
.B(n_3808),
.Y(n_3992)
);

INVx3_ASAP7_75t_L g3993 ( 
.A(n_3861),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3900),
.B(n_288),
.Y(n_3994)
);

OAI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3915),
.A2(n_290),
.B(n_291),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3873),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3874),
.Y(n_3997)
);

OAI22xp5_ASAP7_75t_L g3998 ( 
.A1(n_3915),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3906),
.Y(n_3999)
);

INVx2_ASAP7_75t_SL g4000 ( 
.A(n_3834),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3860),
.Y(n_4001)
);

OR2x2_ASAP7_75t_L g4002 ( 
.A(n_3913),
.B(n_292),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3894),
.Y(n_4003)
);

HB1xp67_ASAP7_75t_L g4004 ( 
.A(n_3850),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3894),
.Y(n_4005)
);

OAI21xp33_ASAP7_75t_L g4006 ( 
.A1(n_3854),
.A2(n_293),
.B(n_294),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3923),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3861),
.B(n_295),
.Y(n_4008)
);

INVx2_ASAP7_75t_SL g4009 ( 
.A(n_3834),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3916),
.B(n_295),
.Y(n_4010)
);

AOI33xp33_ASAP7_75t_L g4011 ( 
.A1(n_3908),
.A2(n_296),
.A3(n_297),
.B1(n_298),
.B2(n_299),
.B3(n_300),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3841),
.B(n_296),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3898),
.B(n_297),
.Y(n_4013)
);

OR2x2_ASAP7_75t_L g4014 ( 
.A(n_3904),
.B(n_300),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3892),
.Y(n_4015)
);

BUFx2_ASAP7_75t_L g4016 ( 
.A(n_3892),
.Y(n_4016)
);

INVx1_ASAP7_75t_SL g4017 ( 
.A(n_3882),
.Y(n_4017)
);

NOR2xp33_ASAP7_75t_L g4018 ( 
.A(n_3966),
.B(n_3916),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3927),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3928),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3946),
.B(n_3870),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3966),
.B(n_3917),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3958),
.B(n_3934),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3964),
.B(n_3917),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_4004),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3937),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3963),
.B(n_3914),
.Y(n_4027)
);

INVxp67_ASAP7_75t_L g4028 ( 
.A(n_4016),
.Y(n_4028)
);

INVxp67_ASAP7_75t_L g4029 ( 
.A(n_3960),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3932),
.B(n_3866),
.Y(n_4030)
);

NOR3x1_ASAP7_75t_L g4031 ( 
.A(n_3957),
.B(n_3886),
.C(n_3891),
.Y(n_4031)
);

BUFx2_ASAP7_75t_L g4032 ( 
.A(n_3993),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3955),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_4017),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3977),
.B(n_4000),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_4009),
.B(n_3882),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3961),
.B(n_3910),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_3962),
.B(n_3864),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3993),
.B(n_3847),
.Y(n_4039)
);

O2A1O1Ixp33_ASAP7_75t_L g4040 ( 
.A1(n_3995),
.A2(n_3902),
.B(n_3866),
.C(n_3905),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3970),
.B(n_3978),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3956),
.Y(n_4042)
);

BUFx3_ASAP7_75t_L g4043 ( 
.A(n_3942),
.Y(n_4043)
);

INVx3_ASAP7_75t_L g4044 ( 
.A(n_4017),
.Y(n_4044)
);

OR2x4_ASAP7_75t_L g4045 ( 
.A(n_3938),
.B(n_3918),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3929),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3968),
.A2(n_3905),
.B1(n_3909),
.B2(n_3925),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3969),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3981),
.B(n_3902),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3970),
.B(n_3922),
.Y(n_4050)
);

NOR3xp33_ASAP7_75t_L g4051 ( 
.A(n_3968),
.B(n_3925),
.C(n_3920),
.Y(n_4051)
);

AOI31xp33_ASAP7_75t_L g4052 ( 
.A1(n_3995),
.A2(n_3896),
.A3(n_3890),
.B(n_3888),
.Y(n_4052)
);

INVx3_ASAP7_75t_L g4053 ( 
.A(n_3978),
.Y(n_4053)
);

INVx2_ASAP7_75t_SL g4054 ( 
.A(n_3967),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3984),
.B(n_3877),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3939),
.Y(n_4056)
);

AND2x4_ASAP7_75t_L g4057 ( 
.A(n_4015),
.B(n_3878),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3992),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3985),
.B(n_3881),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3940),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3936),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3941),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3975),
.B(n_3883),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_4001),
.B(n_3884),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3974),
.B(n_301),
.Y(n_4065)
);

BUFx2_ASAP7_75t_SL g4066 ( 
.A(n_3949),
.Y(n_4066)
);

INVx1_ASAP7_75t_SL g4067 ( 
.A(n_3943),
.Y(n_4067)
);

BUFx3_ASAP7_75t_L g4068 ( 
.A(n_3931),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3944),
.Y(n_4069)
);

NAND2x1p5_ASAP7_75t_L g4070 ( 
.A(n_4008),
.B(n_302),
.Y(n_4070)
);

INVxp67_ASAP7_75t_L g4071 ( 
.A(n_3951),
.Y(n_4071)
);

OAI33xp33_ASAP7_75t_L g4072 ( 
.A1(n_3933),
.A2(n_303),
.A3(n_304),
.B1(n_305),
.B2(n_306),
.B3(n_307),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3950),
.Y(n_4073)
);

INVx3_ASAP7_75t_L g4074 ( 
.A(n_3990),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3983),
.B(n_303),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3952),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3998),
.B(n_305),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3930),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_4007),
.B(n_308),
.Y(n_4079)
);

INVx3_ASAP7_75t_L g4080 ( 
.A(n_3988),
.Y(n_4080)
);

HB1xp67_ASAP7_75t_L g4081 ( 
.A(n_3982),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_3959),
.B(n_309),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3945),
.B(n_309),
.Y(n_4083)
);

AND2x4_ASAP7_75t_L g4084 ( 
.A(n_3982),
.B(n_310),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3999),
.B(n_310),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3998),
.B(n_4010),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3976),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_3971),
.B(n_311),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_4011),
.B(n_312),
.Y(n_4089)
);

INVx2_ASAP7_75t_SL g4090 ( 
.A(n_4002),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3953),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_3954),
.B(n_312),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3935),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3965),
.B(n_313),
.Y(n_4094)
);

OR2x2_ASAP7_75t_L g4095 ( 
.A(n_3987),
.B(n_313),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_4006),
.B(n_3986),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3980),
.B(n_314),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3953),
.Y(n_4098)
);

AND4x1_ASAP7_75t_L g4099 ( 
.A(n_4006),
.B(n_314),
.C(n_315),
.D(n_316),
.Y(n_4099)
);

OR2x2_ASAP7_75t_L g4100 ( 
.A(n_3972),
.B(n_3979),
.Y(n_4100)
);

NAND2x1_ASAP7_75t_L g4101 ( 
.A(n_3996),
.B(n_315),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3989),
.B(n_316),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_4035),
.B(n_3973),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_4081),
.B(n_3994),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4035),
.B(n_3991),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_L g4106 ( 
.A1(n_4051),
.A2(n_3933),
.B1(n_4013),
.B2(n_3972),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_4044),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_4053),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4053),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_4030),
.A2(n_4014),
.B1(n_4012),
.B2(n_3948),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4053),
.Y(n_4111)
);

OR2x2_ASAP7_75t_L g4112 ( 
.A(n_4050),
.B(n_3947),
.Y(n_4112)
);

HB1xp67_ASAP7_75t_L g4113 ( 
.A(n_4081),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4036),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4036),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_4032),
.Y(n_4116)
);

OR2x2_ASAP7_75t_L g4117 ( 
.A(n_4067),
.B(n_3947),
.Y(n_4117)
);

OR2x2_ASAP7_75t_L g4118 ( 
.A(n_4024),
.B(n_3948),
.Y(n_4118)
);

AND2x4_ASAP7_75t_L g4119 ( 
.A(n_4074),
.B(n_3997),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_4023),
.B(n_4003),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4027),
.B(n_4005),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_4044),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_4037),
.B(n_4012),
.Y(n_4123)
);

NOR2xp67_ASAP7_75t_SL g4124 ( 
.A(n_4066),
.B(n_317),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4044),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_4084),
.Y(n_4126)
);

INVx1_ASAP7_75t_SL g4127 ( 
.A(n_4041),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4037),
.B(n_319),
.Y(n_4128)
);

OR2x2_ASAP7_75t_L g4129 ( 
.A(n_4054),
.B(n_319),
.Y(n_4129)
);

INVx2_ASAP7_75t_SL g4130 ( 
.A(n_4057),
.Y(n_4130)
);

OR2x2_ASAP7_75t_L g4131 ( 
.A(n_4054),
.B(n_320),
.Y(n_4131)
);

HB1xp67_ASAP7_75t_L g4132 ( 
.A(n_4101),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_4049),
.B(n_320),
.Y(n_4133)
);

HB1xp67_ASAP7_75t_L g4134 ( 
.A(n_4074),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_4028),
.B(n_321),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_4043),
.B(n_322),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4043),
.B(n_323),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_4038),
.B(n_4068),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4074),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4080),
.Y(n_4140)
);

NOR2x1_ASAP7_75t_L g4141 ( 
.A(n_4084),
.B(n_323),
.Y(n_4141)
);

OAI22xp5_ASAP7_75t_L g4142 ( 
.A1(n_4047),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4080),
.Y(n_4143)
);

OR2x2_ASAP7_75t_L g4144 ( 
.A(n_4022),
.B(n_324),
.Y(n_4144)
);

NAND3xp33_ASAP7_75t_L g4145 ( 
.A(n_4047),
.B(n_325),
.C(n_326),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_4038),
.B(n_327),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4049),
.B(n_329),
.Y(n_4147)
);

INVx1_ASAP7_75t_SL g4148 ( 
.A(n_4068),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_4048),
.B(n_329),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4048),
.B(n_330),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4093),
.B(n_331),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4093),
.B(n_331),
.Y(n_4152)
);

BUFx2_ASAP7_75t_L g4153 ( 
.A(n_4080),
.Y(n_4153)
);

OAI22xp5_ASAP7_75t_L g4154 ( 
.A1(n_4040),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_4154)
);

OAI32xp33_ASAP7_75t_L g4155 ( 
.A1(n_4030),
.A2(n_332),
.A3(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4057),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_4087),
.B(n_338),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_4029),
.B(n_338),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_4084),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4018),
.B(n_339),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4087),
.B(n_340),
.Y(n_4161)
);

INVx2_ASAP7_75t_SL g4162 ( 
.A(n_4057),
.Y(n_4162)
);

NAND2x1p5_ASAP7_75t_L g4163 ( 
.A(n_4025),
.B(n_340),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4018),
.B(n_341),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4046),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4055),
.Y(n_4166)
);

HB1xp67_ASAP7_75t_L g4167 ( 
.A(n_4070),
.Y(n_4167)
);

INVx1_ASAP7_75t_SL g4168 ( 
.A(n_4059),
.Y(n_4168)
);

OR2x2_ASAP7_75t_L g4169 ( 
.A(n_4039),
.B(n_4086),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4033),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_4153),
.B(n_4130),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4130),
.B(n_4162),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_4162),
.B(n_4102),
.Y(n_4173)
);

NOR3xp33_ASAP7_75t_L g4174 ( 
.A(n_4142),
.B(n_4021),
.C(n_4096),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_4148),
.B(n_4052),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4134),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_4138),
.B(n_4042),
.Y(n_4177)
);

AOI22xp33_ASAP7_75t_L g4178 ( 
.A1(n_4145),
.A2(n_4073),
.B1(n_4069),
.B2(n_4056),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4113),
.Y(n_4179)
);

NOR2xp33_ASAP7_75t_L g4180 ( 
.A(n_4132),
.B(n_4167),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4107),
.Y(n_4181)
);

AOI32xp33_ASAP7_75t_L g4182 ( 
.A1(n_4106),
.A2(n_4154),
.A3(n_4110),
.B1(n_4138),
.B2(n_4104),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4124),
.B(n_4026),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4156),
.Y(n_4184)
);

AND2x2_ASAP7_75t_L g4185 ( 
.A(n_4120),
.B(n_4121),
.Y(n_4185)
);

NOR2x1_ASAP7_75t_L g4186 ( 
.A(n_4141),
.B(n_4100),
.Y(n_4186)
);

INVxp67_ASAP7_75t_L g4187 ( 
.A(n_4104),
.Y(n_4187)
);

AOI211x1_ASAP7_75t_L g4188 ( 
.A1(n_4155),
.A2(n_4058),
.B(n_4099),
.C(n_4019),
.Y(n_4188)
);

AOI21x1_ASAP7_75t_L g4189 ( 
.A1(n_4119),
.A2(n_4034),
.B(n_4026),
.Y(n_4189)
);

INVx2_ASAP7_75t_SL g4190 ( 
.A(n_4119),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_4103),
.B(n_4078),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4107),
.Y(n_4192)
);

NOR2xp33_ASAP7_75t_L g4193 ( 
.A(n_4127),
.B(n_4071),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4122),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4122),
.Y(n_4195)
);

NAND3xp33_ASAP7_75t_L g4196 ( 
.A(n_4106),
.B(n_4061),
.C(n_4076),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_4116),
.B(n_4088),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_4120),
.B(n_4083),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_SL g4199 ( 
.A(n_4126),
.B(n_4090),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4103),
.B(n_4078),
.Y(n_4200)
);

NAND3xp33_ASAP7_75t_L g4201 ( 
.A(n_4110),
.B(n_4060),
.C(n_4062),
.Y(n_4201)
);

HB1xp67_ASAP7_75t_L g4202 ( 
.A(n_4119),
.Y(n_4202)
);

INVxp67_ASAP7_75t_L g4203 ( 
.A(n_4105),
.Y(n_4203)
);

NOR2x2_ASAP7_75t_L g4204 ( 
.A(n_4126),
.B(n_4060),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4105),
.B(n_4097),
.Y(n_4205)
);

OR2x2_ASAP7_75t_L g4206 ( 
.A(n_4112),
.B(n_4090),
.Y(n_4206)
);

OR2x2_ASAP7_75t_L g4207 ( 
.A(n_4168),
.B(n_4095),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4159),
.B(n_4085),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4139),
.Y(n_4209)
);

OAI21xp33_ASAP7_75t_L g4210 ( 
.A1(n_4169),
.A2(n_4063),
.B(n_4062),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_4117),
.B(n_4072),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4159),
.B(n_4085),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4140),
.B(n_4031),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_4143),
.B(n_4075),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4108),
.Y(n_4215)
);

BUFx3_ASAP7_75t_L g4216 ( 
.A(n_4163),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4121),
.B(n_4166),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4109),
.Y(n_4218)
);

AOI221xp5_ASAP7_75t_L g4219 ( 
.A1(n_4133),
.A2(n_4098),
.B1(n_4091),
.B2(n_4034),
.C(n_4020),
.Y(n_4219)
);

NOR2xp67_ASAP7_75t_L g4220 ( 
.A(n_4125),
.B(n_4064),
.Y(n_4220)
);

NAND2x1p5_ASAP7_75t_L g4221 ( 
.A(n_4111),
.B(n_4075),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4123),
.B(n_4082),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4114),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_4128),
.B(n_4092),
.Y(n_4224)
);

A2O1A1Ixp33_ASAP7_75t_L g4225 ( 
.A1(n_4158),
.A2(n_4077),
.B(n_4089),
.C(n_4092),
.Y(n_4225)
);

OR2x2_ASAP7_75t_L g4226 ( 
.A(n_4147),
.B(n_4065),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4123),
.B(n_4064),
.Y(n_4227)
);

AOI22xp33_ASAP7_75t_L g4228 ( 
.A1(n_4118),
.A2(n_4079),
.B1(n_4094),
.B2(n_4070),
.Y(n_4228)
);

NAND3xp33_ASAP7_75t_L g4229 ( 
.A(n_4165),
.B(n_4094),
.C(n_4045),
.Y(n_4229)
);

NAND2x1_ASAP7_75t_L g4230 ( 
.A(n_4136),
.B(n_4045),
.Y(n_4230)
);

AND2x2_ASAP7_75t_L g4231 ( 
.A(n_4146),
.B(n_341),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4115),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4128),
.B(n_342),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4185),
.B(n_4190),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4202),
.Y(n_4235)
);

OAI32xp33_ASAP7_75t_L g4236 ( 
.A1(n_4213),
.A2(n_4144),
.A3(n_4170),
.B1(n_4164),
.B2(n_4160),
.Y(n_4236)
);

OAI21xp33_ASAP7_75t_L g4237 ( 
.A1(n_4213),
.A2(n_4158),
.B(n_4152),
.Y(n_4237)
);

OAI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_4196),
.A2(n_4186),
.B(n_4201),
.Y(n_4238)
);

AO22x2_ASAP7_75t_L g4239 ( 
.A1(n_4230),
.A2(n_4129),
.B1(n_4131),
.B2(n_4151),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4189),
.Y(n_4240)
);

AOI21xp33_ASAP7_75t_L g4241 ( 
.A1(n_4180),
.A2(n_4152),
.B(n_4151),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4174),
.A2(n_4146),
.B1(n_4135),
.B2(n_4157),
.Y(n_4242)
);

AO221x1_ASAP7_75t_L g4243 ( 
.A1(n_4203),
.A2(n_4163),
.B1(n_4135),
.B2(n_4157),
.C(n_4161),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_4216),
.B(n_4136),
.Y(n_4244)
);

OAI21xp33_ASAP7_75t_SL g4245 ( 
.A1(n_4182),
.A2(n_4161),
.B(n_4137),
.Y(n_4245)
);

AOI222xp33_ASAP7_75t_L g4246 ( 
.A1(n_4211),
.A2(n_4150),
.B1(n_4149),
.B2(n_4137),
.C1(n_347),
.C2(n_349),
.Y(n_4246)
);

OAI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_4183),
.A2(n_4149),
.B1(n_4150),
.B2(n_346),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4198),
.B(n_344),
.Y(n_4248)
);

INVxp67_ASAP7_75t_L g4249 ( 
.A(n_4171),
.Y(n_4249)
);

NOR2xp33_ASAP7_75t_L g4250 ( 
.A(n_4224),
.B(n_345),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4171),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4172),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4222),
.B(n_4217),
.Y(n_4253)
);

AND2x2_ASAP7_75t_L g4254 ( 
.A(n_4227),
.B(n_349),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_4220),
.B(n_350),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4172),
.Y(n_4256)
);

INVxp67_ASAP7_75t_L g4257 ( 
.A(n_4199),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4228),
.B(n_350),
.Y(n_4258)
);

INVxp67_ASAP7_75t_L g4259 ( 
.A(n_4191),
.Y(n_4259)
);

AOI211xp5_ASAP7_75t_L g4260 ( 
.A1(n_4175),
.A2(n_352),
.B(n_353),
.C(n_354),
.Y(n_4260)
);

AOI211xp5_ASAP7_75t_L g4261 ( 
.A1(n_4210),
.A2(n_352),
.B(n_353),
.C(n_355),
.Y(n_4261)
);

OAI21xp33_ASAP7_75t_L g4262 ( 
.A1(n_4193),
.A2(n_355),
.B(n_356),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4221),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4221),
.Y(n_4264)
);

AOI21xp33_ASAP7_75t_SL g4265 ( 
.A1(n_4206),
.A2(n_356),
.B(n_357),
.Y(n_4265)
);

AOI222xp33_ASAP7_75t_L g4266 ( 
.A1(n_4229),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.C1(n_362),
.C2(n_364),
.Y(n_4266)
);

NAND4xp25_ASAP7_75t_L g4267 ( 
.A(n_4188),
.B(n_359),
.C(n_364),
.D(n_393),
.Y(n_4267)
);

OAI21xp33_ASAP7_75t_L g4268 ( 
.A1(n_4178),
.A2(n_4177),
.B(n_4205),
.Y(n_4268)
);

OAI221xp5_ASAP7_75t_SL g4269 ( 
.A1(n_4187),
.A2(n_394),
.B1(n_396),
.B2(n_399),
.C(n_401),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4204),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4224),
.Y(n_4271)
);

AOI222xp33_ASAP7_75t_L g4272 ( 
.A1(n_4219),
.A2(n_402),
.B1(n_411),
.B2(n_413),
.C1(n_414),
.C2(n_419),
.Y(n_4272)
);

AOI22xp5_ASAP7_75t_L g4273 ( 
.A1(n_4176),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_4273)
);

INVx3_ASAP7_75t_L g4274 ( 
.A(n_4181),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4179),
.B(n_425),
.Y(n_4275)
);

OR2x2_ASAP7_75t_L g4276 ( 
.A(n_4200),
.B(n_435),
.Y(n_4276)
);

OAI21xp33_ASAP7_75t_L g4277 ( 
.A1(n_4225),
.A2(n_436),
.B(n_439),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_4207),
.B(n_1261),
.Y(n_4278)
);

OAI22xp33_ASAP7_75t_L g4279 ( 
.A1(n_4208),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4212),
.Y(n_4280)
);

AO221x1_ASAP7_75t_L g4281 ( 
.A1(n_4184),
.A2(n_444),
.B1(n_446),
.B2(n_448),
.C(n_449),
.Y(n_4281)
);

OAI22xp33_ASAP7_75t_L g4282 ( 
.A1(n_4197),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_4282)
);

O2A1O1Ixp33_ASAP7_75t_L g4283 ( 
.A1(n_4173),
.A2(n_454),
.B(n_455),
.C(n_457),
.Y(n_4283)
);

OAI22xp33_ASAP7_75t_L g4284 ( 
.A1(n_4173),
.A2(n_462),
.B1(n_463),
.B2(n_466),
.Y(n_4284)
);

AOI21xp33_ASAP7_75t_L g4285 ( 
.A1(n_4238),
.A2(n_4214),
.B(n_4195),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4239),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4240),
.B(n_4194),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_SL g4288 ( 
.A(n_4245),
.B(n_4257),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4239),
.Y(n_4289)
);

AOI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_4253),
.A2(n_4215),
.B1(n_4218),
.B2(n_4209),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4234),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4235),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4274),
.Y(n_4293)
);

AOI211xp5_ASAP7_75t_L g4294 ( 
.A1(n_4241),
.A2(n_4214),
.B(n_4192),
.C(n_4223),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_4274),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4254),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4243),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_4270),
.B(n_4263),
.Y(n_4298)
);

OR2x2_ASAP7_75t_L g4299 ( 
.A(n_4264),
.B(n_4226),
.Y(n_4299)
);

AND2x2_ASAP7_75t_L g4300 ( 
.A(n_4242),
.B(n_4231),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4248),
.B(n_4232),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_SL g4302 ( 
.A(n_4245),
.B(n_4233),
.Y(n_4302)
);

OAI22xp33_ASAP7_75t_L g4303 ( 
.A1(n_4267),
.A2(n_467),
.B1(n_469),
.B2(n_471),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4258),
.B(n_473),
.Y(n_4304)
);

OR2x2_ASAP7_75t_L g4305 ( 
.A(n_4244),
.B(n_474),
.Y(n_4305)
);

CKINVDCx20_ASAP7_75t_R g4306 ( 
.A(n_4249),
.Y(n_4306)
);

INVx3_ASAP7_75t_L g4307 ( 
.A(n_4252),
.Y(n_4307)
);

AOI21xp33_ASAP7_75t_L g4308 ( 
.A1(n_4246),
.A2(n_477),
.B(n_480),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_L g4309 ( 
.A(n_4237),
.B(n_484),
.Y(n_4309)
);

INVx2_ASAP7_75t_SL g4310 ( 
.A(n_4256),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4265),
.B(n_485),
.Y(n_4311)
);

AOI21xp33_ASAP7_75t_L g4312 ( 
.A1(n_4247),
.A2(n_486),
.B(n_487),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4255),
.Y(n_4313)
);

INVxp67_ASAP7_75t_L g4314 ( 
.A(n_4250),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4251),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4271),
.B(n_488),
.Y(n_4316)
);

NOR2xp33_ASAP7_75t_SL g4317 ( 
.A(n_4268),
.B(n_489),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4280),
.Y(n_4318)
);

OAI31xp33_ASAP7_75t_L g4319 ( 
.A1(n_4259),
.A2(n_491),
.A3(n_496),
.B(n_498),
.Y(n_4319)
);

INVx2_ASAP7_75t_SL g4320 ( 
.A(n_4281),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4276),
.Y(n_4321)
);

OR2x2_ASAP7_75t_L g4322 ( 
.A(n_4275),
.B(n_499),
.Y(n_4322)
);

OAI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4288),
.A2(n_4260),
.B(n_4266),
.Y(n_4323)
);

NOR2xp33_ASAP7_75t_L g4324 ( 
.A(n_4302),
.B(n_4262),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4286),
.B(n_4261),
.Y(n_4325)
);

INVx1_ASAP7_75t_SL g4326 ( 
.A(n_4298),
.Y(n_4326)
);

AND2x2_ASAP7_75t_L g4327 ( 
.A(n_4300),
.B(n_4236),
.Y(n_4327)
);

AOI21xp5_ASAP7_75t_L g4328 ( 
.A1(n_4285),
.A2(n_4277),
.B(n_4278),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4289),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4287),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4296),
.B(n_4272),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4287),
.Y(n_4332)
);

O2A1O1Ixp33_ASAP7_75t_L g4333 ( 
.A1(n_4285),
.A2(n_4283),
.B(n_4284),
.C(n_4279),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4301),
.Y(n_4334)
);

AOI22xp33_ASAP7_75t_SL g4335 ( 
.A1(n_4306),
.A2(n_4317),
.B1(n_4292),
.B2(n_4297),
.Y(n_4335)
);

OR2x2_ASAP7_75t_L g4336 ( 
.A(n_4301),
.B(n_4299),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4293),
.B(n_4282),
.Y(n_4337)
);

OAI221xp5_ASAP7_75t_SL g4338 ( 
.A1(n_4290),
.A2(n_4273),
.B1(n_4269),
.B2(n_504),
.C(n_506),
.Y(n_4338)
);

INVxp67_ASAP7_75t_L g4339 ( 
.A(n_4317),
.Y(n_4339)
);

INVx1_ASAP7_75t_SL g4340 ( 
.A(n_4295),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4307),
.Y(n_4341)
);

AOI221xp5_ASAP7_75t_L g4342 ( 
.A1(n_4308),
.A2(n_4273),
.B1(n_503),
.B2(n_507),
.C(n_508),
.Y(n_4342)
);

AOI21xp33_ASAP7_75t_L g4343 ( 
.A1(n_4291),
.A2(n_500),
.B(n_1230),
.Y(n_4343)
);

INVxp67_ASAP7_75t_SL g4344 ( 
.A(n_4307),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4320),
.B(n_1290),
.Y(n_4345)
);

AOI221xp5_ASAP7_75t_L g4346 ( 
.A1(n_4308),
.A2(n_1236),
.B1(n_1261),
.B2(n_1256),
.C(n_1159),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_4310),
.B(n_1159),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4327),
.B(n_4304),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4344),
.Y(n_4349)
);

AOI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4326),
.A2(n_4303),
.B1(n_4314),
.B2(n_4309),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_L g4351 ( 
.A1(n_4329),
.A2(n_4321),
.B1(n_4313),
.B2(n_4318),
.Y(n_4351)
);

XNOR2x1_ASAP7_75t_L g4352 ( 
.A(n_4336),
.B(n_4305),
.Y(n_4352)
);

AOI221xp5_ASAP7_75t_L g4353 ( 
.A1(n_4340),
.A2(n_4315),
.B1(n_4294),
.B2(n_4312),
.C(n_4316),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4341),
.Y(n_4354)
);

XNOR2x1_ASAP7_75t_L g4355 ( 
.A(n_4323),
.B(n_4322),
.Y(n_4355)
);

XOR2x2_ASAP7_75t_L g4356 ( 
.A(n_4324),
.B(n_4311),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4340),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4335),
.B(n_4311),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4339),
.B(n_4312),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4334),
.Y(n_4360)
);

NAND2x1_ASAP7_75t_L g4361 ( 
.A(n_4330),
.B(n_4319),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_4332),
.B(n_1290),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_4325),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4357),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4348),
.B(n_4345),
.Y(n_4365)
);

NAND4xp75_ASAP7_75t_L g4366 ( 
.A(n_4353),
.B(n_4337),
.C(n_4328),
.D(n_4331),
.Y(n_4366)
);

NAND2x1_ASAP7_75t_SL g4367 ( 
.A(n_4349),
.B(n_4347),
.Y(n_4367)
);

NOR3xp33_ASAP7_75t_L g4368 ( 
.A(n_4363),
.B(n_4333),
.C(n_4338),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_4354),
.B(n_4342),
.Y(n_4369)
);

NOR3xp33_ASAP7_75t_L g4370 ( 
.A(n_4358),
.B(n_4343),
.C(n_4346),
.Y(n_4370)
);

NOR2x1_ASAP7_75t_L g4371 ( 
.A(n_4352),
.B(n_1236),
.Y(n_4371)
);

NOR2x1_ASAP7_75t_L g4372 ( 
.A(n_4361),
.B(n_1236),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4356),
.Y(n_4373)
);

NAND4xp75_ASAP7_75t_L g4374 ( 
.A(n_4359),
.B(n_1236),
.C(n_1261),
.D(n_1256),
.Y(n_4374)
);

NOR2xp67_ASAP7_75t_L g4375 ( 
.A(n_4364),
.B(n_4350),
.Y(n_4375)
);

OA22x2_ASAP7_75t_L g4376 ( 
.A1(n_4373),
.A2(n_4361),
.B1(n_4360),
.B2(n_4362),
.Y(n_4376)
);

NAND4xp75_ASAP7_75t_L g4377 ( 
.A(n_4372),
.B(n_4355),
.C(n_4351),
.D(n_1256),
.Y(n_4377)
);

AOI222xp33_ASAP7_75t_L g4378 ( 
.A1(n_4365),
.A2(n_1236),
.B1(n_1261),
.B2(n_1256),
.C1(n_1290),
.C2(n_1286),
.Y(n_4378)
);

AOI221xp5_ASAP7_75t_SL g4379 ( 
.A1(n_4369),
.A2(n_1256),
.B1(n_1261),
.B2(n_1159),
.C(n_1290),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4366),
.Y(n_4380)
);

A2O1A1Ixp33_ASAP7_75t_L g4381 ( 
.A1(n_4368),
.A2(n_1286),
.B(n_1275),
.C(n_1271),
.Y(n_4381)
);

NOR4xp75_ASAP7_75t_L g4382 ( 
.A(n_4377),
.B(n_4367),
.C(n_4374),
.D(n_4370),
.Y(n_4382)
);

NOR2x1_ASAP7_75t_L g4383 ( 
.A(n_4375),
.B(n_4371),
.Y(n_4383)
);

NOR2x1_ASAP7_75t_L g4384 ( 
.A(n_4380),
.B(n_1290),
.Y(n_4384)
);

AND2x2_ASAP7_75t_L g4385 ( 
.A(n_4376),
.B(n_1286),
.Y(n_4385)
);

NAND3x1_ASAP7_75t_SL g4386 ( 
.A(n_4381),
.B(n_1286),
.C(n_1275),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_SL g4387 ( 
.A1(n_4385),
.A2(n_4379),
.B1(n_4378),
.B2(n_1271),
.Y(n_4387)
);

AOI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_4383),
.A2(n_1286),
.B(n_1275),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4387),
.Y(n_4389)
);

OAI311xp33_ASAP7_75t_L g4390 ( 
.A1(n_4388),
.A2(n_4382),
.A3(n_4386),
.B1(n_4384),
.C1(n_1271),
.Y(n_4390)
);

OAI221xp5_ASAP7_75t_L g4391 ( 
.A1(n_4389),
.A2(n_1271),
.B1(n_1275),
.B2(n_997),
.C(n_1053),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4391),
.Y(n_4392)
);

AND2x4_ASAP7_75t_L g4393 ( 
.A(n_4392),
.B(n_4390),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4393),
.B(n_1271),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4394),
.Y(n_4395)
);

OAI22xp5_ASAP7_75t_SL g4396 ( 
.A1(n_4395),
.A2(n_1275),
.B1(n_997),
.B2(n_1019),
.Y(n_4396)
);

OAI22xp5_ASAP7_75t_SL g4397 ( 
.A1(n_4396),
.A2(n_997),
.B1(n_1013),
.B2(n_1019),
.Y(n_4397)
);

OAI22xp33_ASAP7_75t_SL g4398 ( 
.A1(n_4397),
.A2(n_997),
.B1(n_1013),
.B2(n_1019),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4398),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_4399),
.B(n_1013),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4400),
.Y(n_4401)
);

OAI22xp33_ASAP7_75t_L g4402 ( 
.A1(n_4400),
.A2(n_1013),
.B1(n_1019),
.B2(n_1016),
.Y(n_4402)
);

OR2x6_ASAP7_75t_L g4403 ( 
.A(n_4401),
.B(n_1053),
.Y(n_4403)
);

AOI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4403),
.A2(n_4402),
.B(n_1053),
.Y(n_4404)
);

AOI211xp5_ASAP7_75t_L g4405 ( 
.A1(n_4404),
.A2(n_1013),
.B(n_1019),
.C(n_4380),
.Y(n_4405)
);


endmodule