module fake_jpeg_16851_n_354 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_70),
.B1(n_74),
.B2(n_40),
.Y(n_76)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_40),
.B1(n_17),
.B2(n_48),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_62),
.B1(n_73),
.B2(n_37),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_29),
.B1(n_35),
.B2(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_71),
.Y(n_80)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_24),
.B1(n_32),
.B2(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_32),
.B1(n_24),
.B2(n_33),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_47),
.B1(n_45),
.B2(n_39),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_55),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_48),
.B1(n_38),
.B2(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_47),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_96),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_98),
.B1(n_54),
.B2(n_64),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_100),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_37),
.Y(n_96)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_60),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_57),
.C(n_71),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_115),
.C(n_120),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_106),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_65),
.B1(n_67),
.B2(n_56),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_127),
.B1(n_89),
.B2(n_69),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_37),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_116),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_58),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_30),
.B(n_46),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_121),
.B(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_88),
.B1(n_91),
.B2(n_81),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_46),
.C(n_42),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_46),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_20),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_130),
.C(n_44),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_68),
.B1(n_64),
.B2(n_54),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_46),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_44),
.C(n_42),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_128),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_135),
.B1(n_107),
.B2(n_137),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_139),
.A2(n_143),
.B1(n_152),
.B2(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_144),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_88),
.B1(n_43),
.B2(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_89),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_18),
.B(n_21),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_20),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_159),
.C(n_118),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_105),
.B1(n_107),
.B2(n_130),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_113),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_156),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_129),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_75),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_36),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_27),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_43),
.B1(n_17),
.B2(n_51),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_163),
.B1(n_114),
.B2(n_25),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_36),
.C(n_33),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_25),
.B1(n_33),
.B2(n_15),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_168),
.B(n_172),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_173),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_177),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_120),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_183),
.C(n_79),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_110),
.B(n_122),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_188),
.B(n_19),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_119),
.B1(n_127),
.B2(n_132),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_194),
.B1(n_158),
.B2(n_149),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_27),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_131),
.B1(n_117),
.B2(n_18),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_180),
.B(n_190),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_163),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_97),
.C(n_79),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_191),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_18),
.B(n_21),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_51),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_97),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_0),
.B(n_2),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g194 ( 
.A1(n_147),
.A2(n_154),
.B1(n_155),
.B2(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_195),
.B(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_R g198 ( 
.A(n_181),
.B(n_134),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_198),
.A2(n_193),
.B(n_22),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_199),
.A2(n_202),
.B1(n_210),
.B2(n_215),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_209),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_159),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_212),
.C(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_138),
.B1(n_131),
.B2(n_94),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_94),
.B1(n_90),
.B2(n_97),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_90),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_27),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_223),
.C(n_22),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_178),
.C(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_164),
.B1(n_191),
.B2(n_168),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_194),
.B1(n_175),
.B2(n_187),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_194),
.B1(n_174),
.B2(n_180),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_170),
.B1(n_173),
.B2(n_188),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_170),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_244),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_199),
.B(n_198),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_247),
.B1(n_249),
.B2(n_197),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_246),
.C(n_210),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_79),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_28),
.C(n_22),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_202),
.A2(n_28),
.B1(n_22),
.B2(n_19),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_28),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_253),
.B(n_261),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_262),
.C(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_216),
.C(n_222),
.Y(n_262)
);

INVxp33_ASAP7_75t_SL g263 ( 
.A(n_225),
.Y(n_263)
);

AO221x1_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_249),
.B1(n_250),
.B2(n_238),
.C(n_5),
.Y(n_291)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_218),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_218),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_231),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_214),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_28),
.C(n_19),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_252),
.B(n_8),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_19),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_245),
.B(n_8),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_2),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_268),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_235),
.B(n_251),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_260),
.B(n_259),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_243),
.C(n_246),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_283),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_242),
.C(n_234),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_238),
.C(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_8),
.B(n_13),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_10),
.B(n_15),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_295),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_302),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_269),
.B(n_254),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_304),
.B(n_284),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_269),
.B1(n_270),
.B2(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_303),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_259),
.B(n_276),
.Y(n_303)
);

OAI21x1_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_282),
.B(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_260),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_278),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_320),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_277),
.C(n_280),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_322),
.C(n_325),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_317),
.B(n_296),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_299),
.B(n_298),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_285),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_287),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_277),
.C(n_288),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_323),
.A2(n_7),
.B(n_11),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_309),
.B(n_301),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_307),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_2),
.C(n_3),
.Y(n_325)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_329),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_330),
.B(n_316),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_333),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_305),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_7),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

OA21x2_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_320),
.B(n_312),
.Y(n_338)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_342),
.B(n_12),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_325),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_339),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_10),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_331),
.C(n_4),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_345),
.A2(n_348),
.B(n_3),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_12),
.C(n_5),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_346),
.A2(n_339),
.B(n_337),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_350),
.C(n_347),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_341),
.Y(n_352)
);

AOI32xp33_ASAP7_75t_SL g353 ( 
.A1(n_352),
.A2(n_5),
.A3(n_6),
.B1(n_344),
.B2(n_348),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_5),
.Y(n_354)
);


endmodule