module fake_jpeg_5430_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_41),
.B1(n_21),
.B2(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_59),
.B1(n_66),
.B2(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_57),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_34),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_31),
.Y(n_83)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_49),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_46),
.B(n_38),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_86),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_62),
.B(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_41),
.B1(n_28),
.B2(n_29),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_59),
.B1(n_28),
.B2(n_29),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

NOR2x1_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_56),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_94),
.B(n_97),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_96),
.B1(n_103),
.B2(n_104),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_62),
.B(n_36),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_42),
.B1(n_54),
.B2(n_36),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_100),
.B(n_107),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_101),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_42),
.B(n_51),
.C(n_30),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_30),
.B1(n_51),
.B2(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_30),
.B1(n_51),
.B2(n_63),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_30),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_80),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_40),
.B(n_32),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_26),
.B(n_15),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_25),
.B1(n_26),
.B2(n_19),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_68),
.C(n_35),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_74),
.C(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_115),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_126),
.C(n_109),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_127),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_80),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_95),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_124),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_57),
.B1(n_68),
.B2(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_121),
.B1(n_58),
.B2(n_60),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_100),
.B1(n_91),
.B2(n_106),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_79),
.B1(n_81),
.B2(n_64),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_97),
.B(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_82),
.B(n_35),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_105),
.B(n_102),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_35),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_100),
.B1(n_93),
.B2(n_106),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_152),
.B1(n_115),
.B2(n_124),
.Y(n_165)
);

OAI21x1_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_98),
.B(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_130),
.B(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_139),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_140),
.C(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_60),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_107),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_154),
.B(n_127),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_93),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_108),
.CI(n_101),
.CON(n_146),
.SN(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_150),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_35),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_151),
.C(n_113),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_67),
.B1(n_89),
.B2(n_81),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_89),
.C(n_58),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_33),
.B1(n_44),
.B2(n_24),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_24),
.B(n_33),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_123),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_27),
.Y(n_199)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_162),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_111),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_169),
.C(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_174),
.B1(n_132),
.B2(n_131),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_173),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_132),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_112),
.B(n_120),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_112),
.B(n_25),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_33),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_89),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_198),
.B1(n_169),
.B2(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_72),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_194),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_132),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_164),
.B1(n_157),
.B2(n_168),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_138),
.C(n_148),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_160),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_146),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_154),
.B1(n_72),
.B2(n_85),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_161),
.C(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_207),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_157),
.B1(n_156),
.B2(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_209),
.B1(n_218),
.B2(n_215),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_72),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_210),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_213),
.C(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_171),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_163),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_165),
.B1(n_183),
.B2(n_180),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_163),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_178),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_195),
.B(n_200),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_12),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_196),
.B1(n_198),
.B2(n_184),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_226),
.B1(n_12),
.B2(n_11),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_225),
.B1(n_232),
.B2(n_11),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_190),
.B1(n_199),
.B2(n_19),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_9),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_85),
.C(n_18),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_231),
.C(n_235),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_85),
.C(n_18),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_18),
.C(n_16),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_16),
.C(n_14),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_0),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_1),
.C(n_5),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_233),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_11),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_245),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_246),
.B(n_247),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_10),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_16),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_250),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_231),
.A2(n_10),
.B1(n_9),
.B2(n_4),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_236),
.B1(n_2),
.B2(n_4),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_10),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_221),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_259),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_221),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_255),
.B(n_239),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_14),
.B1(n_2),
.B2(n_5),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_14),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_249),
.C(n_7),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_268),
.C(n_270),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_240),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_267),
.C(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_260),
.B(n_6),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_6),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_272),
.B(n_261),
.C(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_251),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_277),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_275),
.B1(n_279),
.B2(n_265),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_6),
.B(n_7),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_8),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_275),
.A2(n_8),
.B(n_27),
.Y(n_282)
);

NAND2x1_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_278),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_280),
.B(n_283),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_27),
.Y(n_289)
);


endmodule