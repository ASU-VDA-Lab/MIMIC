module fake_jpeg_3432_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_54),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_43),
.B1(n_41),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_56),
.B1(n_49),
.B2(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_43),
.B1(n_41),
.B2(n_34),
.Y(n_56)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_71),
.B1(n_33),
.B2(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_13),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_35),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_58),
.B1(n_46),
.B2(n_3),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_16),
.C(n_30),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.C(n_65),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_14),
.C(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_89),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_62),
.B1(n_5),
.B2(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_92),
.Y(n_98)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.C(n_7),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_85),
.A3(n_17),
.B1(n_19),
.B2(n_31),
.C1(n_11),
.C2(n_12),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_103),
.B(n_8),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_22),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_8),
.B(n_9),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_111),
.B1(n_98),
.B2(n_104),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_110),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_86),
.C(n_91),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_106),
.CI(n_101),
.CON(n_113),
.SN(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_112),
.C(n_113),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_10),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_10),
.Y(n_120)
);


endmodule