module fake_jpeg_31405_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_17),
.B1(n_36),
.B2(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_3),
.Y(n_65)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_52),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_54),
.Y(n_74)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_4),
.Y(n_66)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_64),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_5),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_48),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_6),
.B(n_7),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_43),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_88),
.Y(n_95)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_89),
.Y(n_104)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_92),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_62),
.B1(n_50),
.B2(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_19),
.B1(n_33),
.B2(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_8),
.B(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_18),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_16),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_21),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_6),
.B(n_7),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

XNOR2x2_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_10),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_88),
.B(n_85),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_11),
.C(n_13),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.C(n_20),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_14),
.B(n_15),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_111),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.C(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_39),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_119),
.C(n_116),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_95),
.B1(n_99),
.B2(n_110),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.C(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_97),
.C(n_96),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_108),
.B1(n_117),
.B2(n_109),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);


endmodule