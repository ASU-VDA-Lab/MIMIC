module fake_jpeg_27841_n_76 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

BUFx12_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_14),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_33),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_16),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_16),
.B(n_13),
.C(n_14),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_23),
.B1(n_19),
.B2(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_47),
.B1(n_12),
.B2(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_23),
.B1(n_12),
.B2(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

A2O1A1O1Ixp25_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_29),
.B(n_9),
.C(n_8),
.D(n_21),
.Y(n_50)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_55),
.B(n_42),
.C(n_44),
.D(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_12),
.B1(n_8),
.B2(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_5),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_22),
.C(n_18),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_40),
.C(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_53),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_48),
.C(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_56),
.B1(n_57),
.B2(n_50),
.Y(n_65)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_61),
.C(n_62),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_1),
.A3(n_2),
.B1(n_6),
.B2(n_65),
.C1(n_66),
.C2(n_68),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_67),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_68),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_6),
.Y(n_76)
);


endmodule