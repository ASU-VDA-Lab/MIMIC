module real_jpeg_13084_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx10_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_26),
.B1(n_28),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_20),
.B1(n_24),
.B2(n_45),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_4),
.A2(n_26),
.B1(n_28),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_5),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_5),
.A2(n_30),
.B1(n_60),
.B2(n_72),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_5),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_7),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_7),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_9),
.B(n_23),
.C(n_26),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_20),
.B1(n_24),
.B2(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_41),
.B1(n_54),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_75),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_49),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_16),
.B(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_34),
.C(n_40),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_17)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_18),
.A2(n_29),
.B1(n_33),
.B2(n_85),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

OA22x2_ASAP7_75t_SL g37 ( 
.A1(n_20),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_20),
.A2(n_39),
.B(n_59),
.C(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_SL g23 ( 
.A(n_21),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_25)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_38),
.C(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_25),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_26),
.Y(n_28)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_33),
.B(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_59),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_37),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_39),
.B1(n_60),
.B2(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_46),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_41),
.A2(n_54),
.B1(n_88),
.B2(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_47),
.B(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_43),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_63),
.B1(n_64),
.B2(n_74),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_61),
.CON(n_59),
.SN(n_59)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_101),
.B(n_106),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_90),
.B(n_100),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_86),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_86),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_96),
.B(n_99),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_98),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);


endmodule