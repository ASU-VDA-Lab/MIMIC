module fake_netlist_6_4177_n_736 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_736);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_736;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_465;
wire n_367;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_449;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_643;
wire n_349;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_400;
wire n_284;
wire n_337;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_238;
wire n_573;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_447;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_535;
wire n_691;
wire n_250;
wire n_544;
wire n_372;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_611;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_624;
wire n_451;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_523;
wire n_322;
wire n_707;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_556;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_254;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_515;
wire n_434;
wire n_427;
wire n_288;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_484;
wire n_262;
wire n_613;
wire n_501;
wire n_531;
wire n_508;
wire n_663;
wire n_361;
wire n_379;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_112),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_15),
.Y(n_220)
);

INVxp33_ASAP7_75t_SL g221 ( 
.A(n_38),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_131),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_22),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_47),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_95),
.Y(n_229)
);

INVxp33_ASAP7_75t_SL g230 ( 
.A(n_158),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_101),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_11),
.B(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_109),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_30),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_16),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_50),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_20),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_53),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_113),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_136),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_8),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_23),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_86),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_69),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_159),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_90),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_150),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_42),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_98),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_198),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_108),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_57),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_92),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_51),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_4),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g275 ( 
.A(n_182),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_45),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_106),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_33),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_78),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_129),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_132),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_7),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_93),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_70),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_160),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_65),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_89),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_3),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_82),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_87),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_144),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_54),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_58),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_125),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_173),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_59),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_211),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_77),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_155),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_62),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_147),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_209),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_67),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_56),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_64),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_169),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_61),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_187),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_81),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_55),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_185),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_107),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_118),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_63),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_110),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_46),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_203),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_201),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_156),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_17),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_157),
.B(n_76),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_148),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_91),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_60),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_96),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_124),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_145),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_25),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_137),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_84),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_10),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_43),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_212),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_68),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_121),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_48),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_21),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_162),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_13),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_170),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_120),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_72),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_152),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_139),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_0),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_143),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_83),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_213),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_39),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_151),
.B(n_104),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_119),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_142),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_206),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_9),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_28),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_167),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_66),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_122),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_36),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_171),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_115),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_44),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_73),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_197),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_37),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_0),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_192),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_228),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_245),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_269),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_272),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_1),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_291),
.B(n_2),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_375),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_285),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_294),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_226),
.B(n_290),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_354),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_3),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_216),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_217),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_248),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_226),
.B(n_5),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_218),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_368),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_224),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_225),
.A2(n_5),
.B(n_6),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_219),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_220),
.B(n_6),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_227),
.Y(n_399)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_223),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_244),
.B(n_7),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_229),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_233),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_236),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_241),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_243),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_246),
.B(n_12),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_247),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_250),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_222),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_251),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_252),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_234),
.B(n_19),
.Y(n_413)
);

NAND2x1p5_ASAP7_75t_L g414 ( 
.A(n_329),
.B(n_24),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_254),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_26),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_255),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_256),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_257),
.A2(n_29),
.B(n_31),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_258),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_278),
.B(n_34),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_259),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_260),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_261),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_356),
.A2(n_337),
.B1(n_289),
.B2(n_327),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_264),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_265),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_267),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_268),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_270),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_287),
.B(n_317),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_355),
.A2(n_274),
.B(n_271),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_276),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_279),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_280),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_281),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_309),
.B(n_35),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_283),
.A2(n_40),
.B(n_41),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_286),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_273),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_292),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_293),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_340),
.B(n_49),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_295),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_296),
.Y(n_445)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_235),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_297),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_299),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_300),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_301),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_303),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_304),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_238),
.B(n_71),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_308),
.A2(n_74),
.B(n_75),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_311),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_312),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_315),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_316),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_319),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_242),
.B(n_79),
.Y(n_460)
);

AND2x4_ASAP7_75t_SL g461 ( 
.A(n_232),
.B(n_80),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_321),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_394),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_322),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_325),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_328),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_417),
.B(n_331),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_386),
.A2(n_266),
.B(n_249),
.C(n_344),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_459),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_323),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_359),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_421),
.B(n_332),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_221),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_380),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_431),
.B(n_238),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_460),
.B(n_302),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_382),
.B(n_400),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_410),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_425),
.B(n_230),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_398),
.B(n_333),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_407),
.B(n_231),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_413),
.B(n_334),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_400),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_377),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_416),
.B(n_358),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_408),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_381),
.B(n_376),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_446),
.A2(n_437),
.B1(n_388),
.B2(n_443),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_381),
.B(n_401),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_401),
.B(n_277),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_392),
.B(n_336),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_453),
.B(n_237),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_422),
.B(n_310),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_435),
.B(n_275),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_378),
.Y(n_511)
);

NAND2x1p5_ASAP7_75t_L g512 ( 
.A(n_432),
.B(n_341),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_429),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_414),
.B(n_439),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_379),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_389),
.B(n_343),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_439),
.B(n_318),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_442),
.B(n_338),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_436),
.B(n_390),
.Y(n_519)
);

BUFx4f_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_403),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_484),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_409),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_512),
.A2(n_454),
.B(n_438),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_474),
.A2(n_396),
.B1(n_447),
.B2(n_411),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_474),
.B(n_420),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_478),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_470),
.B(n_472),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_470),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_473),
.B(n_461),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_384),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_480),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_522),
.Y(n_537)
);

AND3x1_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_384),
.C(n_385),
.Y(n_538)
);

BUFx4f_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_469),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_475),
.B(n_412),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_491),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_483),
.B(n_347),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_506),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_482),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_502),
.B(n_424),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_484),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_489),
.A2(n_335),
.B1(n_350),
.B2(n_240),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_499),
.B(n_418),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_482),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_496),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_500),
.B(n_262),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_477),
.B(n_428),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_495),
.B(n_385),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_493),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_476),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_506),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_467),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_492),
.A2(n_486),
.B1(n_505),
.B2(n_494),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_479),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_477),
.B(n_441),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_503),
.A2(n_396),
.B1(n_448),
.B2(n_445),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_463),
.B(n_239),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_533),
.B(n_477),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_535),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_561),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_555),
.B(n_464),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_542),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_571),
.B(n_490),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_561),
.Y(n_579)
);

BUFx4_ASAP7_75t_SL g580 ( 
.A(n_548),
.Y(n_580)
);

BUFx2_ASAP7_75t_SL g581 ( 
.A(n_531),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_570),
.A2(n_419),
.B1(n_514),
.B2(n_326),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_538),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_535),
.B(n_521),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_565),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_556),
.Y(n_589)
);

BUFx4f_ASAP7_75t_SL g590 ( 
.A(n_553),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_571),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_568),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_527),
.A2(n_419),
.B1(n_330),
.B2(n_326),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_551),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_556),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_528),
.A2(n_239),
.B1(n_330),
.B2(n_360),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_567),
.A2(n_552),
.B1(n_539),
.B2(n_525),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_566),
.Y(n_598)
);

CKINVDCx6p67_ASAP7_75t_R g599 ( 
.A(n_541),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_559),
.B(n_569),
.C(n_560),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_545),
.A2(n_360),
.B1(n_240),
.B2(n_516),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_536),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_566),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_543),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_550),
.A2(n_465),
.B(n_466),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_SL g608 ( 
.A(n_530),
.B(n_346),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_534),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_589),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_583),
.A2(n_529),
.B1(n_572),
.B2(n_540),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_582),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_602),
.Y(n_616)
);

NAND2x1_ASAP7_75t_L g617 ( 
.A(n_612),
.B(n_544),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_584),
.A2(n_530),
.B1(n_540),
.B2(n_546),
.Y(n_618)
);

AOI222xp33_ASAP7_75t_L g619 ( 
.A1(n_597),
.A2(n_449),
.B1(n_452),
.B2(n_450),
.C1(n_444),
.C2(n_434),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_582),
.Y(n_620)
);

OAI222xp33_ASAP7_75t_L g621 ( 
.A1(n_596),
.A2(n_601),
.B1(n_593),
.B2(n_611),
.C1(n_578),
.C2(n_577),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_577),
.B(n_562),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_576),
.B(n_517),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_591),
.A2(n_540),
.B1(n_530),
.B2(n_298),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_SL g626 ( 
.A1(n_573),
.A2(n_600),
.B(n_298),
.C(n_263),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_600),
.A2(n_372),
.B1(n_374),
.B2(n_351),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_599),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_587),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_585),
.B(n_563),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_596),
.A2(n_434),
.B1(n_433),
.B2(n_458),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_607),
.B(n_508),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_574),
.B(n_564),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_601),
.A2(n_339),
.B1(n_263),
.B2(n_253),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_591),
.A2(n_433),
.B1(n_430),
.B2(n_458),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_592),
.A2(n_430),
.B1(n_253),
.B2(n_339),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

NAND2x1_ASAP7_75t_L g638 ( 
.A(n_612),
.B(n_554),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_610),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_634),
.A2(n_574),
.B1(n_603),
.B2(n_595),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_634),
.A2(n_579),
.B1(n_575),
.B2(n_598),
.C(n_594),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_632),
.A2(n_590),
.B1(n_586),
.B2(n_588),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_616),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_622),
.A2(n_603),
.B1(n_357),
.B2(n_366),
.Y(n_644)
);

OAI211xp5_ASAP7_75t_SL g645 ( 
.A1(n_619),
.A2(n_605),
.B(n_518),
.C(n_468),
.Y(n_645)
);

AO21x2_ASAP7_75t_L g646 ( 
.A1(n_626),
.A2(n_526),
.B(n_625),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_624),
.A2(n_581),
.B1(n_604),
.B2(n_282),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_629),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_SL g649 ( 
.A1(n_623),
.A2(n_370),
.B1(n_373),
.B2(n_353),
.Y(n_649)
);

OAI211xp5_ASAP7_75t_SL g650 ( 
.A1(n_636),
.A2(n_504),
.B(n_481),
.C(n_485),
.Y(n_650)
);

OAI211xp5_ASAP7_75t_L g651 ( 
.A1(n_613),
.A2(n_383),
.B(n_362),
.C(n_364),
.Y(n_651)
);

NAND2x1_ASAP7_75t_L g652 ( 
.A(n_633),
.B(n_586),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_617),
.A2(n_371),
.B(n_367),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_633),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_638),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_630),
.B(n_586),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_637),
.B(n_588),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_628),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_627),
.A2(n_369),
.B1(n_345),
.B2(n_588),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_639),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_615),
.B(n_554),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_620),
.Y(n_662)
);

AO21x2_ASAP7_75t_L g663 ( 
.A1(n_646),
.A2(n_621),
.B(n_614),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_656),
.B(n_618),
.Y(n_664)
);

NOR4xp25_ASAP7_75t_L g665 ( 
.A(n_645),
.B(n_621),
.C(n_650),
.D(n_651),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_660),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_643),
.Y(n_667)
);

AOI33xp33_ASAP7_75t_L g668 ( 
.A1(n_641),
.A2(n_636),
.A3(n_631),
.B1(n_640),
.B2(n_635),
.B3(n_383),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_654),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_656),
.B(n_631),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_648),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_647),
.A2(n_547),
.B1(n_554),
.B2(n_306),
.Y(n_672)
);

AOI221xp5_ASAP7_75t_L g673 ( 
.A1(n_649),
.A2(n_635),
.B1(n_423),
.B2(n_498),
.C(n_488),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_662),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_657),
.B(n_509),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_658),
.B(n_513),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_659),
.A2(n_510),
.B1(n_455),
.B2(n_456),
.C(n_451),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_661),
.B(n_580),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_644),
.A2(n_342),
.B1(n_288),
.B2(n_305),
.Y(n_679)
);

AOI221xp5_ASAP7_75t_L g680 ( 
.A1(n_642),
.A2(n_451),
.B1(n_457),
.B2(n_456),
.C(n_455),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_663),
.A2(n_653),
.B(n_608),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_670),
.B(n_661),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_667),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_664),
.B(n_652),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_671),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_674),
.Y(n_686)
);

NOR3xp33_ASAP7_75t_L g687 ( 
.A(n_672),
.B(n_652),
.C(n_532),
.Y(n_687)
);

AOI221xp5_ASAP7_75t_L g688 ( 
.A1(n_665),
.A2(n_457),
.B1(n_324),
.B2(n_361),
.C(n_352),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_664),
.A2(n_655),
.B1(n_349),
.B2(n_320),
.Y(n_689)
);

OAI33xp33_ASAP7_75t_L g690 ( 
.A1(n_675),
.A2(n_314),
.A3(n_313),
.B1(n_307),
.B2(n_284),
.B3(n_102),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_676),
.B(n_655),
.Y(n_691)
);

OAI211xp5_ASAP7_75t_L g692 ( 
.A1(n_665),
.A2(n_655),
.B(n_94),
.C(n_99),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_685),
.B(n_668),
.Y(n_693)
);

NAND5xp2_ASAP7_75t_L g694 ( 
.A(n_688),
.B(n_680),
.C(n_677),
.D(n_673),
.E(n_679),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_682),
.B(n_666),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_683),
.B(n_675),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_691),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_684),
.B(n_678),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_686),
.B(n_669),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_681),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_692),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_688),
.B(n_677),
.C(n_669),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_692),
.B(n_663),
.Y(n_703)
);

AND4x1_ASAP7_75t_L g704 ( 
.A(n_689),
.B(n_85),
.C(n_100),
.D(n_103),
.Y(n_704)
);

AOI21xp33_ASAP7_75t_SL g705 ( 
.A1(n_698),
.A2(n_687),
.B(n_681),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_697),
.B(n_105),
.Y(n_706)
);

AOI211xp5_ASAP7_75t_L g707 ( 
.A1(n_694),
.A2(n_690),
.B(n_114),
.C(n_116),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_697),
.B(n_215),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_696),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_703),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_695),
.B(n_111),
.Y(n_711)
);

XNOR2x1_ASAP7_75t_L g712 ( 
.A(n_706),
.B(n_698),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_709),
.B(n_701),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_709),
.B(n_700),
.Y(n_714)
);

OAI211xp5_ASAP7_75t_L g715 ( 
.A1(n_707),
.A2(n_702),
.B(n_693),
.C(n_699),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_710),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_714),
.B(n_705),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_712),
.Y(n_718)
);

AO22x1_ASAP7_75t_L g719 ( 
.A1(n_713),
.A2(n_711),
.B1(n_708),
.B2(n_704),
.Y(n_719)
);

OA22x2_ASAP7_75t_L g720 ( 
.A1(n_715),
.A2(n_713),
.B1(n_716),
.B2(n_130),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_123),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_719),
.B(n_214),
.C(n_133),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_717),
.A2(n_127),
.B(n_134),
.C(n_138),
.Y(n_723)
);

OAI211xp5_ASAP7_75t_SL g724 ( 
.A1(n_722),
.A2(n_720),
.B(n_141),
.C(n_149),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

AOI221xp5_ASAP7_75t_L g726 ( 
.A1(n_721),
.A2(n_140),
.B1(n_153),
.B2(n_163),
.C(n_164),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_SL g727 ( 
.A(n_722),
.B(n_165),
.C(n_168),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_725),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_728),
.Y(n_729)
);

AND3x4_ASAP7_75t_L g730 ( 
.A(n_729),
.B(n_724),
.C(n_727),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_730),
.B(n_174),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_730),
.B(n_726),
.C(n_179),
.Y(n_732)
);

AOI222xp33_ASAP7_75t_L g733 ( 
.A1(n_731),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.C1(n_184),
.C2(n_190),
.Y(n_733)
);

OA22x2_ASAP7_75t_L g734 ( 
.A1(n_732),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_734)
);

XNOR2xp5_ASAP7_75t_L g735 ( 
.A(n_734),
.B(n_200),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_735),
.A2(n_733),
.B(n_204),
.Y(n_736)
);


endmodule