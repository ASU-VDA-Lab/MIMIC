module fake_netlist_5_844_n_1939 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1939);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1939;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1817;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_7),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_143),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_34),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

INVxp33_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_48),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_145),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_90),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_24),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_150),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_179),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_57),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_137),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_84),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_112),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_110),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_2),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_72),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_89),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_182),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_0),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_25),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_68),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_134),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_105),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_96),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_77),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_34),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_133),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_91),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_7),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_27),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_57),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_20),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_35),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_126),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_36),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_161),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_62),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_194),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_55),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_99),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_111),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_177),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_29),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_38),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_70),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_189),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_38),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_11),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_46),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_51),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_26),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_140),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_18),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_86),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_71),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

BUFx2_ASAP7_75t_SL g295 ( 
.A(n_83),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_119),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_14),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_37),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_118),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_12),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_73),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_37),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_61),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_65),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_155),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_26),
.Y(n_308)
);

BUFx2_ASAP7_75t_SL g309 ( 
.A(n_107),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_92),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_65),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_163),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_185),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_4),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_184),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_48),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_42),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_3),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_116),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_178),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_78),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_15),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_11),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_29),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_55),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_171),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_9),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_149),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_128),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_159),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_80),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_81),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_42),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_151),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_113),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_132),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_30),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_176),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_122),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_191),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_75),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_47),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_68),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_168),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_50),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_82),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_43),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_20),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_123),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_98),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_32),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_35),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_53),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_31),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_172),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_15),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_193),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_54),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_61),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_6),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_40),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_49),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_67),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_9),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_124),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_66),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_21),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_24),
.Y(n_370)
);

BUFx8_ASAP7_75t_SL g371 ( 
.A(n_54),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_1),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_64),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_139),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_5),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_173),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_39),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_97),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_152),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_79),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_195),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_66),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_16),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_16),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_87),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_93),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_85),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_59),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_1),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_45),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_136),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_36),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_160),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_18),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_371),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_301),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_318),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_199),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_218),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_218),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_239),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_237),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_251),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_254),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_245),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_205),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_218),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_248),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_249),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_250),
.Y(n_410)
);

BUFx6f_ASAP7_75t_SL g411 ( 
.A(n_208),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_240),
.B(n_6),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_233),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_252),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_218),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_253),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_218),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_205),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_262),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_316),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_315),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_315),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_312),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_316),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_275),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_323),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_264),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_310),
.B(n_8),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_267),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_274),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_271),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_197),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_386),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_234),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_310),
.B(n_8),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_271),
.B(n_10),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_276),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_281),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_292),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_293),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

INVx4_ASAP7_75t_R g448 ( 
.A(n_374),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_301),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_300),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_198),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_307),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_320),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_328),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_242),
.B(n_10),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_330),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_331),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_332),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_333),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_385),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_208),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_334),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_374),
.B(n_226),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_226),
.B(n_12),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_366),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_366),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_336),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_301),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_337),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_212),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_301),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_212),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_338),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_208),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_341),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_346),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_348),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_375),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_351),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_200),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_214),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_244),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_200),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_247),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_260),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_214),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_261),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_202),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_236),
.B(n_13),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_263),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_301),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_406),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_396),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_497),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_375),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_466),
.B(n_375),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_449),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_449),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_421),
.B(n_202),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_431),
.B(n_204),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_400),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_471),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_487),
.B(n_225),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_455),
.B(n_442),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_475),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_415),
.B(n_204),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_475),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_397),
.B(n_259),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_225),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_437),
.B(n_236),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_420),
.B(n_206),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_397),
.B(n_259),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_424),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_474),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_437),
.B(n_246),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_422),
.B(n_242),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_422),
.B(n_354),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_426),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_429),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_429),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_432),
.B(n_206),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_207),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_246),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_447),
.Y(n_558)
);

NAND2x1_ASAP7_75t_L g559 ( 
.A(n_448),
.B(n_321),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_458),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_493),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_486),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_496),
.B(n_270),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_451),
.B(n_303),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_468),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_402),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_442),
.B(n_354),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_398),
.B(n_256),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_469),
.B(n_207),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_469),
.B(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_551),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_507),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_551),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_568),
.B(n_405),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_500),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_520),
.A2(n_455),
.B1(n_495),
.B2(n_467),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_524),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_512),
.B(n_408),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_540),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_551),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_520),
.A2(n_467),
.B1(n_412),
.B2(n_403),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_512),
.B(n_409),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_500),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_574),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_574),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_520),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_451),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_501),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_511),
.B(n_410),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_511),
.B(n_303),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_552),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_545),
.B(n_451),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_520),
.B(n_559),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_498),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_504),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_414),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_575),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_520),
.B(n_416),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_502),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_498),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_520),
.B(n_419),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_513),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_546),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_514),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_L g620 ( 
.A(n_559),
.B(n_395),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_514),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_532),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_520),
.B(n_430),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_518),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_502),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_518),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_546),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_523),
.Y(n_630)
);

AND3x2_ASAP7_75t_L g631 ( 
.A(n_563),
.B(n_403),
.C(n_297),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_519),
.A2(n_445),
.B1(n_446),
.B2(n_443),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_552),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_523),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_569),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_502),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_528),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_502),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_528),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_321),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_569),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_569),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_527),
.A2(n_440),
.B1(n_460),
.B2(n_450),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_530),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_533),
.B(n_543),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_533),
.B(n_321),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_531),
.Y(n_650)
);

AND3x2_ASAP7_75t_L g651 ( 
.A(n_563),
.B(n_413),
.C(n_476),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_531),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_533),
.B(n_321),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_433),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_575),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_520),
.A2(n_441),
.B1(n_462),
.B2(n_427),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_536),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_536),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_538),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_564),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_538),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_540),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_542),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_542),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_547),
.Y(n_666)
);

BUFx4f_ASAP7_75t_L g667 ( 
.A(n_543),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_508),
.B(n_435),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_506),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_452),
.C(n_444),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_547),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_541),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_543),
.B(n_321),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_541),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_543),
.B(n_201),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_537),
.B(n_453),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_548),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_548),
.Y(n_678)
);

XOR2x2_ASAP7_75t_L g679 ( 
.A(n_567),
.B(n_213),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_564),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_556),
.B(n_463),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_567),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_525),
.B(n_454),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_549),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_525),
.B(n_457),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_556),
.B(n_463),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_508),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_556),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_534),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_556),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_534),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_550),
.B(n_476),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_549),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_553),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_553),
.Y(n_695)
);

AND3x2_ASAP7_75t_L g696 ( 
.A(n_570),
.B(n_492),
.C(n_436),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_570),
.B(n_550),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_570),
.B(n_478),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_555),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_570),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_506),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_554),
.A2(n_441),
.B1(n_492),
.B2(n_576),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_554),
.B(n_478),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_561),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_459),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_577),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_506),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_561),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_562),
.B(n_203),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_562),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_565),
.B(n_461),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_565),
.B(n_479),
.C(n_472),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_573),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_573),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_540),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_577),
.B(n_481),
.C(n_436),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_506),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_544),
.B(n_268),
.C(n_266),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_544),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_544),
.Y(n_722)
);

AND2x6_ASAP7_75t_L g723 ( 
.A(n_506),
.B(n_209),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_560),
.B(n_464),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_560),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_560),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_560),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_499),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_499),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_688),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_689),
.A2(n_477),
.B1(n_480),
.B2(n_470),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_687),
.B(n_484),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_687),
.B(n_485),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_607),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_578),
.B(n_581),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_689),
.B(n_488),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_688),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_607),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_597),
.B(n_494),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_595),
.B(n_401),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_692),
.B(n_299),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_586),
.A2(n_373),
.B1(n_372),
.B2(n_230),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_588),
.B(n_540),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_618),
.B(n_210),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_691),
.B(n_411),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_595),
.B(n_404),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_592),
.B(n_540),
.Y(n_747)
);

INVx8_ASAP7_75t_L g748 ( 
.A(n_675),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_670),
.B(n_215),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_657),
.A2(n_591),
.B1(n_667),
.B2(n_702),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_707),
.B(n_557),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_690),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_707),
.B(n_557),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_597),
.B(n_359),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_692),
.B(n_411),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_600),
.B(n_557),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_683),
.A2(n_425),
.B1(n_428),
.B2(n_438),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_690),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_652),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_597),
.B(n_217),
.Y(n_760)
);

INVx8_ASAP7_75t_L g761 ( 
.A(n_675),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_666),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_632),
.B(n_215),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_618),
.B(n_227),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_597),
.B(n_232),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_697),
.B(n_557),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_693),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_667),
.A2(n_290),
.B1(n_322),
.B2(n_313),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_629),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_697),
.B(n_557),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_613),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_685),
.B(n_706),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_629),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_597),
.B(n_238),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_579),
.B(n_241),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_596),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_693),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_596),
.B(n_613),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_580),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_583),
.B(n_557),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_668),
.B(n_557),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_619),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_619),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_700),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_700),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_694),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_604),
.B(n_558),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_604),
.B(n_558),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_694),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_622),
.B(n_233),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_672),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_621),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_699),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_703),
.B(n_411),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_699),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_SL g796 ( 
.A(n_609),
.B(n_257),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_604),
.B(n_558),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_667),
.B(n_258),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_605),
.B(n_269),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_598),
.B(n_558),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_598),
.B(n_558),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_584),
.B(n_558),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_593),
.B(n_558),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_646),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_579),
.B(n_272),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_646),
.A2(n_503),
.B(n_499),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_622),
.B(n_233),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_599),
.B(n_566),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_603),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_608),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_674),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_714),
.Y(n_813)
);

INVx8_ASAP7_75t_L g814 ( 
.A(n_675),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_674),
.B(n_355),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_587),
.B(n_279),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_615),
.B(n_566),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_616),
.B(n_566),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_682),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_680),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_703),
.A2(n_295),
.B1(n_309),
.B2(n_352),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_676),
.A2(n_224),
.B1(n_222),
.B2(n_231),
.Y(n_822)
);

NOR2x1p5_ASAP7_75t_L g823 ( 
.A(n_680),
.B(n_235),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_617),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_682),
.B(n_355),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_661),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_644),
.B(n_277),
.C(n_273),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_587),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_624),
.B(n_566),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_627),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_594),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_630),
.B(n_566),
.Y(n_832)
);

CKINVDCx16_ASAP7_75t_R g833 ( 
.A(n_661),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_714),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_634),
.B(n_566),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_610),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_611),
.B(n_296),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_614),
.A2(n_340),
.B1(n_391),
.B2(n_378),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_700),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_637),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_656),
.B(n_284),
.C(n_283),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_639),
.B(n_566),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_645),
.B(n_571),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_620),
.B(n_211),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_715),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_648),
.B(n_571),
.Y(n_846)
);

BUFx8_ASAP7_75t_L g847 ( 
.A(n_594),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_696),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_679),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_650),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_580),
.Y(n_851)
);

INVx3_ASAP7_75t_R g852 ( 
.A(n_679),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_658),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_659),
.B(n_571),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_717),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_623),
.B(n_342),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_712),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_660),
.B(n_571),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_662),
.B(n_571),
.Y(n_859)
);

AO22x2_ASAP7_75t_L g860 ( 
.A1(n_601),
.A2(n_219),
.B1(n_229),
.B2(n_382),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_713),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_664),
.B(n_571),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_L g863 ( 
.A(n_675),
.B(n_216),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_665),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_671),
.B(n_571),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_655),
.B(n_343),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_677),
.B(n_515),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_724),
.B(n_216),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_L g869 ( 
.A(n_719),
.B(n_220),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_681),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_727),
.B(n_721),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_681),
.B(n_411),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_686),
.A2(n_221),
.B1(n_357),
.B2(n_367),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_686),
.B(n_698),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_698),
.B(n_220),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_601),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_678),
.B(n_355),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_684),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_695),
.B(n_704),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_675),
.A2(n_221),
.B1(n_367),
.B2(n_357),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_705),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_715),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_709),
.A2(n_389),
.B1(n_235),
.B2(n_368),
.C(n_377),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_582),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_675),
.A2(n_376),
.B1(n_379),
.B2(n_380),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_711),
.B(n_515),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_727),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_720),
.B(n_515),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_721),
.B(n_222),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_582),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_722),
.B(n_223),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_725),
.B(n_515),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_726),
.B(n_612),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_628),
.B(n_522),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_628),
.B(n_522),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_590),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_612),
.B(n_223),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_590),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_612),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_778),
.B(n_651),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_784),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_784),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_772),
.B(n_733),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_766),
.A2(n_653),
.B(n_649),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_735),
.B(n_628),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_876),
.B(n_636),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_857),
.B(n_636),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_812),
.B(n_631),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_750),
.B(n_636),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_879),
.B(n_654),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_879),
.B(n_654),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_831),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_733),
.B(n_265),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_770),
.A2(n_589),
.B(n_585),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_756),
.A2(n_589),
.B(n_585),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_874),
.A2(n_710),
.B1(n_653),
.B2(n_673),
.Y(n_916)
);

BUFx4f_ASAP7_75t_L g917 ( 
.A(n_844),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_784),
.B(n_839),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_732),
.B(n_228),
.C(n_224),
.Y(n_919)
);

AOI21x1_ASAP7_75t_L g920 ( 
.A1(n_871),
.A2(n_673),
.B(n_649),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_743),
.A2(n_589),
.B(n_585),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_828),
.B(n_243),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_747),
.A2(n_663),
.B(n_647),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_866),
.A2(n_800),
.B(n_801),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_784),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_740),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_802),
.A2(n_663),
.B(n_647),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_360),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_741),
.B(n_360),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_808),
.B(n_362),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_742),
.A2(n_394),
.B1(n_306),
.B2(n_311),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_875),
.A2(n_654),
.B(n_669),
.C(n_718),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_759),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_820),
.B(n_796),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_776),
.B(n_669),
.Y(n_935)
);

NOR2x2_ASAP7_75t_L g936 ( 
.A(n_844),
.B(n_448),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_759),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_839),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_781),
.A2(n_663),
.B(n_647),
.Y(n_939)
);

BUFx12f_ASAP7_75t_L g940 ( 
.A(n_847),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_782),
.B(n_669),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_780),
.A2(n_625),
.B(n_612),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_887),
.Y(n_943)
);

BUFx12f_ASAP7_75t_L g944 ( 
.A(n_847),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_746),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_742),
.A2(n_860),
.B1(n_866),
.B2(n_805),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_783),
.B(n_701),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_732),
.B(n_319),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_800),
.A2(n_718),
.B(n_701),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_870),
.B(n_344),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_807),
.A2(n_718),
.B(n_701),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_792),
.B(n_710),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_839),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_787),
.A2(n_797),
.B(n_788),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_762),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_899),
.A2(n_625),
.B(n_612),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_831),
.B(n_350),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_798),
.B(n_710),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_751),
.A2(n_626),
.B(n_625),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_753),
.A2(n_626),
.B(n_625),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_875),
.A2(n_635),
.B(n_606),
.C(n_643),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_837),
.A2(n_856),
.B(n_871),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_826),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_762),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_754),
.A2(n_626),
.B(n_625),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_730),
.B(n_710),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_839),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_791),
.B(n_602),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_754),
.A2(n_638),
.B(n_626),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_881),
.B(n_626),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_837),
.A2(n_856),
.B(n_799),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_799),
.A2(n_641),
.B(n_638),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_737),
.B(n_710),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_855),
.B(n_356),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_872),
.A2(n_635),
.B(n_606),
.C(n_643),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_872),
.A2(n_794),
.B(n_821),
.C(n_755),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_752),
.B(n_710),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_828),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_893),
.A2(n_785),
.B(n_761),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_794),
.A2(n_755),
.B(n_745),
.C(n_758),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_810),
.B(n_602),
.Y(n_981)
);

OAI321xp33_ASAP7_75t_L g982 ( 
.A1(n_883),
.A2(n_255),
.A3(n_278),
.B1(n_353),
.B2(n_339),
.C(n_329),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_893),
.A2(n_642),
.B(n_633),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_785),
.A2(n_708),
.B(n_641),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_861),
.B(n_361),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_815),
.B(n_363),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_734),
.B(n_738),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_736),
.B(n_228),
.C(n_231),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_891),
.A2(n_642),
.B(n_633),
.C(n_729),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_811),
.B(n_728),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_748),
.A2(n_638),
.B(n_708),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_836),
.B(n_370),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_769),
.B(n_392),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_739),
.A2(n_387),
.B1(n_376),
.B2(n_379),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_891),
.A2(n_729),
.B(n_728),
.C(n_288),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_889),
.A2(n_304),
.B(n_298),
.C(n_384),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_L g997 ( 
.A1(n_822),
.A2(n_377),
.B(n_363),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_771),
.B(n_352),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_824),
.B(n_638),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_748),
.A2(n_638),
.B(n_708),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_830),
.B(n_840),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_739),
.A2(n_640),
.B1(n_723),
.B2(n_381),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_748),
.A2(n_814),
.B(n_761),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_761),
.A2(n_708),
.B(n_641),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_850),
.B(n_641),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_853),
.B(n_641),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_814),
.A2(n_708),
.B(n_716),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_773),
.A2(n_387),
.B1(n_381),
.B2(n_393),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_L g1009 ( 
.A(n_731),
.B(n_380),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_767),
.A2(n_640),
.B(n_723),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_868),
.A2(n_640),
.B1(n_723),
.B2(n_393),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_864),
.B(n_640),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_744),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_825),
.Y(n_1014)
);

AND2x6_ASAP7_75t_L g1015 ( 
.A(n_877),
.B(n_744),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_878),
.B(n_640),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_814),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_736),
.B(n_364),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_767),
.B(n_716),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_764),
.B(n_640),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_819),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_764),
.B(n_280),
.Y(n_1022)
);

AND2x2_ASAP7_75t_SL g1023 ( 
.A(n_827),
.B(n_863),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_777),
.Y(n_1024)
);

OR2x6_ASAP7_75t_SL g1025 ( 
.A(n_852),
.B(n_364),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_786),
.B(n_522),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_868),
.A2(n_745),
.B(n_838),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_844),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_894),
.A2(n_716),
.B(n_522),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_789),
.B(n_723),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_789),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_819),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_793),
.A2(n_723),
.B(n_539),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_795),
.B(n_259),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_873),
.B(n_285),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_841),
.A2(n_369),
.B(n_368),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_895),
.A2(n_506),
.B(n_510),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_775),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_803),
.A2(n_510),
.B(n_517),
.Y(n_1039)
);

BUFx8_ASAP7_75t_L g1040 ( 
.A(n_848),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_795),
.B(n_510),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_804),
.A2(n_817),
.B(n_809),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_889),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_813),
.B(n_723),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_775),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_834),
.B(n_510),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_749),
.A2(n_473),
.B1(n_482),
.B2(n_490),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_760),
.A2(n_539),
.B(n_503),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_834),
.B(n_539),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_845),
.B(n_510),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_757),
.B(n_286),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_818),
.A2(n_535),
.B(n_510),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_845),
.B(n_503),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_806),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_829),
.A2(n_835),
.B(n_846),
.Y(n_1055)
);

OAI321xp33_ASAP7_75t_L g1056 ( 
.A1(n_768),
.A2(n_388),
.A3(n_305),
.B1(n_326),
.B2(n_282),
.C(n_482),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_869),
.B(n_287),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_833),
.Y(n_1058)
);

AOI22x1_ASAP7_75t_L g1059 ( 
.A1(n_882),
.A2(n_365),
.B1(n_369),
.B2(n_383),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_806),
.Y(n_1060)
);

OAI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_860),
.A2(n_365),
.B(n_383),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_860),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_882),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_816),
.A2(n_347),
.B(n_291),
.C(n_294),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_832),
.A2(n_535),
.B(n_510),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_842),
.A2(n_535),
.B(n_517),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_816),
.A2(n_490),
.B1(n_535),
.B2(n_521),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_843),
.A2(n_535),
.B(n_521),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_854),
.A2(n_535),
.B(n_521),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_849),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_884),
.B(n_505),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_763),
.B(n_823),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_884),
.B(n_505),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_858),
.A2(n_535),
.B(n_521),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_890),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_897),
.A2(n_521),
.B1(n_517),
.B2(n_516),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_880),
.A2(n_345),
.B1(n_302),
.B2(n_308),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_897),
.B(n_389),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_890),
.B(n_390),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_896),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_885),
.B(n_289),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_896),
.B(n_505),
.Y(n_1082)
);

AND2x4_ASAP7_75t_SL g1083 ( 
.A(n_898),
.B(n_517),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_760),
.A2(n_526),
.B(n_516),
.C(n_509),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_903),
.B(n_898),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_963),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_903),
.A2(n_886),
.B(n_867),
.C(n_862),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_925),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1018),
.B(n_314),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_954),
.A2(n_774),
.B(n_765),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_946),
.A2(n_1062),
.B1(n_976),
.B2(n_1035),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1035),
.A2(n_865),
.B(n_859),
.C(n_851),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_928),
.B(n_317),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_925),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1075),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_915),
.A2(n_774),
.B(n_765),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_919),
.B(n_892),
.C(n_888),
.Y(n_1097)
);

AOI22x1_ASAP7_75t_L g1098 ( 
.A1(n_971),
.A2(n_779),
.B1(n_324),
.B2(n_349),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_948),
.A2(n_325),
.B1(n_327),
.B2(n_335),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_925),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_933),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_940),
.B(n_521),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_948),
.B(n_390),
.C(n_516),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1027),
.A2(n_526),
.B(n_509),
.C(n_19),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1043),
.B(n_526),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_937),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_992),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_913),
.A2(n_509),
.B(n_521),
.C(n_517),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_934),
.B(n_517),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_992),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_921),
.A2(n_923),
.B(n_939),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_914),
.A2(n_517),
.B(n_74),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_913),
.A2(n_13),
.B(n_17),
.C(n_19),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1043),
.B(n_17),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_925),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_938),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_930),
.B(n_21),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_905),
.A2(n_101),
.B(n_186),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_985),
.B(n_22),
.Y(n_1119)
);

CKINVDCx14_ASAP7_75t_R g1120 ( 
.A(n_1058),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_986),
.B(n_22),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_950),
.B(n_27),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_985),
.B(n_28),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_980),
.A2(n_31),
.B(n_33),
.C(n_40),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_938),
.B(n_109),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_912),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_951),
.A2(n_108),
.B(n_180),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1045),
.B(n_102),
.Y(n_1128)
);

OAI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_1051),
.A2(n_33),
.B(n_41),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1075),
.Y(n_1130)
);

INVxp67_ASAP7_75t_R g1131 ( 
.A(n_1072),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_942),
.A2(n_94),
.B(n_174),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_931),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_946),
.B(n_114),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_912),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_910),
.B(n_115),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1001),
.B(n_44),
.Y(n_1137)
);

OAI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_1051),
.A2(n_45),
.B(n_49),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1045),
.B(n_125),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1015),
.A2(n_121),
.B1(n_170),
.B2(n_166),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_938),
.B(n_192),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_938),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_974),
.B(n_50),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_988),
.A2(n_52),
.B(n_53),
.C(n_56),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_978),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_1061),
.B(n_52),
.C(n_56),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_916),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1147)
);

NOR2xp67_ASAP7_75t_L g1148 ( 
.A(n_1014),
.B(n_138),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_988),
.A2(n_58),
.B(n_60),
.C(n_62),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_974),
.B(n_950),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1038),
.B(n_156),
.Y(n_1151)
);

AO32x2_ASAP7_75t_L g1152 ( 
.A1(n_1080),
.A2(n_63),
.A3(n_64),
.B1(n_69),
.B2(n_165),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1015),
.A2(n_135),
.B1(n_142),
.B2(n_157),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_901),
.B(n_158),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_926),
.B(n_63),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_955),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_927),
.A2(n_162),
.B(n_69),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_957),
.B(n_993),
.C(n_900),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_932),
.A2(n_909),
.B(n_970),
.C(n_958),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_904),
.A2(n_909),
.B(n_1042),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_953),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_978),
.B(n_945),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_970),
.A2(n_952),
.B(n_973),
.C(n_966),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_978),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_964),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1055),
.A2(n_911),
.B(n_979),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1015),
.A2(n_919),
.B1(n_1013),
.B2(n_1060),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1078),
.A2(n_1015),
.B1(n_957),
.B2(n_1013),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_978),
.B(n_968),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_924),
.A2(n_961),
.B(n_975),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_993),
.B(n_1079),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_943),
.A2(n_1023),
.B1(n_1054),
.B2(n_990),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_953),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1015),
.A2(n_1023),
.B1(n_1054),
.B2(n_1081),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_929),
.B(n_922),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_944),
.B(n_1032),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1024),
.B(n_1031),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_922),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_962),
.A2(n_982),
.B(n_1064),
.C(n_997),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_901),
.B(n_902),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1022),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_917),
.B(n_1028),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1022),
.B(n_908),
.Y(n_1183)
);

O2A1O1Ixp5_ASAP7_75t_L g1184 ( 
.A1(n_918),
.A2(n_1019),
.B(n_1034),
.C(n_1057),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_902),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1034),
.A2(n_1077),
.B(n_994),
.C(n_996),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_984),
.A2(n_1007),
.B(n_1004),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_1040),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_987),
.B(n_998),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_967),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_991),
.A2(n_1000),
.B(n_977),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1036),
.A2(n_1056),
.B(n_995),
.C(n_1008),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1063),
.B(n_906),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1080),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_959),
.A2(n_960),
.B(n_956),
.Y(n_1195)
);

OAI21xp33_ASAP7_75t_SL g1196 ( 
.A1(n_981),
.A2(n_918),
.B(n_1012),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_967),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1017),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1017),
.B(n_1003),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_907),
.A2(n_999),
.B(n_1005),
.C(n_1006),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_935),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1021),
.B(n_1070),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1009),
.B(n_1020),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1040),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_989),
.A2(n_1016),
.B(n_1028),
.C(n_917),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1025),
.A2(n_936),
.B1(n_1002),
.B2(n_1011),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1049),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_941),
.B(n_947),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_949),
.A2(n_1047),
.B1(n_1030),
.B2(n_1044),
.C(n_983),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_SL g1210 ( 
.A(n_1067),
.B(n_1010),
.C(n_965),
.Y(n_1210)
);

BUFx4f_ASAP7_75t_L g1211 ( 
.A(n_1083),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1059),
.A2(n_920),
.B1(n_1053),
.B2(n_972),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1026),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1071),
.A2(n_1073),
.B1(n_1082),
.B2(n_1033),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1048),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_969),
.A2(n_1029),
.B(n_1050),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1041),
.B(n_1050),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1046),
.Y(n_1218)
);

O2A1O1Ixp5_ASAP7_75t_L g1219 ( 
.A1(n_1037),
.A2(n_1039),
.B(n_1052),
.C(n_1065),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1076),
.B(n_1066),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1068),
.B(n_1069),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1074),
.A2(n_597),
.B(n_667),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1084),
.A2(n_597),
.B(n_667),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_903),
.B(n_772),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_925),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_903),
.B(n_772),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_903),
.A2(n_772),
.B(n_1035),
.C(n_868),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_903),
.B(n_772),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_SL g1229 ( 
.A(n_925),
.B(n_784),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1058),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_912),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_954),
.A2(n_597),
.B(n_667),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_912),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1058),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1075),
.Y(n_1235)
);

AO21x1_ASAP7_75t_L g1236 ( 
.A1(n_903),
.A2(n_772),
.B(n_750),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_940),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_903),
.B(n_772),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1228),
.B(n_1238),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1160),
.A2(n_1166),
.B(n_1232),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1236),
.A2(n_1108),
.A3(n_1212),
.B(n_1091),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1212),
.A2(n_1091),
.A3(n_1172),
.B(n_1220),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1086),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1234),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_SL g1246 ( 
.A1(n_1179),
.A2(n_1134),
.B(n_1205),
.C(n_1227),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1238),
.A2(n_1224),
.B1(n_1226),
.B2(n_1150),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1136),
.A2(n_1221),
.B(n_1195),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1095),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1231),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1224),
.A2(n_1226),
.B(n_1170),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1172),
.A2(n_1216),
.A3(n_1092),
.B(n_1214),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1222),
.A2(n_1090),
.B(n_1159),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1231),
.B(n_1126),
.Y(n_1254)
);

AOI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1119),
.A2(n_1123),
.B1(n_1143),
.B2(n_1129),
.C(n_1138),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1219),
.A2(n_1127),
.B(n_1199),
.Y(n_1256)
);

AO32x2_ASAP7_75t_L g1257 ( 
.A1(n_1147),
.A2(n_1133),
.A3(n_1206),
.B1(n_1214),
.B2(n_1152),
.Y(n_1257)
);

OAI22x1_ASAP7_75t_L g1258 ( 
.A1(n_1167),
.A2(n_1122),
.B1(n_1174),
.B2(n_1189),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1229),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1171),
.B(n_1130),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1235),
.B(n_1085),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_SL g1262 ( 
.A1(n_1134),
.A2(n_1113),
.B(n_1128),
.C(n_1139),
.Y(n_1262)
);

OA22x2_ASAP7_75t_L g1263 ( 
.A1(n_1233),
.A2(n_1099),
.B1(n_1147),
.B2(n_1178),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1170),
.A2(n_1136),
.B(n_1163),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1196),
.A2(n_1104),
.B(n_1087),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_L g1266 ( 
.A(n_1173),
.B(n_1158),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1183),
.B(n_1182),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_SL g1268 ( 
.A1(n_1186),
.A2(n_1192),
.B(n_1114),
.C(n_1124),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1208),
.A2(n_1096),
.B(n_1223),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1157),
.A2(n_1210),
.B1(n_1103),
.B2(n_1112),
.C(n_1097),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1135),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1184),
.A2(n_1137),
.B(n_1200),
.C(n_1144),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1211),
.A2(n_1209),
.B(n_1193),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1211),
.A2(n_1193),
.B(n_1199),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1175),
.A2(n_1168),
.B1(n_1089),
.B2(n_1121),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1201),
.A2(n_1109),
.B(n_1207),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1149),
.A2(n_1097),
.B(n_1146),
.C(n_1203),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1117),
.B(n_1093),
.C(n_1098),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1194),
.A2(n_1203),
.B1(n_1165),
.B2(n_1156),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1217),
.A2(n_1177),
.B(n_1132),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1101),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1181),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1169),
.A2(n_1177),
.B(n_1213),
.Y(n_1283)
);

AOI21xp33_ASAP7_75t_L g1284 ( 
.A1(n_1162),
.A2(n_1110),
.B(n_1107),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1106),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1118),
.A2(n_1161),
.B(n_1105),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_L g1287 ( 
.A(n_1173),
.B(n_1164),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1198),
.A2(n_1215),
.B(n_1190),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1088),
.A2(n_1100),
.A3(n_1152),
.B(n_1215),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1151),
.A2(n_1131),
.B1(n_1155),
.B2(n_1148),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1151),
.B(n_1164),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1198),
.A2(n_1215),
.B(n_1190),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1237),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1088),
.A2(n_1100),
.B1(n_1145),
.B2(n_1164),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1125),
.B(n_1188),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1140),
.A2(n_1153),
.B1(n_1218),
.B2(n_1145),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1125),
.A2(n_1094),
.B(n_1115),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1120),
.A2(n_1102),
.B(n_1202),
.C(n_1176),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1145),
.B(n_1230),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1185),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1094),
.A2(n_1115),
.B(n_1116),
.Y(n_1301)
);

AO32x2_ASAP7_75t_L g1302 ( 
.A1(n_1152),
.A2(n_1218),
.A3(n_1125),
.B1(n_1141),
.B2(n_1154),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1218),
.B(n_1197),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1204),
.Y(n_1304)
);

CKINVDCx6p67_ASAP7_75t_R g1305 ( 
.A(n_1176),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1102),
.A2(n_1176),
.B(n_1142),
.C(n_1116),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1102),
.B(n_1185),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1197),
.B(n_1180),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1197),
.A2(n_772),
.B(n_1227),
.C(n_1150),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1225),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1125),
.A2(n_1236),
.A3(n_1108),
.B(n_1212),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1227),
.A2(n_772),
.B(n_1150),
.C(n_903),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1095),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1236),
.A2(n_1108),
.A3(n_1212),
.B(n_1091),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1183),
.B(n_1182),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1179),
.A2(n_976),
.B(n_1134),
.C(n_1205),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1236),
.A2(n_1108),
.A3(n_1212),
.B(n_1091),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1227),
.A2(n_772),
.B(n_1150),
.C(n_903),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1183),
.B(n_1182),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1095),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1198),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1086),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1086),
.Y(n_1326)
);

O2A1O1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1150),
.A2(n_772),
.B(n_1123),
.C(n_1119),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1095),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1227),
.A2(n_772),
.B(n_1160),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1236),
.A2(n_1108),
.A3(n_1212),
.B(n_1091),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1150),
.A2(n_772),
.B(n_1123),
.C(n_1119),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1150),
.A2(n_772),
.B1(n_1123),
.B2(n_1119),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1228),
.A2(n_772),
.B1(n_796),
.B2(n_934),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1150),
.A2(n_772),
.B(n_1027),
.C(n_976),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1150),
.A2(n_772),
.B(n_1123),
.C(n_1119),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1198),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1126),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1150),
.B(n_772),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1228),
.A2(n_772),
.B1(n_1226),
.B2(n_1224),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1086),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1086),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1228),
.B(n_1224),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1228),
.A2(n_772),
.B1(n_796),
.B2(n_934),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1225),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1227),
.A2(n_772),
.B(n_1160),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1150),
.A2(n_772),
.B(n_1123),
.C(n_1119),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1126),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1228),
.B(n_1224),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1095),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1234),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1236),
.A2(n_1108),
.A3(n_1212),
.B(n_1091),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1227),
.A2(n_772),
.B(n_1150),
.C(n_903),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1234),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_L g1364 ( 
.A(n_1097),
.B(n_857),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1228),
.B(n_1224),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1095),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1224),
.B(n_836),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1183),
.B(n_1182),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1236),
.A2(n_1108),
.A3(n_1212),
.B(n_1091),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1170),
.A2(n_1160),
.B(n_1166),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1126),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1150),
.A2(n_772),
.B1(n_1035),
.B2(n_948),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1160),
.A2(n_597),
.B(n_772),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1126),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1377)
);

NAND2xp33_ASAP7_75t_SL g1378 ( 
.A(n_1229),
.B(n_772),
.Y(n_1378)
);

NAND2xp33_ASAP7_75t_L g1379 ( 
.A(n_1228),
.B(n_772),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1150),
.B(n_772),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1225),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1150),
.B(n_934),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1150),
.B(n_772),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1228),
.B(n_1224),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1150),
.A2(n_772),
.B(n_1123),
.C(n_1119),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1198),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1191),
.A2(n_1187),
.B(n_1111),
.Y(n_1389)
);

AO21x1_ASAP7_75t_L g1390 ( 
.A1(n_1227),
.A2(n_772),
.B(n_1091),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1391)
);

BUFx8_ASAP7_75t_L g1392 ( 
.A(n_1341),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1263),
.A2(n_1295),
.B1(n_1247),
.B2(n_1343),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1295),
.A2(n_1302),
.B1(n_1379),
.B2(n_1251),
.Y(n_1394)
);

BUFx8_ASAP7_75t_SL g1395 ( 
.A(n_1245),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1244),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1249),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1334),
.A2(n_1255),
.B1(n_1387),
.B2(n_1327),
.Y(n_1398)
);

AOI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1333),
.A2(n_1351),
.B(n_1337),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1313),
.Y(n_1400)
);

AOI21xp33_ASAP7_75t_L g1401 ( 
.A1(n_1334),
.A2(n_1347),
.B(n_1335),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1325),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1390),
.A2(n_1382),
.B1(n_1251),
.B2(n_1258),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1239),
.B(n_1346),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1331),
.A2(n_1350),
.B1(n_1354),
.B2(n_1386),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1293),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1250),
.B(n_1323),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1369),
.A2(n_1365),
.B1(n_1290),
.B2(n_1320),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1250),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1326),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1348),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1322),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1356),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1275),
.A2(n_1265),
.B1(n_1321),
.B2(n_1370),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1312),
.B(n_1361),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1305),
.Y(n_1416)
);

CKINVDCx11_ASAP7_75t_R g1417 ( 
.A(n_1304),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1260),
.B(n_1261),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1267),
.B(n_1317),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1275),
.A2(n_1267),
.B1(n_1370),
.B2(n_1321),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1290),
.A2(n_1309),
.B1(n_1317),
.B2(n_1278),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1366),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1344),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1278),
.A2(n_1266),
.B1(n_1364),
.B2(n_1273),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1364),
.A2(n_1264),
.B1(n_1330),
.B2(n_1378),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1271),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1284),
.A2(n_1296),
.B1(n_1285),
.B2(n_1281),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1345),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1339),
.B(n_1388),
.Y(n_1429)
);

INVx8_ASAP7_75t_L g1430 ( 
.A(n_1348),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1310),
.Y(n_1431)
);

CKINVDCx9p33_ASAP7_75t_R g1432 ( 
.A(n_1303),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1353),
.Y(n_1433)
);

BUFx4f_ASAP7_75t_L g1434 ( 
.A(n_1381),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1299),
.A2(n_1262),
.B1(n_1362),
.B2(n_1357),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1282),
.A2(n_1279),
.B1(n_1376),
.B2(n_1373),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1308),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1291),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1381),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1289),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1372),
.A2(n_1283),
.B1(n_1276),
.B2(n_1257),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1277),
.A2(n_1268),
.B1(n_1246),
.B2(n_1318),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1372),
.A2(n_1257),
.B1(n_1274),
.B2(n_1280),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1381),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1259),
.A2(n_1300),
.B1(n_1297),
.B2(n_1307),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1307),
.A2(n_1272),
.B1(n_1297),
.B2(n_1287),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1289),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1336),
.A2(n_1242),
.B1(n_1289),
.B2(n_1253),
.Y(n_1448)
);

INVx2_ASAP7_75t_R g1449 ( 
.A(n_1311),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1294),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1301),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1288),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1286),
.A2(n_1269),
.B1(n_1375),
.B2(n_1368),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1306),
.Y(n_1454)
);

BUFx12f_ASAP7_75t_L g1455 ( 
.A(n_1298),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1242),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1242),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1292),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1314),
.A2(n_1338),
.B1(n_1367),
.B2(n_1360),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1270),
.A2(n_1329),
.B1(n_1328),
.B2(n_1324),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1248),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1311),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1352),
.A2(n_1359),
.B1(n_1355),
.B2(n_1240),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1241),
.B(n_1371),
.Y(n_1464)
);

CKINVDCx14_ASAP7_75t_R g1465 ( 
.A(n_1311),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1252),
.B(n_1371),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1316),
.A2(n_1358),
.B1(n_1371),
.B2(n_1319),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1243),
.A2(n_1389),
.B1(n_1315),
.B2(n_1385),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1256),
.B(n_1340),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1332),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1349),
.A2(n_1363),
.B1(n_1377),
.B2(n_1383),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1332),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1358),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1358),
.A2(n_1342),
.B1(n_1384),
.B2(n_1380),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1310),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1250),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1244),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1334),
.A2(n_772),
.B1(n_1384),
.B2(n_1380),
.Y(n_1478)
);

CKINVDCx6p67_ASAP7_75t_R g1479 ( 
.A(n_1293),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1271),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1249),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1249),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1341),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1334),
.A2(n_772),
.B1(n_1374),
.B2(n_1342),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1271),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1254),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1249),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1293),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1374),
.A2(n_796),
.B1(n_1150),
.B2(n_772),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1342),
.B(n_1380),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1249),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1249),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1342),
.A2(n_1133),
.B1(n_931),
.B2(n_1380),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1348),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1342),
.A2(n_1133),
.B1(n_931),
.B2(n_1380),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1293),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1244),
.Y(n_1500)
);

BUFx12f_ASAP7_75t_L g1501 ( 
.A(n_1293),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1342),
.B(n_1380),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1293),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1334),
.A2(n_772),
.B1(n_1374),
.B2(n_1342),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1245),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1250),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1348),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1249),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1380),
.B2(n_1374),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1244),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1323),
.Y(n_1513)
);

AO21x1_ASAP7_75t_L g1514 ( 
.A1(n_1398),
.A2(n_1399),
.B(n_1485),
.Y(n_1514)
);

BUFx2_ASAP7_75t_SL g1515 ( 
.A(n_1458),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1440),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1447),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1456),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1451),
.B(n_1420),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1496),
.A2(n_1498),
.B1(n_1504),
.B2(n_1490),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1457),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1407),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1391),
.B(n_1482),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1491),
.A2(n_1482),
.B(n_1391),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1461),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1455),
.A2(n_1408),
.B1(n_1421),
.B2(n_1502),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1469),
.A2(n_1463),
.B(n_1453),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1469),
.A2(n_1463),
.B(n_1453),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1473),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1490),
.B(n_1493),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1466),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1464),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1394),
.B(n_1465),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1472),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1409),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1467),
.B(n_1470),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1394),
.B(n_1465),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1448),
.Y(n_1538)
);

NAND2x1p5_ASAP7_75t_L g1539 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1403),
.B(n_1474),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1409),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1496),
.B(n_1498),
.C(n_1508),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1403),
.B(n_1474),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1448),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1476),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1397),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1487),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1400),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1462),
.B(n_1405),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1476),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1412),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1413),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1493),
.B(n_1507),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1405),
.B(n_1443),
.Y(n_1554)
);

NAND3xp33_ASAP7_75t_SL g1555 ( 
.A(n_1507),
.B(n_1511),
.C(n_1508),
.Y(n_1555)
);

CKINVDCx6p67_ASAP7_75t_R g1556 ( 
.A(n_1501),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1443),
.B(n_1414),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1422),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1481),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1483),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1488),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1414),
.B(n_1438),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1506),
.B(n_1441),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1506),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1494),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1495),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1392),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1510),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1511),
.A2(n_1492),
.B1(n_1478),
.B2(n_1435),
.Y(n_1569)
);

AND2x4_ASAP7_75t_SL g1570 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1449),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1449),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1415),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1442),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1441),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1425),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1450),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1429),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1460),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1460),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1452),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1459),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1419),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1459),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1424),
.Y(n_1585)
);

AO21x1_ASAP7_75t_SL g1586 ( 
.A1(n_1401),
.A2(n_1427),
.B(n_1436),
.Y(n_1586)
);

AO21x2_ASAP7_75t_L g1587 ( 
.A1(n_1478),
.A2(n_1404),
.B(n_1471),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1433),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1468),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1471),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1427),
.A2(n_1513),
.B(n_1436),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1393),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1432),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1418),
.B(n_1393),
.Y(n_1595)
);

BUFx8_ASAP7_75t_L g1596 ( 
.A(n_1480),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1445),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1437),
.B(n_1486),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1432),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1411),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1430),
.A2(n_1434),
.B(n_1509),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1426),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1439),
.B(n_1509),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1426),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_SL g1605 ( 
.A1(n_1444),
.A2(n_1410),
.B(n_1477),
.C(n_1499),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1395),
.Y(n_1606)
);

NAND2x1p5_ASAP7_75t_L g1607 ( 
.A(n_1581),
.B(n_1475),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1606),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1527),
.A2(n_1505),
.B(n_1509),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1542),
.A2(n_1434),
.B(n_1431),
.Y(n_1610)
);

AO32x2_ASAP7_75t_L g1611 ( 
.A1(n_1564),
.A2(n_1475),
.A3(n_1431),
.B1(n_1392),
.B2(n_1484),
.Y(n_1611)
);

NAND4xp25_ASAP7_75t_L g1612 ( 
.A(n_1520),
.B(n_1428),
.C(n_1396),
.D(n_1423),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1526),
.A2(n_1406),
.B1(n_1503),
.B2(n_1489),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1524),
.A2(n_1430),
.B(n_1497),
.C(n_1484),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1555),
.A2(n_1402),
.B(n_1500),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1545),
.B(n_1479),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1570),
.A2(n_1430),
.B(n_1497),
.C(n_1416),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1550),
.B(n_1497),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1550),
.B(n_1497),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1569),
.A2(n_1417),
.B1(n_1402),
.B2(n_1500),
.C(n_1512),
.Y(n_1620)
);

BUFx12f_ASAP7_75t_L g1621 ( 
.A(n_1567),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1518),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1535),
.B(n_1541),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1583),
.B(n_1549),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1583),
.B(n_1549),
.Y(n_1625)
);

AOI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1514),
.A2(n_1530),
.B(n_1523),
.C(n_1553),
.Y(n_1626)
);

AOI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1514),
.A2(n_1593),
.B1(n_1540),
.B2(n_1543),
.C(n_1579),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1539),
.A2(n_1584),
.B(n_1582),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1540),
.A2(n_1543),
.B1(n_1580),
.B2(n_1579),
.C(n_1585),
.Y(n_1629)
);

BUFx12f_ASAP7_75t_L g1630 ( 
.A(n_1567),
.Y(n_1630)
);

BUFx12f_ASAP7_75t_L g1631 ( 
.A(n_1567),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1597),
.A2(n_1595),
.B1(n_1562),
.B2(n_1585),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1521),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1521),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1563),
.B(n_1534),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1539),
.A2(n_1605),
.B(n_1595),
.C(n_1597),
.Y(n_1636)
);

BUFx8_ASAP7_75t_L g1637 ( 
.A(n_1525),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1580),
.A2(n_1515),
.B(n_1594),
.C(n_1592),
.Y(n_1638)
);

AOI22x1_ASAP7_75t_SL g1639 ( 
.A1(n_1599),
.A2(n_1574),
.B1(n_1547),
.B2(n_1544),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1515),
.A2(n_1594),
.B(n_1592),
.C(n_1576),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1563),
.B(n_1532),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1582),
.B(n_1584),
.C(n_1574),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1576),
.A2(n_1557),
.B(n_1554),
.C(n_1537),
.Y(n_1643)
);

AO32x2_ASAP7_75t_L g1644 ( 
.A1(n_1522),
.A2(n_1600),
.A3(n_1532),
.B1(n_1544),
.B2(n_1538),
.Y(n_1644)
);

AOI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1525),
.A2(n_1591),
.B(n_1590),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1538),
.A2(n_1554),
.B1(n_1557),
.B2(n_1539),
.C(n_1575),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1583),
.B(n_1599),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1519),
.A2(n_1598),
.B(n_1573),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1602),
.A2(n_1604),
.B1(n_1588),
.B2(n_1573),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1562),
.B(n_1533),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1519),
.B(n_1603),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1519),
.B(n_1551),
.Y(n_1652)
);

AO21x2_ASAP7_75t_L g1653 ( 
.A1(n_1527),
.A2(n_1528),
.B(n_1589),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1552),
.B(n_1558),
.Y(n_1654)
);

AND2x6_ASAP7_75t_L g1655 ( 
.A(n_1577),
.B(n_1578),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1559),
.B(n_1560),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1601),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_R g1658 ( 
.A(n_1556),
.B(n_1600),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1596),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1528),
.A2(n_1536),
.B(n_1586),
.C(n_1577),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1641),
.B(n_1536),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1653),
.B(n_1571),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1609),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1653),
.B(n_1644),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1656),
.B(n_1587),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1609),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1655),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1622),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1644),
.B(n_1571),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1644),
.B(n_1572),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1652),
.B(n_1572),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1635),
.B(n_1531),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1613),
.A2(n_1586),
.B1(n_1587),
.B2(n_1596),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1634),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1531),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1650),
.B(n_1529),
.Y(n_1677)
);

NOR2xp67_ASAP7_75t_L g1678 ( 
.A(n_1642),
.B(n_1566),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1655),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1613),
.A2(n_1587),
.B1(n_1546),
.B2(n_1548),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1654),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1639),
.A2(n_1568),
.B1(n_1565),
.B2(n_1561),
.Y(n_1682)
);

BUFx8_ASAP7_75t_L g1683 ( 
.A(n_1611),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1655),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1647),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1657),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1668),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1665),
.B(n_1618),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1680),
.B(n_1626),
.C(n_1627),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1669),
.B(n_1624),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1669),
.B(n_1619),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1661),
.B(n_1672),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1625),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1662),
.A2(n_1645),
.B(n_1640),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1673),
.A2(n_1620),
.B1(n_1646),
.B2(n_1629),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1674),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1670),
.B(n_1664),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1670),
.B(n_1664),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1680),
.A2(n_1643),
.B1(n_1636),
.B2(n_1632),
.C(n_1612),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1675),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1675),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1632),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_1685),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1675),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1657),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1681),
.B(n_1628),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1687),
.A2(n_1638),
.B1(n_1648),
.B2(n_1615),
.C(n_1610),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1671),
.B(n_1516),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1674),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1677),
.B(n_1517),
.Y(n_1712)
);

BUFx8_ASAP7_75t_SL g1713 ( 
.A(n_1686),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1679),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1621),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1695),
.B(n_1678),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1698),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1696),
.B(n_1684),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1704),
.B(n_1677),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1699),
.B(n_1663),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1699),
.B(n_1663),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1707),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1709),
.B(n_1682),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1699),
.B(n_1663),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1700),
.B(n_1663),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1700),
.B(n_1663),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1704),
.B(n_1677),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1708),
.B(n_1711),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1663),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1693),
.B(n_1676),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1708),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1696),
.B(n_1684),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1702),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1690),
.B(n_1630),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1689),
.B(n_1676),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1702),
.Y(n_1739)
);

NAND2x1p5_ASAP7_75t_L g1740 ( 
.A(n_1714),
.B(n_1679),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1697),
.A2(n_1682),
.B1(n_1673),
.B2(n_1678),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1688),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_1676),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1714),
.B(n_1667),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1663),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1714),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1705),
.B(n_1666),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1696),
.B(n_1684),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1688),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1703),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1739),
.A2(n_1706),
.B(n_1703),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1717),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1736),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1723),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1736),
.Y(n_1757)
);

AOI21xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1715),
.A2(n_1616),
.B(n_1607),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1736),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1717),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1727),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1751),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1737),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1730),
.B(n_1692),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1727),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1729),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1733),
.B(n_1712),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1729),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1740),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1751),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1733),
.B(n_1710),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1741),
.A2(n_1701),
.B1(n_1709),
.B2(n_1687),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1751),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1742),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1719),
.B(n_1710),
.Y(n_1775)
);

AND2x4_ASAP7_75t_SL g1776 ( 
.A(n_1744),
.B(n_1679),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1719),
.B(n_1728),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1742),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1780)
);

NAND4xp75_ASAP7_75t_L g1781 ( 
.A(n_1716),
.B(n_1701),
.C(n_1687),
.D(n_1659),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1730),
.B(n_1692),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1784)
);

OAI31xp33_ASAP7_75t_L g1785 ( 
.A1(n_1741),
.A2(n_1614),
.A3(n_1617),
.B(n_1649),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1749),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1716),
.B(n_1714),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1750),
.B(n_1666),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1738),
.B(n_1743),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1738),
.B(n_1692),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1734),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1746),
.B(n_1667),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1760),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1756),
.B(n_1718),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1756),
.B(n_1718),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1776),
.B(n_1722),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1760),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1774),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1767),
.B(n_1743),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1774),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1789),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1772),
.B(n_1735),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1779),
.Y(n_1807)
);

NAND2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1788),
.B(n_1666),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1779),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1786),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_SL g1811 ( 
.A(n_1785),
.B(n_1725),
.C(n_1726),
.D(n_1731),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1786),
.Y(n_1812)
);

NAND2xp33_ASAP7_75t_SL g1813 ( 
.A(n_1781),
.B(n_1750),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1790),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1783),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1767),
.B(n_1732),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1763),
.B(n_1735),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1776),
.B(n_1722),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1781),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1783),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1776),
.B(n_1783),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1784),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1763),
.B(n_1748),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1790),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1785),
.A2(n_1740),
.B(n_1744),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1788),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1754),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1754),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1784),
.B(n_1722),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1784),
.B(n_1722),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1792),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1761),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1778),
.B(n_1748),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1787),
.B(n_1744),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1813),
.A2(n_1758),
.B(n_1752),
.Y(n_1835)
);

OAI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1819),
.A2(n_1758),
.B1(n_1793),
.B2(n_1666),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1834),
.B(n_1787),
.Y(n_1837)
);

OAI322xp33_ASAP7_75t_L g1838 ( 
.A1(n_1819),
.A2(n_1782),
.A3(n_1764),
.B1(n_1793),
.B2(n_1765),
.C1(n_1766),
.C2(n_1761),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1811),
.A2(n_1777),
.B(n_1752),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1801),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1806),
.B(n_1787),
.Y(n_1841)
);

NOR4xp25_ASAP7_75t_SL g1842 ( 
.A(n_1797),
.B(n_1765),
.C(n_1766),
.D(n_1768),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1817),
.B(n_1791),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1802),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1823),
.A2(n_1740),
.B1(n_1793),
.B2(n_1744),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1797),
.Y(n_1846)
);

NAND5xp2_ASAP7_75t_L g1847 ( 
.A(n_1825),
.B(n_1777),
.C(n_1752),
.D(n_1780),
.E(n_1740),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1808),
.Y(n_1848)
);

AOI222xp33_ASAP7_75t_L g1849 ( 
.A1(n_1798),
.A2(n_1777),
.B1(n_1780),
.B2(n_1792),
.C1(n_1724),
.C2(n_1725),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1804),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1834),
.B(n_1821),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1799),
.A2(n_1780),
.B(n_1771),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1821),
.B(n_1800),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1800),
.B(n_1791),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1826),
.A2(n_1768),
.B(n_1796),
.Y(n_1856)
);

OAI321xp33_ASAP7_75t_L g1857 ( 
.A1(n_1808),
.A2(n_1764),
.A3(n_1782),
.B1(n_1771),
.B2(n_1794),
.C(n_1791),
.Y(n_1857)
);

AOI222xp33_ASAP7_75t_L g1858 ( 
.A1(n_1805),
.A2(n_1731),
.B1(n_1726),
.B2(n_1725),
.C1(n_1795),
.C2(n_1683),
.Y(n_1858)
);

AOI21xp33_ASAP7_75t_SL g1859 ( 
.A1(n_1808),
.A2(n_1831),
.B(n_1832),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1833),
.B(n_1764),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1826),
.A2(n_1769),
.B(n_1782),
.C(n_1794),
.Y(n_1861)
);

NAND2x1p5_ASAP7_75t_L g1862 ( 
.A(n_1840),
.B(n_1818),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1840),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1835),
.A2(n_1818),
.B(n_1815),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1846),
.Y(n_1865)
);

OAI211xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1861),
.A2(n_1827),
.B(n_1828),
.C(n_1807),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1852),
.B(n_1815),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1852),
.B(n_1820),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1841),
.B(n_1803),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1854),
.B(n_1820),
.Y(n_1870)
);

AO21x1_ASAP7_75t_L g1871 ( 
.A1(n_1846),
.A2(n_1828),
.B(n_1827),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1839),
.A2(n_1822),
.B(n_1829),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1844),
.Y(n_1873)
);

OAI321xp33_ASAP7_75t_L g1874 ( 
.A1(n_1836),
.A2(n_1822),
.A3(n_1803),
.B1(n_1829),
.B2(n_1830),
.C(n_1816),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1850),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1851),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1854),
.Y(n_1877)
);

OAI32xp33_ASAP7_75t_L g1878 ( 
.A1(n_1856),
.A2(n_1769),
.A3(n_1816),
.B1(n_1830),
.B2(n_1814),
.Y(n_1878)
);

AOI21xp33_ASAP7_75t_L g1879 ( 
.A1(n_1857),
.A2(n_1807),
.B(n_1804),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1855),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1837),
.B(n_1795),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1837),
.Y(n_1882)
);

AOI21xp33_ASAP7_75t_L g1883 ( 
.A1(n_1878),
.A2(n_1859),
.B(n_1848),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1880),
.A2(n_1877),
.B1(n_1868),
.B2(n_1867),
.Y(n_1884)
);

OAI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1882),
.A2(n_1847),
.B(n_1843),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1870),
.B(n_1855),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1863),
.B(n_1838),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1870),
.B(n_1867),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1871),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1862),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1871),
.Y(n_1891)
);

AOI322xp5_ASAP7_75t_L g1892 ( 
.A1(n_1879),
.A2(n_1842),
.A3(n_1726),
.B1(n_1731),
.B2(n_1795),
.C1(n_1747),
.C2(n_1745),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1874),
.A2(n_1853),
.B(n_1849),
.Y(n_1893)
);

NOR4xp25_ASAP7_75t_L g1894 ( 
.A(n_1889),
.B(n_1866),
.C(n_1865),
.D(n_1875),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1888),
.B(n_1880),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1888),
.Y(n_1896)
);

NAND3xp33_ASAP7_75t_SL g1897 ( 
.A(n_1893),
.B(n_1862),
.C(n_1864),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1890),
.B(n_1868),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1884),
.Y(n_1899)
);

AOI211xp5_ASAP7_75t_L g1900 ( 
.A1(n_1887),
.A2(n_1872),
.B(n_1845),
.C(n_1876),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_L g1901 ( 
.A(n_1887),
.B(n_1876),
.C(n_1873),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1886),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1891),
.A2(n_1869),
.B(n_1881),
.Y(n_1903)
);

OAI21xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1894),
.A2(n_1883),
.B(n_1892),
.Y(n_1904)
);

NAND4xp25_ASAP7_75t_L g1905 ( 
.A(n_1900),
.B(n_1885),
.C(n_1858),
.D(n_1860),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1896),
.Y(n_1906)
);

INVxp67_ASAP7_75t_L g1907 ( 
.A(n_1898),
.Y(n_1907)
);

NAND2x1_ASAP7_75t_L g1908 ( 
.A(n_1902),
.B(n_1809),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_SL g1909 ( 
.A1(n_1897),
.A2(n_1860),
.B(n_1810),
.C(n_1824),
.Y(n_1909)
);

AOI222xp33_ASAP7_75t_L g1910 ( 
.A1(n_1904),
.A2(n_1901),
.B1(n_1899),
.B2(n_1895),
.C1(n_1903),
.C2(n_1824),
.Y(n_1910)
);

O2A1O1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1909),
.A2(n_1814),
.B(n_1812),
.C(n_1810),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1905),
.A2(n_1907),
.B1(n_1906),
.B2(n_1908),
.C(n_1812),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1909),
.B(n_1809),
.Y(n_1913)
);

AOI221x1_ASAP7_75t_L g1914 ( 
.A1(n_1906),
.A2(n_1769),
.B1(n_1794),
.B2(n_1796),
.C(n_1759),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1904),
.A2(n_1769),
.B1(n_1773),
.B2(n_1770),
.C(n_1755),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1909),
.B(n_1796),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1916),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1913),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1910),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1915),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1912),
.B(n_1775),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1914),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1917),
.A2(n_1631),
.B1(n_1796),
.B2(n_1637),
.Y(n_1923)
);

NAND4xp75_ASAP7_75t_L g1924 ( 
.A(n_1919),
.B(n_1911),
.C(n_1753),
.D(n_1745),
.Y(n_1924)
);

NOR3xp33_ASAP7_75t_L g1925 ( 
.A(n_1918),
.B(n_1608),
.C(n_1658),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1918),
.B(n_1796),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1926),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_1925),
.B1(n_1923),
.B2(n_1919),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1928),
.A2(n_1919),
.B1(n_1921),
.B2(n_1920),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1928),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1930),
.A2(n_1920),
.B1(n_1922),
.B2(n_1924),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1929),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1931),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1932),
.A2(n_1746),
.B1(n_1753),
.B2(n_1757),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1933),
.A2(n_1757),
.B(n_1755),
.Y(n_1935)
);

AO21x2_ASAP7_75t_L g1936 ( 
.A1(n_1935),
.A2(n_1934),
.B(n_1757),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1936),
.A2(n_1762),
.B1(n_1755),
.B2(n_1759),
.C(n_1773),
.Y(n_1937)
);

OAI221xp5_ASAP7_75t_R g1938 ( 
.A1(n_1937),
.A2(n_1759),
.B1(n_1762),
.B2(n_1773),
.C(n_1770),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1938),
.A2(n_1658),
.B(n_1762),
.C(n_1770),
.Y(n_1939)
);


endmodule