module fake_jpeg_22733_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_21),
.Y(n_42)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_28),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_21),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_52),
.B(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_57),
.B1(n_20),
.B2(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_53),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_63),
.B(n_75),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_57),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_19),
.B(n_39),
.C(n_33),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_70),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_33),
.B1(n_41),
.B2(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_50),
.B1(n_52),
.B2(n_49),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_72),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_54),
.B1(n_51),
.B2(n_44),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_38),
.B1(n_35),
.B2(n_2),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_59),
.C(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_56),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_51),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_89),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_38),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_90),
.B1(n_66),
.B2(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_49),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_35),
.B1(n_44),
.B2(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_25),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_97),
.B(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_95),
.B1(n_76),
.B2(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_43),
.B1(n_33),
.B2(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_25),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_66),
.B(n_56),
.C(n_70),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_105),
.B1(n_117),
.B2(n_83),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_108),
.B1(n_109),
.B2(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_96),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_79),
.B1(n_78),
.B2(n_69),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_87),
.B1(n_80),
.B2(n_97),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_76),
.B(n_64),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_113),
.B(n_94),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_78),
.B(n_54),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_78),
.B1(n_46),
.B2(n_72),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_86),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_2),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_46),
.B(n_71),
.C(n_0),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_122),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_85),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_92),
.C(n_100),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_133),
.C(n_134),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_132),
.B(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_106),
.B1(n_117),
.B2(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_93),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_84),
.C(n_93),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_93),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_98),
.C(n_46),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_137),
.C(n_114),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_1),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_115),
.B(n_117),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_110),
.C(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_144),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_126),
.C(n_113),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_152),
.B1(n_25),
.B2(n_4),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_104),
.C(n_106),
.Y(n_149)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_117),
.B(n_136),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_151),
.B(n_154),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_111),
.B(n_117),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_102),
.B1(n_120),
.B2(n_117),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_159),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_154),
.C(n_148),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_128),
.B(n_134),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_161),
.B(n_164),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_162),
.C(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_113),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_163),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_142),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_150),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_143),
.B(n_153),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_3),
.B(n_5),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_167),
.B1(n_166),
.B2(n_164),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_153),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_144),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.C(n_158),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_148),
.C(n_4),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_177),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_183),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_182),
.C(n_3),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_166),
.C(n_155),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_167),
.B1(n_155),
.B2(n_6),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_173),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_9),
.B(n_10),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_8),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_193),
.B1(n_12),
.B2(n_13),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_201),
.B(n_198),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_10),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

OAI211xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_198),
.B(n_13),
.C(n_14),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_10),
.Y(n_206)
);


endmodule