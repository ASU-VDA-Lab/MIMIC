module fake_ariane_2897_n_333 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_333);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_333;

wire n_295;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_124;
wire n_119;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_183;
wire n_299;
wire n_133;
wire n_205;
wire n_109;
wire n_245;
wire n_319;
wire n_283;
wire n_187;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_189;
wire n_286;
wire n_117;
wire n_139;
wire n_130;
wire n_214;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_327;
wire n_279;
wire n_207;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_320;
wire n_309;
wire n_115;
wire n_331;
wire n_267;
wire n_291;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_128;
wire n_224;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_108;
wire n_303;
wire n_168;
wire n_206;
wire n_238;
wire n_136;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_104;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_221;
wire n_321;
wire n_149;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_287;
wire n_302;
wire n_284;
wire n_249;
wire n_123;
wire n_212;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_150;
wire n_113;
wire n_114;
wire n_324;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_246;
wire n_159;
wire n_105;
wire n_131;
wire n_263;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_258;
wire n_121;
wire n_118;
wire n_241;
wire n_191;
wire n_211;
wire n_322;
wire n_251;
wire n_116;
wire n_155;
wire n_127;

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_39),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_15),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_61),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_5),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_57),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_20),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_72),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_65),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_41),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_53),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_35),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_47),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_31),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_44),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_40),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_18),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_36),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_49),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_37),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_50),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_0),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_106),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_0),
.B(n_1),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_2),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_134),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_128),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_147),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_108),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_132),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_160),
.B1(n_134),
.B2(n_132),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_178),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_160),
.B1(n_147),
.B2(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_128),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_159),
.C(n_130),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_164),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_156),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_169),
.B(n_104),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_131),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NAND2x1p5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_135),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_139),
.C(n_137),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_136),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_140),
.B(n_141),
.C(n_152),
.Y(n_216)
);

AND3x2_ASAP7_75t_SL g217 ( 
.A(n_190),
.B(n_154),
.C(n_146),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_203),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_143),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_111),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_144),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_113),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_145),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_150),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

BUFx4f_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_192),
.A2(n_151),
.B1(n_120),
.B2(n_122),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_142),
.B(n_149),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_199),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_187),
.B1(n_108),
.B2(n_138),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_232),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_153),
.B(n_133),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_187),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_233),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_7),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_124),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_119),
.B1(n_118),
.B2(n_115),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_218),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_225),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_216),
.B1(n_210),
.B2(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_103),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_14),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_258),
.B(n_252),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_235),
.B(n_231),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_231),
.B(n_228),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_265),
.B(n_257),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_223),
.B(n_246),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_225),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_226),
.B(n_17),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_226),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_217),
.B(n_19),
.Y(n_279)
);

OAI211xp5_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_16),
.B(n_22),
.C(n_24),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_28),
.B(n_29),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_R g284 ( 
.A(n_248),
.B(n_100),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_253),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_259),
.B1(n_260),
.B2(n_250),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx5_ASAP7_75t_SL g288 ( 
.A(n_274),
.Y(n_288)
);

AOI221xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_241),
.B1(n_251),
.B2(n_254),
.C(n_38),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_269),
.B(n_268),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

AOI221xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_254),
.B1(n_32),
.B2(n_33),
.C(n_43),
.Y(n_293)
);

AOI221xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.C(n_48),
.Y(n_294)
);

AO31x2_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_281),
.A3(n_283),
.B(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_278),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_282),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_276),
.B1(n_273),
.B2(n_284),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_287),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_277),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_294),
.C(n_289),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_293),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

AND4x1_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_289),
.C(n_280),
.D(n_295),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

OAI33xp33_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_295),
.A3(n_51),
.B1(n_52),
.B2(n_62),
.B3(n_63),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_68),
.Y(n_321)
);

AO22x1_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_318),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_317),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

NAND4xp25_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_312),
.C(n_309),
.D(n_315),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_71),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_74),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

AOI222xp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.C1(n_80),
.C2(n_81),
.Y(n_331)
);

AO21x2_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_91),
.B(n_95),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_333)
);


endmodule