module fake_jpeg_15578_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_48),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_24),
.B1(n_22),
.B2(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_47),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_22),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_84)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_29),
.B1(n_33),
.B2(n_30),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_63),
.B1(n_68),
.B2(n_21),
.Y(n_89)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_15),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_30),
.B1(n_36),
.B2(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_69),
.Y(n_73)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_36),
.B1(n_31),
.B2(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_45),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_81),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_38),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_56),
.B(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_21),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_52),
.B1(n_65),
.B2(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_12),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_53),
.B1(n_20),
.B2(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_0),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_105),
.B(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_15),
.B(n_20),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_88),
.B1(n_74),
.B2(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_127),
.Y(n_140)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_89),
.B1(n_81),
.B2(n_75),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_115),
.B1(n_118),
.B2(n_97),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_108),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_75),
.B1(n_80),
.B2(n_83),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_75),
.B1(n_73),
.B2(n_52),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_85),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_97),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_90),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_105),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_23),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_87),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_107),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_102),
.B(n_100),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_132),
.B(n_141),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_115),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_143),
.B1(n_137),
.B2(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_103),
.B1(n_88),
.B2(n_55),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_74),
.B(n_76),
.C(n_55),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_76),
.B(n_23),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_151),
.B(n_49),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_79),
.Y(n_148)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_118),
.Y(n_167)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_55),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_113),
.B1(n_117),
.B2(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_174),
.B1(n_176),
.B2(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_122),
.C(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_134),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_114),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_49),
.Y(n_195)
);

NAND2x1_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_130),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_174),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_61),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_151),
.Y(n_180)
);

HB1xp67_ASAP7_75t_SL g172 ( 
.A(n_139),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_175),
.B(n_151),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_145),
.B1(n_144),
.B2(n_135),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_66),
.B1(n_64),
.B2(n_55),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_64),
.B1(n_17),
.B2(n_14),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_149),
.C(n_142),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_194),
.C(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_189),
.B1(n_196),
.B2(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_150),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_141),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_146),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_49),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_49),
.C(n_43),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_67),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_158),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_213),
.C(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_197),
.A2(n_162),
.B1(n_177),
.B2(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_205),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_162),
.B1(n_165),
.B2(n_160),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_168),
.B1(n_184),
.B2(n_159),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_0),
.B(n_1),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_165),
.B1(n_161),
.B2(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_40),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_175),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_67),
.C(n_40),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_211),
.B(n_184),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_219),
.B(n_224),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_227),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_191),
.B(n_193),
.C(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_195),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.C(n_201),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_11),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_237),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_214),
.C(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_206),
.B1(n_213),
.B2(n_203),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_203),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_236),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_10),
.B(n_17),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_17),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_34),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_230),
.B1(n_232),
.B2(n_229),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_249),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_219),
.B1(n_222),
.B2(n_17),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_238),
.A2(n_219),
.B1(n_10),
.B2(n_6),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_219),
.B(n_5),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_235),
.B(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_233),
.C(n_35),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_23),
.B(n_5),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_35),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_4),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_247),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_243),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_261),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_247),
.C(n_248),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_6),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_263),
.A2(n_255),
.B1(n_258),
.B2(n_8),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_8),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_260),
.A3(n_261),
.B1(n_8),
.B2(n_9),
.C1(n_6),
.C2(n_7),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_269),
.A2(n_266),
.B(n_264),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_35),
.C(n_9),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_35),
.Y(n_273)
);


endmodule