module real_jpeg_23135_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_1),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_119),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_119),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_1),
.A2(n_67),
.B1(n_68),
.B2(n_119),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_67),
.B1(n_68),
.B2(n_84),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_45),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_33),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_107),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_68),
.C(n_80),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_57),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_3),
.A2(n_65),
.B1(n_234),
.B2(n_241),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_5),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_5),
.A2(n_43),
.B1(n_67),
.B2(n_68),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_8),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_8),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_8),
.A2(n_26),
.B1(n_67),
.B2(n_68),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_51),
.B1(n_67),
.B2(n_68),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_12),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_155)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_20),
.B(n_120),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_90),
.C(n_102),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_21),
.B(n_90),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_24),
.B(n_47),
.C(n_63),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_42),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_118),
.Y(n_117)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_30),
.B(n_35),
.C(n_37),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_31),
.A2(n_42),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_31),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_32),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_32),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_158)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_35),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_34),
.A2(n_38),
.B(n_106),
.C(n_108),
.Y(n_105)
);

HAxp5_ASAP7_75t_SL g190 ( 
.A(n_34),
.B(n_107),
.CON(n_190),
.SN(n_190)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_35),
.A2(n_56),
.A3(n_59),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_46),
.B(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_60),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_50),
.B(n_57),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_52),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_52),
.A2(n_115),
.B1(n_140),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_52),
.A2(n_140),
.B1(n_157),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_53),
.B(n_61),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_53),
.A2(n_57),
.B1(n_181),
.B2(n_190),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AO22x1_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_55),
.B(n_58),
.Y(n_191)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_59),
.B1(n_80),
.B2(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_59),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_64),
.B(n_78),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_74),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_128),
.B(n_130),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_65),
.A2(n_74),
.B(n_130),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_65),
.A2(n_93),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_65),
.A2(n_128),
.B1(n_231),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_66),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_68),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_67),
.B(n_245),
.Y(n_244)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_77),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B(n_85),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_79),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_79),
.B(n_107),
.Y(n_239)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_100),
.B(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_125),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_86),
.A2(n_99),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_86),
.A2(n_196),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_86),
.A2(n_99),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_86),
.A2(n_99),
.B1(n_195),
.B2(n_216),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_101),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_101),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_96),
.A2(n_112),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_102),
.A2(n_103),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.C(n_117),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_107),
.B(n_128),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_118),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_145),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_131),
.B1(n_143),
.B2(n_144),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_142),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_182),
.B(n_260),
.C(n_265),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_168),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_168),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_165),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_163),
.B2(n_164),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_151),
.B(n_164),
.C(n_165),
.Y(n_261)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_169),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_172),
.B(n_174),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_201),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_255),
.B(n_259),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_210),
.B(n_254),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_187),
.B(n_197),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.C(n_194),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_192),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_193),
.B(n_194),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_205),
.C(n_209),
.Y(n_256)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_249),
.B(n_253),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_227),
.B(n_248),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_219),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_219),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_237),
.B(n_247),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_236),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_246),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);


endmodule