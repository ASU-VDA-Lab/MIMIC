module fake_netlist_1_7118_n_750 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_750);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_750;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_165;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_716;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_16), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_18), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_38), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_6), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_4), .Y(n_84) );
INVxp33_ASAP7_75t_L g85 ( .A(n_53), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_19), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_71), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_40), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_56), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_17), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_76), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_65), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_58), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_8), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_17), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_35), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_72), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_14), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_78), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_31), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_29), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_14), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_5), .B(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_55), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_62), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_3), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_16), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_51), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_75), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_0), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_24), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_68), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_85), .B(n_0), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_123), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_103), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_103), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
INVx2_ASAP7_75t_SL g136 ( .A(n_120), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_97), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_106), .B(n_1), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_111), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_111), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_82), .B(n_1), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
CKINVDCx11_ASAP7_75t_R g144 ( .A(n_79), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_123), .B(n_2), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_82), .B(n_2), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
OR2x2_ASAP7_75t_L g148 ( .A(n_84), .B(n_4), .Y(n_148) );
NAND2xp33_ASAP7_75t_L g149 ( .A(n_107), .B(n_42), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_128), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
BUFx8_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_88), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_108), .B(n_5), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_90), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_125), .B(n_6), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_107), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_84), .B(n_7), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_86), .B(n_7), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_90), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_107), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_86), .B(n_8), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_91), .B(n_9), .Y(n_167) );
INVxp67_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_107), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_92), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_92), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_93), .B(n_116), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_93), .B(n_9), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_160), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_172), .B(n_116), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_130), .B(n_110), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_130), .B(n_98), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_168), .B(n_102), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_162), .A2(n_102), .B1(n_122), .B2(n_105), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_166), .B(n_105), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_168), .B(n_99), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_141), .B(n_113), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_171), .B(n_113), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_141), .B(n_112), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_163), .B(n_112), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_143), .B(n_114), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_150), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_172), .B(n_80), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_129), .B(n_122), .Y(n_205) );
BUFx4f_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_129), .B(n_119), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_155), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_137), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_129), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_148), .A2(n_126), .B1(n_109), .B2(n_96), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_138), .B(n_158), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_172), .B(n_118), .Y(n_213) );
AND2x6_ASAP7_75t_L g214 ( .A(n_173), .B(n_114), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_138), .B(n_110), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_163), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_173), .B(n_115), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_173), .B(n_115), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_131), .Y(n_221) );
AND2x4_ASAP7_75t_SL g222 ( .A(n_138), .B(n_104), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_144), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_158), .B(n_104), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_143), .B(n_94), .Y(n_226) );
INVx8_ASAP7_75t_L g227 ( .A(n_145), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_145), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_131), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_173), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_131), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_131), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_151), .B(n_94), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_166), .Y(n_237) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_171), .B(n_95), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_166), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_152), .B(n_95), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_177), .B(n_148), .Y(n_243) );
CKINVDCx11_ASAP7_75t_R g244 ( .A(n_224), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_188), .Y(n_245) );
BUFx12f_ASAP7_75t_SL g246 ( .A(n_177), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_185), .A2(n_154), .B1(n_152), .B2(n_171), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_207), .B(n_155), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_188), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g250 ( .A(n_208), .B(n_155), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_185), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_208), .B(n_155), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_185), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_222), .B(n_148), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_210), .A2(n_136), .B1(n_154), .B2(n_146), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
CKINVDCx8_ASAP7_75t_R g260 ( .A(n_204), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_184), .B(n_142), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_240), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_240), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_222), .B(n_142), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_240), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_212), .B(n_146), .Y(n_266) );
INVx4_ASAP7_75t_SL g267 ( .A(n_196), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
NOR2xp33_ASAP7_75t_R g269 ( .A(n_209), .B(n_144), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_241), .Y(n_270) );
NAND2xp33_ASAP7_75t_L g271 ( .A(n_196), .B(n_214), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
AO22x1_ASAP7_75t_L g273 ( .A1(n_196), .A2(n_167), .B1(n_124), .B2(n_100), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_218), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_229), .B(n_153), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_202), .B(n_167), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_205), .B(n_157), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_218), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_220), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_220), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_183), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_194), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_225), .B(n_171), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_215), .B(n_170), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_196), .B(n_170), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_201), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_220), .B(n_170), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_238), .B(n_136), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_196), .B(n_157), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_214), .B(n_157), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_206), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_214), .B(n_159), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_182), .B(n_164), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_174), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_181), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_211), .A2(n_136), .B1(n_164), .B2(n_156), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_179), .B(n_156), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_214), .B(n_159), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_201), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_189), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_201), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_206), .Y(n_306) );
BUFx4f_ASAP7_75t_SL g307 ( .A(n_209), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_214), .B(n_159), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_190), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_193), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_238), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_179), .B(n_156), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_199), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_203), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_206), .B(n_216), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_266), .B(n_217), .Y(n_317) );
BUFx8_ASAP7_75t_SL g318 ( .A(n_258), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_303), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_246), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_248), .A2(n_195), .B(n_198), .C(n_226), .Y(n_321) );
AND2x6_ASAP7_75t_L g322 ( .A(n_303), .B(n_232), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_243), .B(n_236), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_277), .B(n_235), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_259), .Y(n_325) );
CKINVDCx11_ASAP7_75t_R g326 ( .A(n_260), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_309), .B(n_191), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_284), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_261), .B(n_242), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_300), .A2(n_176), .B1(n_230), .B2(n_226), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_274), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_254), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_275), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_300), .B(n_192), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_250), .A2(n_176), .B(n_230), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_279), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_254), .B(n_176), .Y(n_340) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_283), .B(n_191), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_282), .A2(n_198), .B1(n_195), .B2(n_239), .C(n_192), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_243), .B(n_176), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_309), .B(n_230), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_250), .A2(n_230), .B(n_239), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_264), .B(n_127), .Y(n_347) );
AOI21x1_ASAP7_75t_L g348 ( .A1(n_273), .A2(n_231), .B(n_233), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_278), .B(n_164), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_244), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_254), .B(n_153), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
BUFx12f_ASAP7_75t_L g353 ( .A(n_256), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_245), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_269), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_305), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_289), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_262), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_278), .B(n_153), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_280), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_281), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_311), .Y(n_362) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_264), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_249), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_286), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_307), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_307), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_267), .B(n_132), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_286), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_267), .B(n_132), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_293), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_267), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_251), .A2(n_140), .B1(n_139), .B2(n_135), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_263), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_328), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_365), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_369), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_363), .A2(n_253), .B1(n_247), .B2(n_255), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_374), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_374), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_319), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_319), .Y(n_384) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_326), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_333), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_SL g387 ( .A1(n_321), .A2(n_252), .B(n_248), .C(n_287), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_324), .B(n_247), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_324), .A2(n_272), .B1(n_268), .B2(n_270), .C(n_329), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_338), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_363), .A2(n_306), .B1(n_289), .B2(n_295), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_353), .A2(n_276), .B1(n_271), .B2(n_295), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_364), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_327), .A2(n_304), .B1(n_276), .B2(n_313), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_321), .A2(n_304), .B(n_316), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_352), .B(n_306), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_360), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_325), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_329), .A2(n_257), .B1(n_298), .B2(n_285), .C(n_299), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_323), .B(n_296), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_323), .B(n_297), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_348), .A2(n_301), .B(n_291), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_341), .B(n_310), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_336), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_341), .B(n_314), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_317), .A2(n_315), .B1(n_311), .B2(n_294), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_388), .B(n_357), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_389), .A2(n_318), .B1(n_353), .B2(n_326), .Y(n_411) );
OAI211xp5_ASAP7_75t_L g412 ( .A1(n_400), .A2(n_347), .B(n_366), .C(n_367), .Y(n_412) );
BUFx4f_ASAP7_75t_SL g413 ( .A(n_385), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_388), .A2(n_318), .B1(n_357), .B2(n_344), .Y(n_414) );
NOR4xp25_ASAP7_75t_L g415 ( .A(n_376), .B(n_124), .C(n_100), .D(n_121), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_375), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_376), .B(n_357), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_406), .A2(n_357), .B1(n_344), .B2(n_343), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_387), .A2(n_337), .B(n_346), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_349), .B1(n_354), .B2(n_357), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_380), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_377), .B(n_359), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_403), .A2(n_355), .B1(n_320), .B2(n_373), .C(n_330), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
OAI22xp33_ASAP7_75t_SL g425 ( .A1(n_378), .A2(n_350), .B1(n_355), .B2(n_351), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_393), .B(n_351), .Y(n_426) );
AO31x2_ASAP7_75t_L g427 ( .A1(n_395), .A2(n_140), .A3(n_132), .B(n_135), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_381), .Y(n_429) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_385), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_403), .A2(n_350), .B1(n_345), .B2(n_135), .C(n_139), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_375), .A2(n_335), .B1(n_332), .B2(n_339), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
OAI31xp33_ASAP7_75t_SL g434 ( .A1(n_393), .A2(n_370), .A3(n_368), .B(n_340), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_377), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_409), .A2(n_290), .B(n_358), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_406), .A2(n_322), .B1(n_371), .B2(n_356), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_379), .A2(n_322), .B1(n_371), .B2(n_356), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_421), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_421), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_426), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_435), .B(n_382), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_416), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_424), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_412), .A2(n_418), .B1(n_414), .B2(n_423), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_428), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_428), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_411), .B(n_385), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_429), .B(n_401), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g452 ( .A1(n_434), .A2(n_408), .B(n_392), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_415), .A2(n_391), .B(n_378), .C(n_398), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_420), .A2(n_402), .B1(n_407), .B2(n_405), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_438), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_429), .B(n_405), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_433), .B(n_407), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_431), .A2(n_386), .B1(n_399), .B2(n_398), .C(n_397), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_435), .B(n_117), .C(n_382), .D(n_397), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_425), .A2(n_399), .B1(n_390), .B2(n_386), .C(n_140), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_433), .B(n_390), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_425), .A2(n_396), .B1(n_322), .B2(n_384), .Y(n_462) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_419), .A2(n_404), .B(n_139), .Y(n_463) );
BUFx4f_ASAP7_75t_L g464 ( .A(n_426), .Y(n_464) );
OAI33xp33_ASAP7_75t_L g465 ( .A1(n_432), .A2(n_101), .A3(n_118), .B1(n_121), .B2(n_265), .B3(n_233), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_438), .B(n_383), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_430), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_410), .A2(n_396), .B1(n_322), .B2(n_368), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_439), .A2(n_101), .B1(n_356), .B2(n_291), .C(n_292), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_410), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_422), .B(n_383), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_437), .A2(n_396), .B1(n_342), .B2(n_292), .C(n_294), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_436), .B(n_149), .C(n_134), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_448), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_440), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_471), .B(n_427), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_442), .B(n_427), .Y(n_480) );
OAI33xp33_ASAP7_75t_L g481 ( .A1(n_459), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_15), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g482 ( .A1(n_450), .A2(n_413), .B1(n_430), .B2(n_396), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_459), .B(n_149), .C(n_169), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_440), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_447), .A2(n_335), .B1(n_332), .B2(n_362), .C(n_312), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_441), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_447), .B(n_368), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_448), .Y(n_489) );
NAND4xp25_ASAP7_75t_SL g490 ( .A(n_462), .B(n_11), .C(n_12), .D(n_13), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_468), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g492 ( .A1(n_465), .A2(n_332), .B(n_370), .C(n_340), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_452), .A2(n_322), .B1(n_383), .B2(n_384), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_471), .B(n_427), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g495 ( .A1(n_452), .A2(n_134), .B(n_161), .C(n_165), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
NAND2xp33_ASAP7_75t_SL g497 ( .A(n_454), .B(n_372), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_467), .B(n_427), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_472), .B(n_384), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_458), .A2(n_322), .B1(n_133), .B2(n_147), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_458), .A2(n_335), .B1(n_334), .B2(n_319), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_456), .B(n_18), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_460), .B(n_169), .C(n_131), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_472), .B(n_20), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g507 ( .A(n_453), .B(n_372), .C(n_301), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_476), .B(n_169), .C(n_133), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_443), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_464), .A2(n_335), .B1(n_334), .B2(n_319), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_451), .B(n_20), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_442), .B(n_370), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_451), .B(n_169), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_446), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_169), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_446), .B(n_169), .C(n_133), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_464), .A2(n_319), .B1(n_334), .B2(n_362), .Y(n_518) );
OAI31xp33_ASAP7_75t_L g519 ( .A1(n_454), .A2(n_340), .A3(n_362), .B(n_287), .Y(n_519) );
OAI31xp33_ASAP7_75t_L g520 ( .A1(n_470), .A2(n_308), .A3(n_342), .B(n_134), .Y(n_520) );
AOI21xp5_ASAP7_75t_SL g521 ( .A1(n_457), .A2(n_470), .B(n_449), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_475), .A2(n_334), .B1(n_308), .B2(n_372), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_442), .B(n_334), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_449), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_449), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_457), .B(n_131), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_461), .B(n_131), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_444), .B(n_131), .Y(n_529) );
OAI222xp33_ASAP7_75t_L g530 ( .A1(n_511), .A2(n_444), .B1(n_473), .B2(n_469), .C1(n_474), .C2(n_455), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_479), .B(n_474), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_480), .B(n_517), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_477), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_480), .B(n_474), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_480), .B(n_455), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_496), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_524), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_494), .B(n_455), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_484), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_511), .B(n_473), .Y(n_542) );
INVxp67_ASAP7_75t_L g543 ( .A(n_524), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_523), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_487), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_497), .B(n_464), .Y(n_546) );
INVx4_ASAP7_75t_L g547 ( .A(n_512), .Y(n_547) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_490), .B(n_466), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_506), .B(n_464), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_501), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_506), .B(n_475), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_509), .B(n_463), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_485), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_514), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_485), .Y(n_556) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_488), .B(n_165), .C(n_161), .D(n_134), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_483), .B(n_169), .C(n_147), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_481), .A2(n_134), .B1(n_161), .B2(n_165), .C(n_133), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_489), .B(n_463), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_525), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_491), .Y(n_563) );
NOR2xp67_ASAP7_75t_L g564 ( .A(n_507), .B(n_147), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_525), .B(n_463), .Y(n_565) );
INVx5_ASAP7_75t_L g566 ( .A(n_513), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_482), .B(n_23), .Y(n_567) );
NOR3xp33_ASAP7_75t_SL g568 ( .A(n_488), .B(n_25), .C(n_30), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_526), .B(n_463), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_526), .B(n_133), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_515), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_515), .B(n_133), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_499), .B(n_133), .Y(n_574) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_502), .A2(n_404), .B(n_231), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_513), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_504), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_521), .B(n_161), .C(n_165), .D(n_178), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_497), .A2(n_161), .B(n_165), .C(n_133), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_529), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_528), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_521), .B(n_147), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_512), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_512), .B(n_147), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_493), .B(n_147), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_492), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_493), .Y(n_591) );
AOI22xp5_ASAP7_75t_SL g592 ( .A1(n_577), .A2(n_518), .B1(n_519), .B2(n_495), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_540), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_571), .B(n_500), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_540), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_537), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_531), .B(n_500), .Y(n_597) );
CKINVDCx16_ASAP7_75t_R g598 ( .A(n_563), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_541), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_566), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_578), .A2(n_486), .B(n_520), .C(n_505), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_541), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_544), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_531), .B(n_522), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_545), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_554), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_571), .B(n_147), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_590), .A2(n_508), .B(n_200), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_590), .A2(n_200), .B(n_228), .Y(n_609) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_547), .B(n_147), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_566), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_536), .B(n_32), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_538), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_545), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_532), .B(n_169), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_530), .A2(n_543), .B(n_546), .C(n_567), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_554), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_550), .B(n_187), .Y(n_619) );
NAND4xp25_ASAP7_75t_SL g620 ( .A(n_548), .B(n_33), .C(n_34), .D(n_37), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_552), .Y(n_621) );
CKINVDCx16_ASAP7_75t_R g622 ( .A(n_547), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_538), .B(n_228), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_564), .A2(n_178), .B(n_197), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_532), .B(n_39), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_586), .B(n_43), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_544), .B(n_44), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_581), .B(n_219), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_555), .B(n_187), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_555), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_581), .B(n_219), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_535), .B(n_46), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_553), .B(n_187), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_560), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_535), .Y(n_636) );
NAND2xp33_ASAP7_75t_R g637 ( .A(n_568), .B(n_47), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_560), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_574), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_542), .B(n_197), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_585), .A2(n_49), .B(n_50), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_582), .B(n_583), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_551), .A2(n_234), .B1(n_221), .B2(n_187), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_582), .B(n_52), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_553), .B(n_186), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_547), .B(n_54), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_616), .A2(n_588), .B1(n_591), .B2(n_534), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_610), .A2(n_579), .B(n_588), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_613), .B(n_580), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_642), .B(n_580), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_593), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_595), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_596), .B(n_591), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_599), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_603), .B(n_583), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_647), .B(n_534), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_615), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_598), .B(n_557), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_602), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_636), .B(n_569), .Y(n_661) );
AO22x2_ASAP7_75t_L g662 ( .A1(n_605), .A2(n_533), .B1(n_539), .B2(n_556), .Y(n_662) );
INVx4_ASAP7_75t_L g663 ( .A(n_622), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_639), .B(n_572), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_600), .B(n_539), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_604), .B(n_606), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_614), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_618), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_617), .B(n_621), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_625), .B(n_572), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_631), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_635), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_611), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_638), .B(n_576), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_612), .B(n_587), .Y(n_675) );
AOI31xp33_ASAP7_75t_L g676 ( .A1(n_592), .A2(n_646), .A3(n_641), .B(n_601), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_594), .B(n_576), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_594), .B(n_569), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_626), .B(n_566), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_607), .B(n_561), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_607), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_634), .B(n_561), .Y(n_682) );
NOR2x1p5_ASAP7_75t_SL g683 ( .A(n_644), .B(n_584), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_597), .B(n_562), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_634), .B(n_565), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_645), .B(n_562), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_633), .B(n_566), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_628), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_620), .A2(n_585), .B(n_589), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_619), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_641), .A2(n_559), .B(n_549), .C(n_566), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_637), .A2(n_566), .B1(n_573), .B2(n_589), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_609), .A2(n_584), .B1(n_573), .B2(n_565), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_640), .A2(n_570), .B(n_556), .Y(n_694) );
AO21x1_ASAP7_75t_L g695 ( .A1(n_643), .A2(n_533), .B(n_575), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_619), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_630), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_630), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_645), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_627), .A2(n_558), .B1(n_570), .B2(n_575), .Y(n_700) );
OAI322xp33_ASAP7_75t_L g701 ( .A1(n_632), .A2(n_186), .A3(n_180), .B1(n_63), .B2(n_64), .C1(n_66), .C2(n_69), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_609), .B(n_186), .C(n_180), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_623), .B(n_186), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g704 ( .A1(n_643), .A2(n_180), .B(n_234), .C(n_221), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_629), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_608), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_608), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_624), .B(n_180), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_636), .B(n_57), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_616), .A2(n_61), .B1(n_70), .B2(n_73), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_642), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_648), .B(n_678), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_676), .A2(n_659), .B(n_683), .C(n_689), .Y(n_713) );
AOI211x1_ASAP7_75t_SL g714 ( .A1(n_654), .A2(n_656), .B(n_691), .C(n_649), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_663), .A2(n_679), .B(n_708), .Y(n_715) );
OAI22xp33_ASAP7_75t_SL g716 ( .A1(n_663), .A2(n_679), .B1(n_673), .B2(n_711), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_651), .A2(n_663), .B1(n_658), .B2(n_678), .C(n_659), .Y(n_717) );
AOI311xp33_ASAP7_75t_L g718 ( .A1(n_699), .A2(n_694), .A3(n_675), .B(n_705), .C(n_652), .Y(n_718) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_710), .A2(n_692), .B(n_693), .C(n_675), .Y(n_719) );
OAI31xp33_ASAP7_75t_L g720 ( .A1(n_688), .A2(n_662), .A3(n_665), .B(n_709), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_696), .B(n_698), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_693), .A2(n_706), .B(n_677), .C(n_684), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_661), .B(n_668), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_662), .Y(n_724) );
XNOR2xp5_ASAP7_75t_L g725 ( .A(n_666), .B(n_657), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_708), .A2(n_662), .B(n_695), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_721), .Y(n_727) );
AOI31xp33_ASAP7_75t_L g728 ( .A1(n_713), .A2(n_706), .A3(n_704), .B(n_700), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_718), .A2(n_665), .B1(n_702), .B2(n_650), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g730 ( .A1(n_716), .A2(n_664), .B(n_669), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_723), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_720), .B(n_661), .Y(n_732) );
AOI221xp5_ASAP7_75t_SL g733 ( .A1(n_717), .A2(n_669), .B1(n_655), .B2(n_671), .C(n_653), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g734 ( .A1(n_712), .A2(n_680), .B(n_697), .Y(n_734) );
OAI221xp5_ASAP7_75t_L g735 ( .A1(n_714), .A2(n_660), .B1(n_667), .B2(n_690), .C(n_672), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_727), .B(n_722), .Y(n_736) );
INVxp33_ASAP7_75t_SL g737 ( .A(n_729), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_728), .B(n_719), .C(n_726), .Y(n_738) );
NAND4xp25_ASAP7_75t_SL g739 ( .A(n_733), .B(n_715), .C(n_726), .D(n_687), .Y(n_739) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_730), .B(n_701), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_738), .A2(n_732), .B1(n_734), .B2(n_735), .Y(n_741) );
AOI222xp33_ASAP7_75t_L g742 ( .A1(n_737), .A2(n_736), .B1(n_740), .B2(n_732), .C1(n_724), .C2(n_739), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_738), .A2(n_731), .B1(n_725), .B2(n_681), .Y(n_743) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_742), .A2(n_731), .B1(n_665), .B2(n_707), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_743), .B(n_703), .C(n_670), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_745), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g747 ( .A1(n_744), .A2(n_741), .B1(n_674), .B2(n_686), .C(n_680), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_746), .A2(n_682), .B(n_685), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_748), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_749), .A2(n_747), .B(n_682), .Y(n_750) );
endmodule