module real_jpeg_30661_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_0),
.Y(n_255)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_0),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_1),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_69),
.B1(n_99),
.B2(n_103),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_69),
.B1(n_219),
.B2(n_224),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_1),
.A2(n_69),
.B1(n_342),
.B2(n_346),
.Y(n_341)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_3),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_3),
.A2(n_141),
.B1(n_287),
.B2(n_290),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_4),
.B(n_114),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g351 ( 
.A1(n_4),
.A2(n_352),
.A3(n_357),
.B1(n_359),
.B2(n_364),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_4),
.A2(n_190),
.B1(n_383),
.B2(n_386),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_4),
.A2(n_257),
.B(n_419),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_5),
.A2(n_63),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_5),
.A2(n_63),
.B1(n_375),
.B2(n_379),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_5),
.A2(n_63),
.B1(n_411),
.B2(n_415),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_6),
.A2(n_204),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_6),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_13),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_11),
.A2(n_248),
.B1(n_251),
.B2(n_253),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_11),
.Y(n_253)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_12),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_14),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_14),
.A2(n_109),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_14),
.A2(n_109),
.B1(n_368),
.B2(n_371),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_14),
.A2(n_109),
.B1(n_317),
.B2(n_464),
.Y(n_463)
);

AOI22x1_ASAP7_75t_L g206 ( 
.A1(n_15),
.A2(n_207),
.B1(n_213),
.B2(n_214),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_15),
.A2(n_213),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_15),
.A2(n_213),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_16),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_17),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_17),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_17),
.A2(n_132),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_299),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_258),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_173),
.C(n_233),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_25),
.A2(n_26),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_115),
.B1(n_116),
.B2(n_172),
.Y(n_26)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_75),
.B2(n_76),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_28),
.B(n_75),
.C(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_59),
.B(n_66),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_30),
.A2(n_184),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_30),
.A2(n_66),
.B(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_31),
.A2(n_176),
.B1(n_182),
.B2(n_183),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g314 ( 
.A(n_31),
.B(n_68),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_45),
.Y(n_31)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_35),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_36),
.Y(n_223)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_40),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_41),
.Y(n_245)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_50),
.B(n_53),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_48),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_49),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_49),
.Y(n_168)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_52),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_57),
.Y(n_388)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g385 ( 
.A(n_62),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_68),
.Y(n_268)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_73),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_74),
.Y(n_356)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_107),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_98),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_78),
.B(n_188),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_78),
.A2(n_108),
.B1(n_114),
.B2(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_95),
.Y(n_280)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_114),
.Y(n_186)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_104),
.Y(n_277)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_149),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_117),
.B(n_149),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_125),
.B1(n_137),
.B2(n_140),
.Y(n_117)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_118),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_118),
.B(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_118),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_120),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_121),
.Y(n_250)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_121),
.Y(n_467)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_124),
.Y(n_298)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_124),
.Y(n_421)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_126),
.A2(n_257),
.B1(n_316),
.B2(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_131),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_131),
.Y(n_345)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_135),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_136),
.Y(n_349)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_136),
.Y(n_418)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_145),
.Y(n_320)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_148),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_155),
.B1(n_161),
.B2(n_165),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_173),
.A2(n_174),
.B1(n_233),
.B2(n_234),
.Y(n_304)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_185),
.C(n_192),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_175),
.B(n_192),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_176),
.Y(n_313)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_179),
.Y(n_274)
);

BUFx4f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g312 ( 
.A1(n_184),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_184),
.B(n_190),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_185),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B(n_191),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_190),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_190),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_190),
.B(n_437),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_190),
.B(n_236),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_190),
.B(n_476),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_205),
.B1(n_218),
.B2(n_226),
.Y(n_192)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_193),
.B(n_218),
.Y(n_392)
);

AO22x2_ASAP7_75t_SL g406 ( 
.A1(n_193),
.A2(n_218),
.B1(n_226),
.B2(n_407),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_228),
.Y(n_227)
);

OAI22x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_200),
.B2(n_203),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_215),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_197),
.Y(n_446)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_227),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_211),
.Y(n_370)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_212),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_212),
.Y(n_438)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_217),
.Y(n_380)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_223),
.Y(n_291)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_223),
.Y(n_378)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI211xp5_ASAP7_75t_L g448 ( 
.A1(n_226),
.A2(n_449),
.B(n_450),
.C(n_451),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_227),
.A2(n_236),
.B1(n_237),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_227),
.A2(n_236),
.B1(n_367),
.B2(n_374),
.Y(n_366)
);

OAI21xp33_ASAP7_75t_SL g391 ( 
.A1(n_227),
.A2(n_374),
.B(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_245),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_247),
.A2(n_257),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_254),
.Y(n_480)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_SL g321 ( 
.A(n_255),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_257),
.A2(n_410),
.B(n_419),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_281),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_275),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx4f_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_292),
.B2(n_293),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_290),
.Y(n_450)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_324),
.B(n_494),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_303),
.Y(n_497)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_306),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_307),
.B(n_490),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_309),
.Y(n_491)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.C(n_322),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_312),
.B(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_315),
.A2(n_322),
.B1(n_323),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_316),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI21x1_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_485),
.B(n_492),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_399),
.B(n_484),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_389),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_330),
.B(n_389),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_366),
.C(n_381),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_350),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_351),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_340),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_338),
.Y(n_471)
);

OAI21xp33_ASAP7_75t_L g462 ( 
.A1(n_340),
.A2(n_463),
.B(n_468),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_381),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_367),
.Y(n_407)
);

BUFx4f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_396),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.Y(n_390)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_391),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_393),
.B(n_394),
.C(n_488),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_422),
.B(n_454),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_401),
.B(n_455),
.C(n_458),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_402),
.Y(n_424)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.C(n_409),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_408),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_453),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_410),
.Y(n_481)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx2_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_415),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_452),
.Y(n_422)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_425),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_447),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_447),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_435),
.B1(n_439),
.B2(n_440),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_437),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_452),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_478),
.C(n_482),
.Y(n_458)
);

OA21x2_ASAP7_75t_SL g459 ( 
.A1(n_460),
.A2(n_472),
.B(n_477),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_461),
.B(n_462),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_465),
.B(n_475),
.Y(n_474)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_469),
.Y(n_476)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_489),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_497),
.Y(n_495)
);


endmodule