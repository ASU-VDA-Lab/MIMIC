module fake_jpeg_16470_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_42),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_14),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_35),
.Y(n_106)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_54),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_29),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_24),
.B1(n_23),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_78),
.A2(n_83),
.B1(n_91),
.B2(n_94),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_79),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_96),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_40),
.A2(n_23),
.B1(n_33),
.B2(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_23),
.B1(n_65),
.B2(n_68),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_100),
.B1(n_115),
.B2(n_50),
.Y(n_129)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_36),
.B1(n_31),
.B2(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_28),
.B1(n_36),
.B2(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_38),
.B1(n_34),
.B2(n_18),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_99),
.B1(n_105),
.B2(n_111),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_39),
.A2(n_38),
.B1(n_34),
.B2(n_18),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_22),
.B1(n_34),
.B2(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_108),
.Y(n_125)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_35),
.B1(n_29),
.B2(n_22),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_22),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_3),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g114 ( 
.A(n_45),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_114),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_61),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_2),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_5),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_128),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_146),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_126),
.B(n_133),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_77),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_134),
.B1(n_161),
.B2(n_104),
.Y(n_185)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_73),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_80),
.A2(n_59),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_135),
.B(n_74),
.Y(n_206)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_89),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_140),
.B(n_154),
.Y(n_216)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_58),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_114),
.B(n_105),
.C(n_70),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_58),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_56),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_158),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_49),
.C(n_7),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_155),
.B1(n_119),
.B2(n_70),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_6),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_152),
.Y(n_215)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_7),
.Y(n_154)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_8),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_166),
.B1(n_13),
.B2(n_118),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_9),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_75),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_11),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_13),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_88),
.B(n_12),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_72),
.B(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_13),
.Y(n_168)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_75),
.B1(n_119),
.B2(n_98),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_185),
.B1(n_217),
.B2(n_218),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_193),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_165),
.B1(n_145),
.B2(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_186),
.A2(n_213),
.B1(n_212),
.B2(n_180),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_187),
.A2(n_182),
.B(n_191),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_125),
.B(n_85),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g195 ( 
.A1(n_145),
.A2(n_92),
.B1(n_74),
.B2(n_81),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_169),
.B(n_164),
.C(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_81),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_149),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_208),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_205),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_130),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_195),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_132),
.A2(n_92),
.B1(n_166),
.B2(n_157),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_214),
.B1(n_207),
.B2(n_215),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_136),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_139),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_165),
.A2(n_92),
.B1(n_160),
.B2(n_123),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_144),
.A2(n_166),
.B1(n_157),
.B2(n_164),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_150),
.A2(n_152),
.B1(n_132),
.B2(n_155),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_152),
.A2(n_132),
.B1(n_151),
.B2(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_225),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_146),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_232),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_223),
.A2(n_231),
.B(n_238),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_122),
.B1(n_163),
.B2(n_147),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_224),
.A2(n_234),
.B1(n_248),
.B2(n_192),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_135),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_235),
.C(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_229),
.B(n_236),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_124),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_186),
.A2(n_147),
.B1(n_162),
.B2(n_124),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_178),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_178),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_240),
.A2(n_244),
.B1(n_246),
.B2(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_201),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_242),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_173),
.B(n_177),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_187),
.A3(n_195),
.B1(n_211),
.B2(n_203),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_175),
.B(n_202),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g290 ( 
.A1(n_247),
.A2(n_255),
.B(n_231),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_172),
.B1(n_200),
.B2(n_199),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_190),
.B(n_172),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_254),
.Y(n_288)
);

NAND2x1_ASAP7_75t_SL g255 ( 
.A(n_208),
.B(n_191),
.Y(n_255)
);

XOR2x2_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_209),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_179),
.B(n_196),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_180),
.B(n_184),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_184),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_261),
.B(n_265),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_257),
.B1(n_255),
.B2(n_245),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_181),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_192),
.C(n_181),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_269),
.C(n_275),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_209),
.C(n_241),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_290),
.B(n_238),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_223),
.C(n_222),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_246),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_276),
.B(n_294),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_234),
.A2(n_227),
.B1(n_244),
.B2(n_251),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_278),
.A2(n_286),
.B1(n_290),
.B2(n_292),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_219),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_279),
.B(n_281),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_229),
.C(n_242),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_282),
.C(n_285),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_235),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_220),
.C(n_239),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_260),
.C(n_237),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_244),
.A2(n_231),
.B1(n_246),
.B2(n_253),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_219),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_287),
.B(n_228),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_300),
.B1(n_308),
.B2(n_313),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_302),
.B(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_221),
.Y(n_298)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_267),
.B1(n_290),
.B2(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_254),
.B1(n_236),
.B2(n_230),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_303),
.B(n_317),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_247),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_312),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_245),
.B1(n_230),
.B2(n_250),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_310),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_233),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_316),
.C(n_309),
.Y(n_339)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_250),
.B1(n_247),
.B2(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_315),
.Y(n_335)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_228),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_280),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_268),
.B(n_282),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_269),
.B1(n_294),
.B2(n_275),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_266),
.B(n_276),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_341),
.B(n_336),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_324),
.A2(n_334),
.B1(n_327),
.B2(n_344),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_336),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_265),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_339),
.C(n_340),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_270),
.B1(n_278),
.B2(n_286),
.Y(n_334)
);

AO22x1_ASAP7_75t_SL g336 ( 
.A1(n_297),
.A2(n_270),
.B1(n_271),
.B2(n_225),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_322),
.C(n_309),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_308),
.B1(n_313),
.B2(n_305),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_341),
.A2(n_295),
.B1(n_306),
.B2(n_304),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_322),
.C(n_311),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_344),
.C(n_312),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_300),
.C(n_307),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_345),
.A2(n_351),
.B1(n_362),
.B2(n_330),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_318),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_346),
.B(n_361),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_352),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_315),
.Y(n_350)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_331),
.A2(n_299),
.B1(n_337),
.B2(n_341),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_340),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_354),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_324),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_356),
.A2(n_362),
.B1(n_349),
.B2(n_345),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_323),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_359),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_342),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_325),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_335),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_335),
.Y(n_368)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_329),
.B(n_330),
.Y(n_362)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_374),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_371),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_348),
.B(n_332),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_356),
.C(n_357),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_359),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_354),
.C(n_347),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_379),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_347),
.C(n_352),
.Y(n_379)
);

AO21x1_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_374),
.B(n_368),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_383),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_376),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_358),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_378),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_387),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_382),
.A2(n_365),
.B(n_372),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_364),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_377),
.C(n_364),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_388),
.B(n_389),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_363),
.B1(n_365),
.B2(n_370),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_392),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_366),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_380),
.Y(n_395)
);


endmodule