module fake_jpeg_30653_n_203 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_11),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_22),
.Y(n_52)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_66),
.B1(n_77),
.B2(n_9),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_21),
.B(n_26),
.C(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_67),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_19),
.B1(n_30),
.B2(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_23),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_83),
.C(n_6),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_30),
.B1(n_23),
.B2(n_17),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_80),
.B(n_7),
.C(n_8),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_37),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_10),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_0),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_38),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_5),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_92),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

BUFx2_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_6),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_101),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_96),
.B(n_56),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_8),
.B1(n_51),
.B2(n_58),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_106),
.B1(n_66),
.B2(n_77),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_64),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_51),
.B1(n_54),
.B2(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_72),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_101),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_74),
.A3(n_73),
.B1(n_59),
.B2(n_68),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_68),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_103),
.CI(n_102),
.CON(n_127),
.SN(n_127)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_140),
.B(n_127),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_137),
.A2(n_141),
.B(n_121),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_113),
.B1(n_94),
.B2(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_129),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_87),
.B1(n_108),
.B2(n_107),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_88),
.C(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_92),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_96),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.C(n_124),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_156),
.B(n_134),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_142),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_157),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_114),
.B(n_112),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_131),
.B1(n_126),
.B2(n_125),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_137),
.B1(n_165),
.B2(n_161),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_132),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_134),
.B(n_147),
.C(n_149),
.D(n_135),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_146),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_136),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_172),
.C(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_174),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_167),
.Y(n_185)
);

OA21x2_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_162),
.B(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_156),
.C(n_152),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_166),
.B1(n_169),
.B2(n_173),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_179),
.B1(n_172),
.B2(n_148),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_165),
.B(n_158),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_190),
.B(n_178),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_144),
.B(n_163),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_189),
.B(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_187),
.B(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_185),
.B1(n_133),
.B2(n_135),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_195),
.Y(n_197)
);

OAI21x1_ASAP7_75t_SL g200 ( 
.A1(n_196),
.A2(n_195),
.B(n_193),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_177),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.C(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_122),
.Y(n_202)
);

XNOR2x2_ASAP7_75t_SL g203 ( 
.A(n_202),
.B(n_133),
.Y(n_203)
);


endmodule