module fake_netlist_1_9959_n_41 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
OAI22xp33_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_7), .B1(n_0), .B2(n_6), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_2), .B(n_11), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_2), .B(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_3), .B(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
BUFx2_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_6), .Y(n_18) );
AO22x1_ASAP7_75t_L g19 ( .A1(n_13), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
OAI21xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_13), .B(n_17), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_21), .B(n_17), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_23), .B(n_19), .Y(n_27) );
AOI211xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_12), .B(n_15), .C(n_14), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
OAI22xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_27), .B1(n_15), .B2(n_16), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_29), .B(n_27), .Y(n_31) );
OAI21xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_25), .B(n_28), .Y(n_32) );
AOI32xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_14), .A3(n_16), .B1(n_13), .B2(n_26), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
AOI21xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_13), .B(n_22), .Y(n_35) );
A2O1A1Ixp33_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_18), .B(n_24), .C(n_7), .Y(n_36) );
NOR2x1p5_ASAP7_75t_L g37 ( .A(n_32), .B(n_18), .Y(n_37) );
NOR2x1p5_ASAP7_75t_L g38 ( .A(n_37), .B(n_18), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_35), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_36), .B1(n_24), .B2(n_8), .Y(n_40) );
OAI31xp33_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_38), .A3(n_5), .B(n_8), .Y(n_41) );
endmodule