module fake_jpeg_16397_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_16),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_52),
.B1(n_22),
.B2(n_21),
.Y(n_66)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_36),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_29),
.Y(n_76)
);

AND2x4_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_24),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_33),
.B(n_37),
.C(n_32),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_64),
.B1(n_66),
.B2(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_67),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_75),
.B(n_76),
.Y(n_104)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_31),
.B(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_29),
.B1(n_16),
.B2(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_28),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_2),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_3),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_40),
.B1(n_51),
.B2(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_79),
.B1(n_52),
.B2(n_43),
.Y(n_95)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_78),
.Y(n_80)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_20),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_95),
.B1(n_19),
.B2(n_68),
.Y(n_115)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_89),
.Y(n_117)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_94),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_48),
.C(n_51),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_65),
.C(n_24),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_104),
.B(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_19),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_71),
.B1(n_79),
.B2(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_77),
.B1(n_60),
.B2(n_61),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_124),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_119),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_120),
.C(n_125),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_45),
.B1(n_68),
.B2(n_60),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_123),
.B1(n_96),
.B2(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_92),
.B1(n_97),
.B2(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_3),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_41),
.C(n_24),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_81),
.B1(n_84),
.B2(n_88),
.C(n_87),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_24),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_24),
.C(n_26),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_27),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_27),
.C(n_26),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_103),
.C(n_89),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_140),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_147),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_86),
.B1(n_84),
.B2(n_94),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_136),
.B1(n_149),
.B2(n_118),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_27),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_26),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_96),
.B(n_18),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_105),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_4),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_120),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_157),
.C(n_133),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_125),
.C(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_131),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_110),
.B1(n_116),
.B2(n_114),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_166),
.B1(n_143),
.B2(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_138),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_167),
.B(n_137),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_134),
.B1(n_132),
.B2(n_150),
.Y(n_178)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_144),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_182),
.C(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_180),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_139),
.B1(n_130),
.B2(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_154),
.B1(n_153),
.B2(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_183),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_142),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_141),
.C(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_165),
.Y(n_189)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_187),
.B1(n_192),
.B2(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_157),
.C(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_194),
.C(n_197),
.Y(n_198)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_118),
.B1(n_186),
.B2(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_152),
.C(n_159),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_161),
.C(n_170),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_180),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.C(n_203),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_171),
.C(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_177),
.C(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_140),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_189),
.B(n_196),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_203),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_191),
.B1(n_179),
.B2(n_176),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_198),
.B1(n_193),
.B2(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_219),
.C(n_212),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_126),
.B(n_14),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_111),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_199),
.C(n_149),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_210),
.B1(n_209),
.B2(n_135),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_222),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_214),
.C(n_8),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_226),
.B1(n_11),
.B2(n_13),
.Y(n_228)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

AOI31xp33_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_7),
.A3(n_11),
.B(n_12),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_227),
.B(n_13),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_13),
.Y(n_231)
);


endmodule