module real_aes_8122_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_1), .A2(n_152), .B(n_155), .C(n_158), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_2), .A2(n_178), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g538 ( .A(n_3), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_4), .B(n_201), .Y(n_224) );
AOI21xp33_ASAP7_75t_L g465 ( .A1(n_5), .A2(n_178), .B(n_466), .Y(n_465) );
AND2x6_ASAP7_75t_L g152 ( .A(n_6), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g185 ( .A(n_7), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_41), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_9), .A2(n_232), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_10), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g470 ( .A(n_11), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_12), .B(n_207), .Y(n_509) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g521 ( .A(n_14), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_15), .A2(n_186), .B(n_196), .C(n_199), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_16), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_17), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_18), .B(n_477), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_19), .B(n_178), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_20), .B(n_242), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_21), .A2(n_207), .B(n_208), .C(n_210), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_22), .B(n_201), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_23), .B(n_164), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_24), .A2(n_198), .B(n_199), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_25), .B(n_164), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_26), .Y(n_260) );
INVx1_ASAP7_75t_L g250 ( .A(n_27), .Y(n_250) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_28), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_29), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_30), .B(n_164), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_31), .A2(n_65), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_31), .Y(n_129) );
INVx1_ASAP7_75t_L g237 ( .A(n_32), .Y(n_237) );
INVx1_ASAP7_75t_L g459 ( .A(n_33), .Y(n_459) );
INVx2_ASAP7_75t_L g150 ( .A(n_34), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_35), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_36), .A2(n_207), .B(n_220), .C(n_222), .Y(n_219) );
INVxp67_ASAP7_75t_L g239 ( .A(n_37), .Y(n_239) );
CKINVDCx14_ASAP7_75t_R g218 ( .A(n_38), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_39), .A2(n_155), .B(n_249), .C(n_253), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_40), .A2(n_152), .B(n_155), .C(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g458 ( .A(n_42), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_43), .A2(n_166), .B(n_183), .C(n_184), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_44), .B(n_164), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_45), .A2(n_102), .B1(n_113), .B2(n_732), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_46), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_47), .Y(n_234) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_48), .A2(n_447), .B1(n_722), .B2(n_725), .C1(n_726), .C2(n_728), .Y(n_446) );
INVx1_ASAP7_75t_L g205 ( .A(n_49), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_50), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_51), .B(n_178), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_52), .A2(n_155), .B1(n_210), .B2(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_53), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_54), .Y(n_535) );
CKINVDCx14_ASAP7_75t_R g180 ( .A(n_55), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_56), .A2(n_183), .B(n_222), .C(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_57), .Y(n_501) );
INVx1_ASAP7_75t_L g467 ( .A(n_58), .Y(n_467) );
INVx1_ASAP7_75t_L g153 ( .A(n_59), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_60), .A2(n_78), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_60), .Y(n_724) );
INVx1_ASAP7_75t_L g143 ( .A(n_61), .Y(n_143) );
INVx1_ASAP7_75t_SL g221 ( .A(n_62), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_63), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_64), .B(n_201), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_65), .Y(n_128) );
INVx1_ASAP7_75t_L g263 ( .A(n_66), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_SL g476 ( .A1(n_67), .A2(n_222), .B(n_477), .C(n_478), .Y(n_476) );
INVxp67_ASAP7_75t_L g479 ( .A(n_68), .Y(n_479) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_70), .A2(n_178), .B(n_179), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_71), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_72), .A2(n_178), .B(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_73), .Y(n_462) );
INVx1_ASAP7_75t_L g495 ( .A(n_74), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_75), .A2(n_232), .B(n_233), .Y(n_231) );
INVx1_ASAP7_75t_L g194 ( .A(n_76), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_77), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_78), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_79), .A2(n_152), .B(n_155), .C(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_80), .A2(n_178), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g197 ( .A(n_81), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_82), .B(n_238), .Y(n_489) );
INVx2_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
INVx1_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_85), .B(n_477), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_86), .A2(n_152), .B(n_155), .C(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
OR2x2_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g721 ( .A(n_87), .B(n_123), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_88), .A2(n_155), .B(n_262), .C(n_265), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_89), .B(n_140), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_90), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_91), .A2(n_152), .B(n_155), .C(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_92), .Y(n_513) );
INVx1_ASAP7_75t_L g475 ( .A(n_93), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_94), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_95), .B(n_238), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_96), .B(n_171), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_97), .B(n_171), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g209 ( .A(n_99), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_100), .A2(n_178), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_104), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_111), .Y(n_105) );
OR2x2_ASAP7_75t_L g718 ( .A(n_107), .B(n_123), .Y(n_718) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_107), .B(n_122), .Y(n_730) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g123 ( .A(n_112), .B(n_124), .Y(n_123) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_445), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g731 ( .A(n_118), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_125), .B(n_442), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_121), .Y(n_444) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_130), .A2(n_448), .B1(n_716), .B2(n_719), .Y(n_447) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_131), .A2(n_716), .B1(n_721), .B2(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_397), .Y(n_131) );
NAND5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_309), .C(n_347), .D(n_368), .E(n_385), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_281), .C(n_302), .Y(n_133) );
OAI221xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_213), .B1(n_244), .B2(n_268), .C(n_272), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_173), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_137), .B(n_270), .Y(n_289) );
OR2x2_ASAP7_75t_L g316 ( .A(n_137), .B(n_190), .Y(n_316) );
AND2x2_ASAP7_75t_L g330 ( .A(n_137), .B(n_190), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_137), .B(n_176), .Y(n_344) );
AND2x2_ASAP7_75t_L g382 ( .A(n_137), .B(n_346), .Y(n_382) );
AND2x2_ASAP7_75t_L g411 ( .A(n_137), .B(n_321), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_137), .B(n_293), .Y(n_428) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g308 ( .A(n_138), .B(n_189), .Y(n_308) );
BUFx3_ASAP7_75t_L g333 ( .A(n_138), .Y(n_333) );
AND2x2_ASAP7_75t_L g362 ( .A(n_138), .B(n_190), .Y(n_362) );
AND3x2_ASAP7_75t_L g375 ( .A(n_138), .B(n_376), .C(n_377), .Y(n_375) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_168), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_139), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_139), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_139), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_140), .A2(n_177), .B(n_188), .Y(n_176) );
INVx2_ASAP7_75t_L g243 ( .A(n_140), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_140), .A2(n_147), .B(n_247), .C(n_248), .Y(n_246) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_140), .A2(n_516), .B(n_522), .Y(n_515) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g172 ( .A(n_141), .B(n_142), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_154), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_147), .A2(n_260), .B(n_261), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_147), .A2(n_187), .B1(n_456), .B2(n_460), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_147), .A2(n_495), .B(n_496), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_147), .A2(n_535), .B(n_536), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AND2x4_ASAP7_75t_L g178 ( .A(n_148), .B(n_152), .Y(n_178) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g240 ( .A(n_149), .Y(n_240) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
INVx3_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
INVx1_ASAP7_75t_L g477 ( .A(n_151), .Y(n_477) );
INVx4_ASAP7_75t_SL g187 ( .A(n_152), .Y(n_187) );
BUFx3_ASAP7_75t_L g253 ( .A(n_152), .Y(n_253) );
INVx5_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx3_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_156), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_163), .C(n_165), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_160), .A2(n_165), .B(n_263), .C(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_161), .A2(n_162), .B1(n_458), .B2(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx4_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
INVx2_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
INVx4_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_165), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_165), .A2(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx3_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_170), .B(n_255), .Y(n_254) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_170), .A2(n_259), .B(n_266), .Y(n_258) );
NOR2xp33_ASAP7_75t_SL g491 ( .A(n_170), .B(n_492), .Y(n_491) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_171), .A2(n_473), .B(n_480), .Y(n_472) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g230 ( .A(n_172), .Y(n_230) );
INVx1_ASAP7_75t_L g298 ( .A(n_173), .Y(n_298) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_189), .Y(n_173) );
AOI32xp33_ASAP7_75t_L g353 ( .A1(n_174), .A2(n_305), .A3(n_354), .B1(n_357), .B2(n_358), .Y(n_353) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g280 ( .A(n_175), .B(n_189), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_175), .B(n_308), .Y(n_351) );
AND2x2_ASAP7_75t_L g358 ( .A(n_175), .B(n_330), .Y(n_358) );
OR2x2_ASAP7_75t_L g364 ( .A(n_175), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_175), .B(n_319), .Y(n_389) );
OR2x2_ASAP7_75t_L g407 ( .A(n_175), .B(n_226), .Y(n_407) );
BUFx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g271 ( .A(n_176), .B(n_202), .Y(n_271) );
INVx2_ASAP7_75t_L g293 ( .A(n_176), .Y(n_293) );
OR2x2_ASAP7_75t_L g315 ( .A(n_176), .B(n_202), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_176), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_176), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g376 ( .A(n_176), .B(n_270), .Y(n_376) );
BUFx2_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_187), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_181), .A2(n_187), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_SL g204 ( .A1(n_181), .A2(n_187), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_181), .A2(n_187), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_181), .A2(n_187), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_181), .A2(n_187), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_181), .A2(n_187), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_181), .A2(n_187), .B(n_518), .C(n_519), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx5_ASAP7_75t_L g238 ( .A(n_186), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_186), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_186), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
INVx1_ASAP7_75t_SL g427 ( .A(n_189), .Y(n_427) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_202), .Y(n_189) );
INVx1_ASAP7_75t_SL g270 ( .A(n_190), .Y(n_270) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_190), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_190), .B(n_356), .Y(n_355) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_190), .B(n_293), .C(n_411), .Y(n_422) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_200), .Y(n_190) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_191), .A2(n_203), .B(n_212), .Y(n_202) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_191), .A2(n_216), .B(n_224), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_198), .B(n_209), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_198), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_198), .B(n_521), .Y(n_520) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_201), .A2(n_465), .B(n_471), .Y(n_464) );
INVx2_ASAP7_75t_L g321 ( .A(n_202), .Y(n_321) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_202), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_207), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g540 ( .A(n_210), .Y(n_540) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
INVx1_ASAP7_75t_L g357 ( .A(n_214), .Y(n_357) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g275 ( .A(n_215), .B(n_257), .Y(n_275) );
INVx2_ASAP7_75t_L g292 ( .A(n_215), .Y(n_292) );
AND2x2_ASAP7_75t_L g297 ( .A(n_215), .B(n_258), .Y(n_297) );
AND2x2_ASAP7_75t_L g312 ( .A(n_215), .B(n_245), .Y(n_312) );
AND2x2_ASAP7_75t_L g324 ( .A(n_215), .B(n_296), .Y(n_324) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_223), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_225), .B(n_340), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_225), .B(n_297), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_225), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_225), .B(n_291), .Y(n_419) );
BUFx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g256 ( .A(n_226), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_226), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g301 ( .A(n_226), .B(n_245), .Y(n_301) );
AND2x2_ASAP7_75t_L g327 ( .A(n_226), .B(n_257), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_226), .B(n_367), .Y(n_366) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_231), .B(n_241), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_228), .A2(n_286), .B(n_287), .Y(n_285) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_228), .A2(n_494), .B(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_SL g485 ( .A1(n_229), .A2(n_486), .B(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_230), .A2(n_455), .B(n_461), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_230), .B(n_462), .Y(n_461) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_230), .A2(n_534), .B(n_541), .Y(n_533) );
INVx1_ASAP7_75t_L g286 ( .A(n_231), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_236), .B(n_240), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_238), .A2(n_250), .B(n_251), .C(n_252), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_238), .A2(n_538), .B(n_539), .C(n_540), .Y(n_537) );
INVx2_ASAP7_75t_L g252 ( .A(n_240), .Y(n_252) );
INVx1_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_243), .B(n_267), .Y(n_266) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_243), .A2(n_505), .B(n_512), .Y(n_504) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_256), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_245), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g291 ( .A(n_245), .B(n_292), .Y(n_291) );
INVx3_ASAP7_75t_SL g296 ( .A(n_245), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_245), .B(n_283), .Y(n_349) );
OR2x2_ASAP7_75t_L g359 ( .A(n_245), .B(n_285), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_245), .B(n_327), .Y(n_387) );
OR2x2_ASAP7_75t_L g417 ( .A(n_245), .B(n_257), .Y(n_417) );
AND2x2_ASAP7_75t_L g421 ( .A(n_245), .B(n_258), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_245), .B(n_297), .Y(n_434) );
AND2x2_ASAP7_75t_L g441 ( .A(n_245), .B(n_323), .Y(n_441) );
OR2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
INVx1_ASAP7_75t_SL g384 ( .A(n_256), .Y(n_384) );
AND2x2_ASAP7_75t_L g323 ( .A(n_257), .B(n_285), .Y(n_323) );
AND2x2_ASAP7_75t_L g337 ( .A(n_257), .B(n_292), .Y(n_337) );
AND2x2_ASAP7_75t_L g340 ( .A(n_257), .B(n_296), .Y(n_340) );
INVx1_ASAP7_75t_L g367 ( .A(n_257), .Y(n_367) );
INVx2_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g279 ( .A(n_258), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_269), .A2(n_315), .B(n_439), .C(n_440), .Y(n_438) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g345 ( .A(n_270), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_271), .B(n_288), .Y(n_303) );
AND2x2_ASAP7_75t_L g329 ( .A(n_271), .B(n_330), .Y(n_329) );
OAI21xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_276), .B(n_280), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_274), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_275), .B(n_296), .Y(n_341) );
AND2x2_ASAP7_75t_L g432 ( .A(n_275), .B(n_283), .Y(n_432) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_279), .B(n_292), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_279), .B(n_290), .Y(n_306) );
OAI322xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_289), .A3(n_290), .B1(n_293), .B2(n_294), .C1(n_298), .C2(n_299), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
AND2x2_ASAP7_75t_L g393 ( .A(n_283), .B(n_305), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_283), .B(n_357), .Y(n_439) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g336 ( .A(n_285), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g402 ( .A(n_289), .B(n_315), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_290), .B(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_291), .B(n_323), .Y(n_380) );
AND2x2_ASAP7_75t_L g326 ( .A(n_292), .B(n_296), .Y(n_326) );
AND2x2_ASAP7_75t_L g334 ( .A(n_293), .B(n_335), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_293), .A2(n_372), .B(n_432), .C(n_433), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_294), .A2(n_307), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_296), .B(n_323), .Y(n_363) );
AND2x2_ASAP7_75t_L g369 ( .A(n_296), .B(n_337), .Y(n_369) );
AND2x2_ASAP7_75t_L g403 ( .A(n_296), .B(n_305), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_297), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_SL g413 ( .A(n_297), .Y(n_413) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_301), .A2(n_329), .B1(n_331), .B2(n_336), .Y(n_328) );
OAI22xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_304), .B1(n_306), .B2(n_307), .Y(n_302) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_303), .A2(n_339), .B1(n_341), .B2(n_342), .Y(n_338) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_308), .A2(n_410), .B1(n_412), .B2(n_414), .C(n_418), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B(n_317), .C(n_338), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
OR2x2_ASAP7_75t_L g379 ( .A(n_315), .B(n_332), .Y(n_379) );
INVx1_ASAP7_75t_L g430 ( .A(n_315), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g317 ( .A1(n_316), .A2(n_318), .B1(n_322), .B2(n_325), .C(n_328), .Y(n_317) );
INVx2_ASAP7_75t_SL g372 ( .A(n_316), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g437 ( .A(n_319), .Y(n_437) );
AND2x2_ASAP7_75t_L g361 ( .A(n_320), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g346 ( .A(n_321), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g408 ( .A(n_324), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_332), .B(n_434), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_336), .A2(n_348), .B(n_350), .C(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g425 ( .A(n_339), .Y(n_425) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_343), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g356 ( .A(n_346), .Y(n_356) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_359), .B1(n_360), .B2(n_363), .C1(n_364), .C2(n_366), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g392 ( .A(n_356), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_359), .B(n_413), .Y(n_412) );
NAND2xp33_ASAP7_75t_SL g390 ( .A(n_360), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g365 ( .A(n_362), .Y(n_365) );
AND2x2_ASAP7_75t_L g429 ( .A(n_362), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g395 ( .A(n_365), .B(n_392), .Y(n_395) );
INVx1_ASAP7_75t_L g424 ( .A(n_366), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_373), .C(n_378), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_372), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
AOI322xp5_ASAP7_75t_L g423 ( .A1(n_375), .A2(n_403), .A3(n_408), .B1(n_424), .B2(n_425), .C1(n_426), .C2(n_429), .Y(n_423) );
AND2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_411), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_381), .B2(n_383), .Y(n_378) );
INVxp33_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B1(n_390), .B2(n_393), .C(n_394), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND5xp2_ASAP7_75t_L g397 ( .A(n_398), .B(n_409), .C(n_423), .D(n_431), .E(n_435), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B(n_404), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp33_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_411), .A2(n_436), .B(n_437), .C(n_438), .Y(n_435) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_413), .A2(n_419), .A3(n_420), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g436 ( .A(n_434), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_442), .B(n_446), .C(n_731), .Y(n_445) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g727 ( .A(n_448), .Y(n_727) );
AND3x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_641), .C(n_690), .Y(n_448) );
NOR3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_548), .C(n_586), .Y(n_449) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_481), .B1(n_523), .B2(n_529), .C1(n_543), .C2(n_546), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_452), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_452), .B(n_591), .Y(n_682) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g559 ( .A(n_453), .B(n_472), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_453), .B(n_464), .Y(n_567) );
AND2x2_ASAP7_75t_L g602 ( .A(n_453), .B(n_579), .Y(n_602) );
OR2x2_ASAP7_75t_L g626 ( .A(n_453), .B(n_464), .Y(n_626) );
OR2x2_ASAP7_75t_L g634 ( .A(n_453), .B(n_533), .Y(n_634) );
AND2x2_ASAP7_75t_L g637 ( .A(n_453), .B(n_472), .Y(n_637) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g531 ( .A(n_454), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g545 ( .A(n_454), .B(n_472), .Y(n_545) );
AND2x2_ASAP7_75t_L g595 ( .A(n_454), .B(n_533), .Y(n_595) );
AND2x2_ASAP7_75t_L g608 ( .A(n_454), .B(n_464), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_454), .B(n_694), .Y(n_715) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_463), .A2(n_634), .B(n_635), .C(n_638), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_463), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_463), .B(n_578), .Y(n_700) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_472), .Y(n_463) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_464), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g558 ( .A(n_464), .Y(n_558) );
AND2x2_ASAP7_75t_L g585 ( .A(n_464), .B(n_579), .Y(n_585) );
INVx1_ASAP7_75t_SL g593 ( .A(n_464), .Y(n_593) );
AND2x2_ASAP7_75t_L g616 ( .A(n_464), .B(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g694 ( .A(n_464), .Y(n_694) );
BUFx2_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
INVx1_ASAP7_75t_L g592 ( .A(n_472), .Y(n_592) );
INVx3_ASAP7_75t_L g617 ( .A(n_472), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_481), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_502), .Y(n_481) );
INVx1_ASAP7_75t_L g613 ( .A(n_482), .Y(n_613) );
OAI32xp33_ASAP7_75t_L g619 ( .A1(n_482), .A2(n_558), .A3(n_620), .B1(n_621), .B2(n_622), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_482), .A2(n_624), .B1(n_627), .B2(n_632), .Y(n_623) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g561 ( .A(n_483), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g639 ( .A(n_483), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g709 ( .A(n_483), .B(n_655), .Y(n_709) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
AND2x2_ASAP7_75t_L g524 ( .A(n_484), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g554 ( .A(n_484), .Y(n_554) );
INVx1_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
OR2x2_ASAP7_75t_L g581 ( .A(n_484), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g588 ( .A(n_484), .B(n_562), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_484), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g609 ( .A(n_484), .B(n_527), .Y(n_609) );
INVx3_ASAP7_75t_L g631 ( .A(n_484), .Y(n_631) );
AND2x2_ASAP7_75t_L g656 ( .A(n_484), .B(n_528), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_484), .B(n_621), .Y(n_704) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
INVx2_ASAP7_75t_L g528 ( .A(n_493), .Y(n_528) );
AND2x2_ASAP7_75t_L g660 ( .A(n_493), .B(n_503), .Y(n_660) );
INVx2_ASAP7_75t_L g702 ( .A(n_502), .Y(n_702) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
INVx1_ASAP7_75t_L g547 ( .A(n_503), .Y(n_547) );
AND2x2_ASAP7_75t_L g574 ( .A(n_503), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_503), .B(n_528), .Y(n_582) );
AND2x2_ASAP7_75t_L g640 ( .A(n_503), .B(n_563), .Y(n_640) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g526 ( .A(n_504), .Y(n_526) );
AND2x2_ASAP7_75t_L g553 ( .A(n_504), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_504), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_504), .B(n_528), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_510), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_514), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g575 ( .A(n_514), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_514), .B(n_528), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_514), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g655 ( .A(n_514), .Y(n_655) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g527 ( .A(n_515), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g563 ( .A(n_515), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_523), .A2(n_533), .B1(n_692), .B2(n_695), .Y(n_691) );
INVx1_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_525), .A2(n_636), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_526), .B(n_631), .Y(n_648) );
INVx1_ASAP7_75t_L g673 ( .A(n_526), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_527), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_553), .Y(n_600) );
INVx2_ASAP7_75t_L g556 ( .A(n_528), .Y(n_556) );
INVx1_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_529), .A2(n_681), .B1(n_698), .B2(n_701), .C(n_703), .Y(n_697) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g568 ( .A(n_530), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_530), .B(n_579), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_531), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g622 ( .A(n_531), .B(n_568), .Y(n_622) );
INVx3_ASAP7_75t_SL g663 ( .A(n_531), .Y(n_663) );
AND2x2_ASAP7_75t_L g607 ( .A(n_532), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g636 ( .A(n_532), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_532), .B(n_545), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_532), .B(n_591), .Y(n_677) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g579 ( .A(n_533), .Y(n_579) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_533), .A2(n_605), .A3(n_627), .B1(n_675), .B2(n_677), .C1(n_678), .C2(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_544), .A2(n_547), .B(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_545), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g646 ( .A(n_545), .B(n_558), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_545), .B(n_585), .Y(n_661) );
INVxp67_ASAP7_75t_L g612 ( .A(n_547), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_547), .A2(n_619), .B(n_623), .C(n_633), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_557), .B1(n_560), .B2(n_564), .C(n_569), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g572 ( .A(n_556), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g689 ( .A(n_556), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_557), .A2(n_706), .B1(n_711), .B2(n_712), .C(n_714), .Y(n_705) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_558), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g605 ( .A(n_558), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_558), .B(n_636), .Y(n_643) );
AND2x2_ASAP7_75t_L g685 ( .A(n_558), .B(n_663), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_559), .B(n_584), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_559), .A2(n_571), .B1(n_681), .B2(n_682), .Y(n_680) );
OR2x2_ASAP7_75t_L g711 ( .A(n_559), .B(n_579), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g688 ( .A(n_562), .Y(n_688) );
AND2x2_ASAP7_75t_L g713 ( .A(n_562), .B(n_656), .Y(n_713) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_SL g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g577 ( .A(n_567), .B(n_578), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_576), .B1(n_580), .B2(n_583), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g644 ( .A(n_572), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_572), .B(n_612), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g603 ( .A1(n_574), .A2(n_604), .A3(n_606), .B1(n_607), .B2(n_609), .C1(n_610), .C2(n_614), .Y(n_603) );
INVxp67_ASAP7_75t_L g597 ( .A(n_575), .Y(n_597) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_577), .A2(n_582), .B1(n_599), .B2(n_601), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_578), .B(n_591), .Y(n_678) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_579), .B(n_617), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_579), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g675 ( .A(n_581), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
NAND3xp33_ASAP7_75t_SL g586 ( .A(n_587), .B(n_603), .C(n_618), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_594), .B2(n_596), .C(n_598), .Y(n_587) );
AND2x2_ASAP7_75t_L g594 ( .A(n_590), .B(n_595), .Y(n_594) );
INVx3_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g604 ( .A(n_595), .B(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_597), .Y(n_676) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_602), .B(n_616), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_605), .B(n_663), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_606), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g681 ( .A(n_609), .Y(n_681) );
AND2x2_ASAP7_75t_L g696 ( .A(n_609), .B(n_673), .Y(n_696) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_620), .A2(n_691), .B(n_697), .C(n_705), .Y(n_690) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g659 ( .A(n_630), .B(n_660), .Y(n_659) );
NAND2x1_ASAP7_75t_SL g701 ( .A(n_631), .B(n_702), .Y(n_701) );
CKINVDCx16_ASAP7_75t_R g671 ( .A(n_634), .Y(n_671) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g666 ( .A(n_640), .Y(n_666) );
AND2x2_ASAP7_75t_L g670 ( .A(n_640), .B(n_656), .Y(n_670) );
NOR5xp2_ASAP7_75t_L g641 ( .A(n_642), .B(n_657), .C(n_674), .D(n_680), .E(n_683), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_645), .B2(n_647), .C(n_649), .Y(n_642) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_646), .B(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g672 ( .A(n_656), .B(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_661), .B1(n_662), .B2(n_664), .C(n_667), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
AOI211xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_686), .B(n_688), .C(n_689), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
CKINVDCx14_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
CKINVDCx14_ASAP7_75t_R g725 ( .A(n_722), .Y(n_725) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx3_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
endmodule