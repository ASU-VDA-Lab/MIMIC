module fake_jpeg_22271_n_284 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_23),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_32),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_16),
.B1(n_23),
.B2(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_32),
.B1(n_39),
.B2(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_15),
.B1(n_22),
.B2(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_19),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_15),
.B1(n_25),
.B2(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NAND2xp67_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_32),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_61),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_35),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_32),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_82),
.C(n_54),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_32),
.B1(n_30),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_72),
.B1(n_73),
.B2(n_41),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_43),
.B1(n_45),
.B2(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_30),
.B(n_24),
.C(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2x1_ASAP7_75t_SL g82 ( 
.A(n_41),
.B(n_24),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_75),
.B1(n_73),
.B2(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_47),
.B1(n_55),
.B2(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_89),
.B1(n_72),
.B2(n_60),
.Y(n_112)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_58),
.B1(n_57),
.B2(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_42),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_82),
.B(n_37),
.Y(n_121)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_120),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_71),
.B(n_73),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_111),
.B(n_119),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_96),
.B1(n_89),
.B2(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_60),
.B1(n_53),
.B2(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_93),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_56),
.B(n_66),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_57),
.B1(n_58),
.B2(n_69),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_92),
.C(n_91),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_69),
.B1(n_53),
.B2(n_79),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_91),
.B1(n_41),
.B2(n_33),
.Y(n_153)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_69),
.B1(n_82),
.B2(n_40),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_128),
.B1(n_107),
.B2(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_79),
.Y(n_125)
);

XOR2x2_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_69),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_90),
.B(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_37),
.B1(n_34),
.B2(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_90),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_148),
.C(n_115),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_105),
.C(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_88),
.B(n_87),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_127),
.B(n_34),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_152),
.B1(n_153),
.B2(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_92),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_164),
.C(n_172),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_158),
.B1(n_165),
.B2(n_168),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_123),
.B1(n_111),
.B2(n_126),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_108),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_166),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_147),
.B1(n_144),
.B2(n_141),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_109),
.B(n_114),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_109),
.CI(n_117),
.CON(n_167),
.SN(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_131),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_127),
.B1(n_120),
.B2(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_175),
.B1(n_177),
.B2(n_134),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_106),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_149),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_77),
.C(n_62),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_24),
.C(n_26),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_100),
.B1(n_103),
.B2(n_40),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_40),
.B1(n_20),
.B2(n_17),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_183),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_190),
.B(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_132),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_130),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_139),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_143),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_137),
.B1(n_136),
.B2(n_98),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_200),
.B1(n_176),
.B2(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_178),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_172),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_158),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.C(n_199),
.Y(n_205)
);

AOI21x1_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_24),
.B(n_1),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_70),
.C(n_98),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_26),
.C(n_21),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_165),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_213),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_157),
.B(n_163),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_SL g235 ( 
.A(n_206),
.B(n_214),
.C(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_157),
.C(n_166),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_176),
.C(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_168),
.C(n_167),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_167),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_21),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_13),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_12),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_180),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_212),
.C(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_196),
.B1(n_197),
.B2(n_20),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_13),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_10),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_12),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_12),
.Y(n_241)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_9),
.Y(n_259)
);

OAI21x1_ASAP7_75t_SL g238 ( 
.A1(n_230),
.A2(n_203),
.B(n_213),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_225),
.B1(n_11),
.B2(n_10),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_205),
.B(n_212),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_221),
.B(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_242),
.C(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_248),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_218),
.C(n_1),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_0),
.C(n_1),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_11),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_255),
.B(n_257),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_231),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_253),
.B(n_0),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_235),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_228),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_11),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_9),
.C(n_2),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_246),
.C(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_0),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_244),
.B1(n_17),
.B2(n_4),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_0),
.C(n_3),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_4),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_4),
.B(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_262),
.B(n_263),
.Y(n_275)
);

AOI321xp33_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_260),
.A3(n_261),
.B1(n_266),
.B2(n_276),
.C(n_7),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_269),
.B(n_264),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_278),
.B(n_272),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_265),
.Y(n_278)
);

AOI222xp33_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_280),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_257),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_5),
.B(n_7),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_7),
.Y(n_284)
);


endmodule