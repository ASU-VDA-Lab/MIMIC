module real_aes_2657_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g512 ( .A(n_0), .B(n_209), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_1), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_2), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g143 ( .A(n_3), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_4), .B(n_515), .Y(n_534) );
NAND2xp33_ASAP7_75t_SL g505 ( .A(n_5), .B(n_164), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_6), .B(n_177), .Y(n_200) );
INVx1_ASAP7_75t_L g497 ( .A(n_7), .Y(n_497) );
INVx1_ASAP7_75t_L g234 ( .A(n_8), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g805 ( .A(n_9), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_10), .Y(n_251) );
AND2x2_ASAP7_75t_L g532 ( .A(n_11), .B(n_133), .Y(n_532) );
INVx2_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_13), .Y(n_110) );
INVx1_ASAP7_75t_L g210 ( .A(n_14), .Y(n_210) );
AOI221x1_ASAP7_75t_L g500 ( .A1(n_15), .A2(n_166), .B1(n_501), .B2(n_503), .C(n_504), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_16), .B(n_515), .Y(n_568) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g207 ( .A(n_18), .Y(n_207) );
INVx1_ASAP7_75t_SL g155 ( .A(n_19), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_20), .B(n_158), .Y(n_180) );
AOI33xp33_ASAP7_75t_L g225 ( .A1(n_21), .A2(n_49), .A3(n_140), .B1(n_151), .B2(n_226), .B3(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_22), .A2(n_503), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_23), .B(n_209), .Y(n_537) );
AOI221xp5_ASAP7_75t_SL g577 ( .A1(n_24), .A2(n_39), .B1(n_503), .B2(n_515), .C(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g244 ( .A(n_25), .Y(n_244) );
OR2x2_ASAP7_75t_L g135 ( .A(n_26), .B(n_88), .Y(n_135) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_26), .A2(n_88), .B(n_134), .Y(n_168) );
INVxp67_ASAP7_75t_L g499 ( .A(n_27), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_28), .B(n_212), .Y(n_572) );
AND2x2_ASAP7_75t_L g526 ( .A(n_29), .B(n_132), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_30), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_31), .A2(n_503), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_32), .B(n_212), .Y(n_579) );
AND2x2_ASAP7_75t_L g145 ( .A(n_33), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g150 ( .A(n_33), .Y(n_150) );
AND2x2_ASAP7_75t_L g164 ( .A(n_33), .B(n_143), .Y(n_164) );
OR2x6_ASAP7_75t_L g112 ( .A(n_34), .B(n_113), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_34), .B(n_804), .C(n_806), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_35), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_36), .B(n_138), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_37), .A2(n_167), .B1(n_173), .B2(n_177), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_38), .B(n_182), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_40), .A2(n_79), .B1(n_148), .B2(n_503), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_41), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_42), .B(n_209), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_43), .A2(n_779), .B1(n_781), .B2(n_783), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_44), .B(n_184), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_45), .B(n_158), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_46), .Y(n_176) );
AND2x2_ASAP7_75t_L g516 ( .A(n_47), .B(n_132), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_48), .B(n_132), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_50), .B(n_158), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_51), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_51), .A2(n_61), .B1(n_423), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g141 ( .A(n_52), .Y(n_141) );
INVx1_ASAP7_75t_L g160 ( .A(n_52), .Y(n_160) );
AND2x2_ASAP7_75t_L g276 ( .A(n_53), .B(n_132), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_54), .A2(n_72), .B1(n_138), .B2(n_148), .C(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_55), .B(n_138), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_56), .B(n_515), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_57), .B(n_167), .Y(n_253) );
AOI21xp5_ASAP7_75t_SL g189 ( .A1(n_58), .A2(n_148), .B(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g553 ( .A(n_59), .B(n_132), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_60), .B(n_212), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_61), .Y(n_798) );
INVx1_ASAP7_75t_L g203 ( .A(n_62), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_63), .B(n_209), .Y(n_551) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_64), .B(n_133), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_65), .A2(n_503), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g274 ( .A(n_66), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_67), .B(n_212), .Y(n_538) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_68), .B(n_184), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_69), .A2(n_148), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g146 ( .A(n_70), .Y(n_146) );
INVx1_ASAP7_75t_L g162 ( .A(n_70), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_71), .B(n_138), .Y(n_228) );
AND2x2_ASAP7_75t_L g165 ( .A(n_73), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g204 ( .A(n_74), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_75), .A2(n_148), .B(n_154), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_76), .A2(n_148), .B(n_179), .C(n_183), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_77), .A2(n_82), .B1(n_138), .B2(n_515), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_78), .B(n_515), .Y(n_552) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_80), .B(n_114), .Y(n_807) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_81), .B(n_166), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_83), .A2(n_148), .B1(n_223), .B2(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_84), .B(n_209), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_85), .B(n_209), .Y(n_580) );
INVxp33_ASAP7_75t_L g809 ( .A(n_86), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_87), .A2(n_503), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g191 ( .A(n_89), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_90), .B(n_212), .Y(n_550) );
AND2x2_ASAP7_75t_L g229 ( .A(n_91), .B(n_166), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_92), .A2(n_242), .B(n_243), .C(n_245), .Y(n_241) );
INVxp67_ASAP7_75t_L g502 ( .A(n_93), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_94), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_95), .B(n_212), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_96), .A2(n_503), .B(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g105 ( .A(n_97), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_98), .B(n_158), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_99), .Y(n_779) );
AOI21xp33_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_800), .B(n_808), .Y(n_100) );
OA21x2_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_117), .B(n_787), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_104), .B(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_107), .A2(n_789), .B(n_799), .Y(n_788) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_116), .Y(n_107) );
BUFx2_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g799 ( .A(n_109), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x6_ASAP7_75t_SL g487 ( .A(n_110), .B(n_112), .Y(n_487) );
OR2x6_ASAP7_75t_SL g778 ( .A(n_110), .B(n_111), .Y(n_778) );
OR2x2_ASAP7_75t_L g786 ( .A(n_110), .B(n_112), .Y(n_786) );
CKINVDCx16_ASAP7_75t_R g806 ( .A(n_110), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_779), .B(n_780), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_486), .B1(n_488), .B2(n_776), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_121), .A2(n_486), .B1(n_489), .B2(n_782), .Y(n_781) );
AND3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_480), .C(n_483), .Y(n_121) );
NAND5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_380), .C(n_410), .D(n_424), .E(n_450), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g480 ( .A1(n_124), .A2(n_423), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g794 ( .A(n_124), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_329), .Y(n_124) );
NOR3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_277), .C(n_311), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_194), .B(n_216), .C(n_255), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_169), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_129), .B(n_267), .Y(n_332) );
AND2x2_ASAP7_75t_L g419 ( .A(n_129), .B(n_197), .Y(n_419) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g215 ( .A(n_130), .B(n_186), .Y(n_215) );
INVx1_ASAP7_75t_L g257 ( .A(n_130), .Y(n_257) );
INVx2_ASAP7_75t_L g262 ( .A(n_130), .Y(n_262) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_130), .Y(n_290) );
INVx1_ASAP7_75t_L g304 ( .A(n_130), .Y(n_304) );
AND2x2_ASAP7_75t_L g308 ( .A(n_130), .B(n_199), .Y(n_308) );
AND2x2_ASAP7_75t_L g389 ( .A(n_130), .B(n_198), .Y(n_389) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_136), .B(n_165), .Y(n_130) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_131), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_131), .A2(n_547), .B(n_553), .Y(n_546) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_131), .A2(n_520), .B(n_526), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_132), .Y(n_131) );
OA21x2_ASAP7_75t_L g576 ( .A1(n_132), .A2(n_577), .B(n_581), .Y(n_576) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g177 ( .A(n_134), .B(n_135), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_147), .Y(n_136) );
INVx1_ASAP7_75t_L g254 ( .A(n_138), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_138), .A2(n_148), .B1(n_496), .B2(n_498), .Y(n_495) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
OR2x6_ASAP7_75t_L g156 ( .A(n_140), .B(n_152), .Y(n_156) );
INVxp33_ASAP7_75t_L g226 ( .A(n_140), .Y(n_226) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g153 ( .A(n_141), .B(n_143), .Y(n_153) );
AND2x4_ASAP7_75t_L g212 ( .A(n_141), .B(n_161), .Y(n_212) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g503 ( .A(n_145), .B(n_153), .Y(n_503) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
AND2x6_ASAP7_75t_L g209 ( .A(n_146), .B(n_159), .Y(n_209) );
INVxp67_ASAP7_75t_L g252 ( .A(n_148), .Y(n_252) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NOR2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx1_ASAP7_75t_L g227 ( .A(n_151), .Y(n_227) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_156), .B(n_157), .C(n_163), .Y(n_154) );
INVx2_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_156), .A2(n_163), .B(n_191), .C(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_156), .A2(n_163), .B(n_234), .C(n_235), .Y(n_233) );
INVxp67_ASAP7_75t_L g242 ( .A(n_156), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_156), .A2(n_163), .B(n_274), .C(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
AND2x4_ASAP7_75t_L g515 ( .A(n_158), .B(n_164), .Y(n_515) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_163), .A2(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_163), .B(n_177), .Y(n_213) );
INVx1_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_163), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_163), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_163), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_163), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_163), .A2(n_571), .B(n_572), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_163), .A2(n_579), .B(n_580), .Y(n_578) );
INVx5_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_164), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_166), .A2(n_241), .B1(n_246), .B2(n_247), .Y(n_240) );
INVx3_ASAP7_75t_L g247 ( .A(n_166), .Y(n_247) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_167), .B(n_250), .Y(n_249) );
AOI21x1_ASAP7_75t_L g508 ( .A1(n_167), .A2(n_509), .B(n_516), .Y(n_508) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_168), .Y(n_184) );
AND2x4_ASAP7_75t_SL g169 ( .A(n_170), .B(n_185), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g214 ( .A(n_171), .Y(n_214) );
AND2x2_ASAP7_75t_L g258 ( .A(n_171), .B(n_199), .Y(n_258) );
AND2x2_ASAP7_75t_L g279 ( .A(n_171), .B(n_186), .Y(n_279) );
INVx1_ASAP7_75t_L g302 ( .A(n_171), .Y(n_302) );
AND2x4_ASAP7_75t_L g369 ( .A(n_171), .B(n_198), .Y(n_369) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_178), .Y(n_171) );
NOR3xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .C(n_176), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_177), .A2(n_189), .B(n_193), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_177), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_177), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_177), .B(n_502), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_177), .B(n_205), .C(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_177), .A2(n_534), .B(n_535), .Y(n_533) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_183), .A2(n_221), .B(n_229), .Y(n_220) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_183), .A2(n_221), .B(n_229), .Y(n_284) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_183), .A2(n_542), .B(n_545), .Y(n_541) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_184), .A2(n_232), .B(n_236), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_184), .A2(n_568), .B(n_569), .Y(n_567) );
AND2x4_ASAP7_75t_L g385 ( .A(n_185), .B(n_302), .Y(n_385) );
OR2x2_ASAP7_75t_L g426 ( .A(n_185), .B(n_427), .Y(n_426) );
NOR2xp67_ASAP7_75t_SL g445 ( .A(n_185), .B(n_318), .Y(n_445) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_185), .B(n_377), .Y(n_463) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2x1_ASAP7_75t_SL g263 ( .A(n_186), .B(n_199), .Y(n_263) );
AND2x4_ASAP7_75t_L g301 ( .A(n_186), .B(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_186), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_186), .B(n_261), .Y(n_339) );
INVx2_ASAP7_75t_L g353 ( .A(n_186), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_186), .B(n_305), .Y(n_375) );
AND2x2_ASAP7_75t_L g467 ( .A(n_186), .B(n_325), .Y(n_467) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_L g195 ( .A(n_196), .B(n_215), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_197), .B(n_304), .Y(n_318) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_197), .B(n_307), .Y(n_327) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_214), .Y(n_197) );
INVx1_ASAP7_75t_L g305 ( .A(n_198), .Y(n_305) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g325 ( .A(n_199), .Y(n_325) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_206), .B(n_213), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_205), .B(n_244), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B1(n_210), .B2(n_211), .Y(n_206) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVxp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g358 ( .A(n_214), .Y(n_358) );
INVx2_ASAP7_75t_SL g403 ( .A(n_215), .Y(n_403) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_237), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_218), .B(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g349 ( .A(n_218), .Y(n_349) );
AND2x2_ASAP7_75t_L g473 ( .A(n_218), .B(n_298), .Y(n_473) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_230), .Y(n_218) );
AND2x4_ASAP7_75t_L g286 ( .A(n_219), .B(n_268), .Y(n_286) );
INVx1_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
AND2x2_ASAP7_75t_L g328 ( .A(n_219), .B(n_283), .Y(n_328) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_220), .B(n_231), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_220), .B(n_269), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_222), .B(n_228), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVxp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
AND2x4_ASAP7_75t_L g334 ( .A(n_231), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g346 ( .A(n_231), .Y(n_346) );
INVx1_ASAP7_75t_L g388 ( .A(n_231), .Y(n_388) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_231), .Y(n_400) );
AND2x2_ASAP7_75t_L g416 ( .A(n_231), .B(n_239), .Y(n_416) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g363 ( .A(n_238), .B(n_321), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_238), .Y(n_365) );
AND2x2_ASAP7_75t_L g386 ( .A(n_238), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x4_ASAP7_75t_L g265 ( .A(n_239), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g293 ( .A(n_239), .Y(n_293) );
INVx2_ASAP7_75t_L g299 ( .A(n_239), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_239), .B(n_269), .Y(n_314) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_248), .Y(n_239) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_247), .A2(n_270), .B(n_276), .Y(n_269) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_247), .A2(n_270), .B(n_276), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_252), .B1(n_253), .B2(n_254), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B(n_264), .Y(n_255) );
INVx1_ASAP7_75t_L g395 ( .A(n_256), .Y(n_395) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
AND2x2_ASAP7_75t_L g371 ( .A(n_258), .B(n_307), .Y(n_371) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g285 ( .A(n_260), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_260), .B(n_301), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_260), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_260), .B(n_385), .Y(n_392) );
AND2x2_ASAP7_75t_L g466 ( .A(n_260), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_261), .Y(n_454) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_262), .Y(n_374) );
AND2x2_ASAP7_75t_L g287 ( .A(n_263), .B(n_288), .Y(n_287) );
OAI21xp33_ASAP7_75t_L g475 ( .A1(n_263), .A2(n_476), .B(n_478), .Y(n_475) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx3_ASAP7_75t_L g361 ( .A(n_265), .Y(n_361) );
NAND2x1_ASAP7_75t_SL g405 ( .A(n_265), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_265), .B(n_286), .Y(n_408) );
AND2x2_ASAP7_75t_L g320 ( .A(n_267), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g457 ( .A(n_267), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g468 ( .A(n_267), .B(n_416), .Y(n_468) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_268), .B(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g399 ( .A(n_269), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
OAI21xp5_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_291), .B(n_294), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B1(n_286), .B2(n_287), .Y(n_278) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_279), .Y(n_336) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_285), .Y(n_280) );
AND2x2_ASAP7_75t_L g309 ( .A(n_281), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g415 ( .A(n_281), .B(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_281), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_281), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g298 ( .A(n_283), .B(n_299), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_283), .B(n_299), .Y(n_379) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_283), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g335 ( .A(n_284), .Y(n_335) );
AND2x2_ASAP7_75t_L g343 ( .A(n_284), .B(n_299), .Y(n_343) );
INVx1_ASAP7_75t_L g406 ( .A(n_284), .Y(n_406) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_289), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g436 ( .A(n_292), .B(n_321), .Y(n_436) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
AND2x2_ASAP7_75t_L g333 ( .A(n_293), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g421 ( .A(n_293), .B(n_328), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_300), .B1(n_306), .B2(n_309), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g429 ( .A(n_296), .B(n_430), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g459 ( .A(n_299), .B(n_346), .Y(n_459) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g326 ( .A(n_301), .Y(n_326) );
OAI21xp33_ASAP7_75t_SL g472 ( .A1(n_301), .A2(n_473), .B(n_474), .Y(n_472) );
AND2x4_ASAP7_75t_SL g303 ( .A(n_304), .B(n_305), .Y(n_303) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_304), .Y(n_462) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_SL g404 ( .A1(n_307), .A2(n_405), .B(n_407), .C(n_409), .Y(n_404) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_308), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g409 ( .A(n_308), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_308), .B(n_385), .Y(n_449) );
INVx1_ASAP7_75t_SL g316 ( .A(n_309), .Y(n_316) );
AND2x2_ASAP7_75t_L g397 ( .A(n_310), .B(n_334), .Y(n_397) );
INVx1_ASAP7_75t_L g442 ( .A(n_310), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_316), .B2(n_317), .C(n_319), .Y(n_311) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_312), .Y(n_431) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g479 ( .A(n_314), .B(n_322), .Y(n_479) );
OR2x2_ASAP7_75t_L g338 ( .A(n_315), .B(n_339), .Y(n_338) );
NOR2x1_ASAP7_75t_L g351 ( .A(n_315), .B(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_315), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g477 ( .A(n_315), .B(n_374), .Y(n_477) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI32xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .A3(n_326), .B1(n_327), .B2(n_328), .Y(n_319) );
INVx1_ASAP7_75t_L g340 ( .A(n_321), .Y(n_340) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_323), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g435 ( .A(n_324), .Y(n_435) );
OAI22xp33_ASAP7_75t_SL g417 ( .A1(n_326), .A2(n_418), .B1(n_420), .B2(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g448 ( .A(n_327), .Y(n_448) );
AOI211x1_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_336), .B(n_337), .C(n_354), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_331), .B(n_416), .Y(n_422) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g378 ( .A(n_334), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g444 ( .A(n_334), .Y(n_444) );
OAI222xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B1(n_341), .B2(n_347), .C1(n_348), .C2(n_350), .Y(n_337) );
INVxp67_ASAP7_75t_L g434 ( .A(n_338), .Y(n_434) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_342), .B(n_427), .Y(n_474) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g390 ( .A(n_343), .B(n_387), .Y(n_390) );
INVx3_ASAP7_75t_L g430 ( .A(n_345), .Y(n_430) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g368 ( .A(n_353), .B(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B1(n_362), .B2(n_367), .C(n_370), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_356), .A2(n_413), .B(n_415), .Y(n_412) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g366 ( .A(n_360), .Y(n_366) );
OR2x2_ASAP7_75t_L g470 ( .A(n_361), .B(n_406), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_364), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_367), .A2(n_396), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_368), .A2(n_440), .B(n_447), .Y(n_446) );
INVx4_ASAP7_75t_L g377 ( .A(n_369), .Y(n_377) );
OAI31xp33_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_372), .A3(n_376), .B(n_378), .Y(n_370) );
INVx1_ASAP7_75t_L g428 ( .A(n_372), .Y(n_428) );
NOR2x1_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g402 ( .A(n_377), .Y(n_402) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_393), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_381), .B(n_393), .C(n_412), .D(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_391), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_389), .B2(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g453 ( .A(n_385), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_386), .B(n_406), .Y(n_414) );
INVx1_ASAP7_75t_SL g427 ( .A(n_389), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_404), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_398), .B2(n_401), .Y(n_394) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_403), .A2(n_466), .B1(n_468), .B2(n_469), .Y(n_465) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_417), .C(n_423), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI21xp33_ASAP7_75t_L g483 ( .A1(n_423), .A2(n_484), .B(n_485), .Y(n_483) );
INVxp33_ASAP7_75t_L g484 ( .A(n_424), .Y(n_484) );
AND2x2_ASAP7_75t_L g793 ( .A(n_424), .B(n_450), .Y(n_793) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_425), .B(n_432), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_429), .B2(n_431), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_429), .A2(n_452), .B(n_455), .Y(n_451) );
INVx2_ASAP7_75t_L g439 ( .A(n_430), .Y(n_439) );
NAND3xp33_ASAP7_75t_SL g432 ( .A(n_433), .B(n_437), .C(n_446), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_443), .B2(n_445), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVxp33_ASAP7_75t_SL g485 ( .A(n_450), .Y(n_485) );
NOR3x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_464), .C(n_471), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g795 ( .A(n_481), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_653), .Y(n_489) );
NOR4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_596), .C(n_635), .D(n_642), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_517), .B1(n_554), .B2(n_563), .C(n_582), .Y(n_491) );
OR2x2_ASAP7_75t_L g726 ( .A(n_492), .B(n_588), .Y(n_726) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g641 ( .A(n_493), .B(n_566), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_493), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_SL g706 ( .A(n_493), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .Y(n_493) );
AND2x4_ASAP7_75t_SL g565 ( .A(n_494), .B(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g587 ( .A(n_494), .Y(n_587) );
AND2x2_ASAP7_75t_L g622 ( .A(n_494), .B(n_595), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_494), .B(n_507), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_494), .B(n_589), .Y(n_674) );
OR2x2_ASAP7_75t_L g752 ( .A(n_494), .B(n_566), .Y(n_752) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .Y(n_494) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g574 ( .A(n_507), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_507), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g600 ( .A(n_507), .Y(n_600) );
OR2x2_ASAP7_75t_L g605 ( .A(n_507), .B(n_589), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_507), .B(n_576), .Y(n_618) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_507), .Y(n_621) );
INVx1_ASAP7_75t_L g633 ( .A(n_507), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_507), .B(n_587), .Y(n_698) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_518), .B(n_527), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g562 ( .A(n_519), .B(n_546), .Y(n_562) );
AND2x4_ASAP7_75t_L g592 ( .A(n_519), .B(n_531), .Y(n_592) );
INVx2_ASAP7_75t_L g626 ( .A(n_519), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_519), .B(n_546), .Y(n_684) );
AND2x2_ASAP7_75t_L g731 ( .A(n_519), .B(n_560), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g719 ( .A1(n_527), .A2(n_591), .B1(n_634), .B2(n_694), .C1(n_720), .C2(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
AND2x2_ASAP7_75t_L g638 ( .A(n_529), .B(n_558), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_529), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g767 ( .A(n_529), .B(n_607), .Y(n_767) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_530), .A2(n_598), .B(n_602), .Y(n_597) );
AND2x2_ASAP7_75t_L g678 ( .A(n_530), .B(n_561), .Y(n_678) );
OR2x2_ASAP7_75t_L g703 ( .A(n_530), .B(n_562), .Y(n_703) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx5_ASAP7_75t_L g557 ( .A(n_531), .Y(n_557) );
AND2x2_ASAP7_75t_L g644 ( .A(n_531), .B(n_626), .Y(n_644) );
AND2x2_ASAP7_75t_L g670 ( .A(n_531), .B(n_546), .Y(n_670) );
OR2x2_ASAP7_75t_L g673 ( .A(n_531), .B(n_560), .Y(n_673) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_531), .Y(n_691) );
AND2x4_ASAP7_75t_SL g748 ( .A(n_531), .B(n_625), .Y(n_748) );
OR2x2_ASAP7_75t_L g757 ( .A(n_531), .B(n_584), .Y(n_757) );
OR2x6_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g590 ( .A(n_539), .Y(n_590) );
AOI221xp5_ASAP7_75t_SL g708 ( .A1(n_539), .A2(n_592), .B1(n_709), .B2(n_711), .C(n_712), .Y(n_708) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
OR2x2_ASAP7_75t_L g647 ( .A(n_540), .B(n_617), .Y(n_647) );
OR2x2_ASAP7_75t_L g657 ( .A(n_540), .B(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g683 ( .A(n_540), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g689 ( .A(n_540), .B(n_608), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_540), .B(n_672), .Y(n_701) );
INVx2_ASAP7_75t_L g714 ( .A(n_540), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_540), .B(n_592), .Y(n_735) );
AND2x2_ASAP7_75t_L g739 ( .A(n_540), .B(n_561), .Y(n_739) );
AND2x2_ASAP7_75t_L g747 ( .A(n_540), .B(n_748), .Y(n_747) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g560 ( .A(n_541), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_546), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g591 ( .A(n_546), .B(n_560), .Y(n_591) );
INVx2_ASAP7_75t_L g608 ( .A(n_546), .Y(n_608) );
AND2x4_ASAP7_75t_L g625 ( .A(n_546), .B(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_546), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g737 ( .A(n_556), .B(n_559), .Y(n_737) );
AND2x4_ASAP7_75t_L g583 ( .A(n_557), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g624 ( .A(n_557), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g651 ( .A(n_557), .B(n_591), .Y(n_651) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g755 ( .A(n_559), .B(n_756), .Y(n_755) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g607 ( .A(n_560), .B(n_608), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g627 ( .A1(n_561), .A2(n_628), .B(n_634), .Y(n_627) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_574), .Y(n_564) );
INVx1_ASAP7_75t_SL g681 ( .A(n_565), .Y(n_681) );
AND2x2_ASAP7_75t_L g711 ( .A(n_565), .B(n_621), .Y(n_711) );
AND2x4_ASAP7_75t_L g722 ( .A(n_565), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g588 ( .A(n_566), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g595 ( .A(n_566), .Y(n_595) );
AND2x4_ASAP7_75t_L g601 ( .A(n_566), .B(n_587), .Y(n_601) );
INVx2_ASAP7_75t_L g612 ( .A(n_566), .Y(n_612) );
INVx1_ASAP7_75t_L g661 ( .A(n_566), .Y(n_661) );
OR2x2_ASAP7_75t_L g682 ( .A(n_566), .B(n_666), .Y(n_682) );
OR2x2_ASAP7_75t_L g696 ( .A(n_566), .B(n_576), .Y(n_696) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_566), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_566), .B(n_618), .Y(n_768) );
OR2x6_ASAP7_75t_L g566 ( .A(n_567), .B(n_573), .Y(n_566) );
INVx1_ASAP7_75t_L g613 ( .A(n_574), .Y(n_613) );
AND2x2_ASAP7_75t_L g746 ( .A(n_574), .B(n_612), .Y(n_746) );
AND2x2_ASAP7_75t_L g771 ( .A(n_574), .B(n_601), .Y(n_771) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g589 ( .A(n_576), .Y(n_589) );
BUFx3_ASAP7_75t_L g631 ( .A(n_576), .Y(n_631) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_576), .Y(n_658) );
INVx1_ASAP7_75t_L g667 ( .A(n_576), .Y(n_667) );
AOI33xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .A3(n_590), .B1(n_591), .B2(n_592), .B3(n_593), .Y(n_582) );
AOI21x1_ASAP7_75t_SL g685 ( .A1(n_583), .A2(n_607), .B(n_669), .Y(n_685) );
INVx2_ASAP7_75t_L g715 ( .A(n_583), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_583), .B(n_714), .Y(n_721) );
AND2x2_ASAP7_75t_L g669 ( .A(n_584), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AND2x2_ASAP7_75t_L g632 ( .A(n_587), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g733 ( .A(n_588), .Y(n_733) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_589), .Y(n_723) );
OAI32xp33_ASAP7_75t_L g772 ( .A1(n_590), .A2(n_592), .A3(n_768), .B1(n_773), .B2(n_775), .Y(n_772) );
AND2x2_ASAP7_75t_L g690 ( .A(n_591), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g680 ( .A(n_592), .Y(n_680) );
AND2x2_ASAP7_75t_L g745 ( .A(n_592), .B(n_689), .Y(n_745) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_606), .B1(n_609), .B2(n_623), .C(n_627), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_600), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_601), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_601), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_601), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g650 ( .A(n_605), .Y(n_650) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_614), .C(n_619), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_611), .A2(n_673), .B1(n_713), .B2(n_716), .Y(n_712) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g616 ( .A(n_612), .Y(n_616) );
NOR2x1p5_ASAP7_75t_L g630 ( .A(n_612), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_612), .Y(n_652) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI322xp33_ASAP7_75t_L g679 ( .A1(n_615), .A2(n_657), .A3(n_680), .B1(n_681), .B2(n_682), .C1(n_683), .C2(n_685), .Y(n_679) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_617), .A2(n_636), .B(n_637), .C(n_639), .Y(n_635) );
OR2x2_ASAP7_75t_L g727 ( .A(n_617), .B(n_681), .Y(n_727) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g634 ( .A(n_618), .B(n_622), .Y(n_634) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g640 ( .A(n_624), .B(n_641), .Y(n_640) );
INVx3_ASAP7_75t_SL g672 ( .A(n_625), .Y(n_672) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_629), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_SL g676 ( .A(n_632), .Y(n_676) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_633), .Y(n_718) );
OR2x6_ASAP7_75t_SL g773 ( .A(n_636), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g763 ( .A1(n_641), .A2(n_764), .B(n_765), .C(n_772), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_645), .B(n_648), .C(n_652), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_643), .A2(n_655), .B(n_662), .C(n_686), .Y(n_654) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_699), .C(n_743), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_658), .Y(n_750) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g705 ( .A(n_661), .Y(n_705) );
NOR3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_675), .C(n_679), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_668), .B1(n_671), .B2(n_674), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g707 ( .A(n_667), .Y(n_707) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_667), .Y(n_774) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g760 ( .A(n_673), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OR2x2_ASAP7_75t_L g710 ( .A(n_676), .B(n_696), .Y(n_710) );
OR2x2_ASAP7_75t_L g761 ( .A(n_676), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g759 ( .A(n_684), .Y(n_759) );
OR2x2_ASAP7_75t_L g775 ( .A(n_684), .B(n_714), .Y(n_775) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .B(n_692), .Y(n_686) );
OAI31xp33_ASAP7_75t_L g700 ( .A1(n_687), .A2(n_701), .A3(n_702), .B(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g732 ( .A(n_697), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND4xp25_ASAP7_75t_SL g699 ( .A(n_700), .B(n_708), .C(n_719), .D(n_724), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_707), .Y(n_742) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B1(n_732), .B2(n_734), .C(n_736), .Y(n_724) );
NAND2xp33_ASAP7_75t_SL g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g769 ( .A(n_728), .Y(n_769) );
AND2x2_ASAP7_75t_SL g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI21xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g764 ( .A(n_738), .Y(n_764) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_744), .B(n_763), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_749), .C(n_753), .Y(n_744) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_758), .B(n_761), .Y(n_753) );
INVxp33_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_777), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
INVx3_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI22xp33_ASAP7_75t_SL g789 ( .A1(n_790), .A2(n_791), .B1(n_796), .B2(n_797), .Y(n_789) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND3x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .C(n_795), .Y(n_792) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
BUFx4f_ASAP7_75t_SL g811 ( .A(n_802), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g802 ( .A(n_803), .B(n_807), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
endmodule