module fake_jpeg_11108_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_37),
.B1(n_42),
.B2(n_33),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_25),
.B1(n_28),
.B2(n_18),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_43),
.B1(n_45),
.B2(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_22),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_20),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_41),
.B1(n_45),
.B2(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_102),
.B1(n_43),
.B2(n_40),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_103),
.B1(n_49),
.B2(n_22),
.Y(n_118)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_33),
.B1(n_37),
.B2(n_19),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_19),
.B(n_20),
.C(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_49),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_99),
.B1(n_42),
.B2(n_31),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_98),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_45),
.B1(n_39),
.B2(n_28),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_42),
.B1(n_36),
.B2(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_39),
.B1(n_32),
.B2(n_28),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_68),
.B1(n_54),
.B2(n_57),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_105),
.A2(n_107),
.B1(n_120),
.B2(n_130),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_57),
.B1(n_65),
.B2(n_40),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_115),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_39),
.B1(n_65),
.B2(n_31),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_121),
.B1(n_99),
.B2(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_111),
.B(n_117),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_32),
.B1(n_31),
.B2(n_26),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_32),
.B1(n_21),
.B2(n_26),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_90),
.C(n_79),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_27),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_17),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_17),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_26),
.B1(n_48),
.B2(n_36),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_76),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_145),
.B1(n_147),
.B2(n_158),
.Y(n_176)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_81),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_75),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_148),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_100),
.B1(n_93),
.B2(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_93),
.B1(n_100),
.B2(n_73),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_75),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_114),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_159),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_86),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_124),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_109),
.A2(n_100),
.B1(n_83),
.B2(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_125),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_100),
.B1(n_83),
.B2(n_32),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_113),
.B1(n_114),
.B2(n_98),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_125),
.B(n_119),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_49),
.B(n_29),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_115),
.B1(n_120),
.B2(n_107),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_164),
.B1(n_88),
.B2(n_77),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_100),
.B1(n_96),
.B2(n_77),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_138),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_137),
.B(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_167),
.A2(n_179),
.B(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_170),
.B(n_148),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_180),
.C(n_186),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_126),
.B(n_112),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_191),
.B(n_142),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_174),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_188),
.B1(n_198),
.B2(n_192),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_112),
.B(n_97),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_91),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_184),
.B1(n_136),
.B2(n_161),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_151),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_114),
.B1(n_97),
.B2(n_98),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_92),
.A3(n_91),
.B1(n_16),
.B2(n_13),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_158),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_48),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_26),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_36),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_22),
.B1(n_49),
.B2(n_92),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_164),
.B1(n_145),
.B2(n_152),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_189),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_13),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_171),
.A3(n_185),
.B1(n_35),
.B2(n_34),
.C1(n_29),
.C2(n_165),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_27),
.B1(n_35),
.B2(n_34),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_174),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_144),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_206),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_200),
.C(n_199),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_208),
.B1(n_216),
.B2(n_210),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_160),
.B(n_149),
.C(n_154),
.D(n_153),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_205),
.B(n_223),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_210),
.B(n_222),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_141),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_15),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_173),
.B1(n_188),
.B2(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_160),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_186),
.C(n_180),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_140),
.B(n_135),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_16),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_13),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_170),
.B(n_140),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_140),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_232),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_176),
.B(n_189),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_238),
.B1(n_215),
.B2(n_204),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_245),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_250),
.B1(n_203),
.B2(n_222),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_174),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_240),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_173),
.B1(n_189),
.B2(n_176),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_30),
.B1(n_17),
.B2(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_189),
.C(n_184),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_242),
.C(n_236),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_241),
.B(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_181),
.C(n_175),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_193),
.B(n_175),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_223),
.B(n_221),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_196),
.B1(n_34),
.B2(n_15),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_14),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_262),
.B1(n_234),
.B2(n_233),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_225),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_239),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_242),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_265),
.B1(n_266),
.B2(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_218),
.B1(n_221),
.B2(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_217),
.C(n_204),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_260),
.C(n_273),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_205),
.B1(n_226),
.B2(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_272),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_231),
.A2(n_14),
.B1(n_22),
.B2(n_30),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_230),
.B1(n_247),
.B2(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_243),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_270),
.B1(n_235),
.B2(n_266),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_248),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_275),
.B(n_289),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_234),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_290),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_282),
.C(n_288),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_232),
.C(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_279),
.C(n_280),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_291),
.B1(n_0),
.B2(n_3),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_244),
.B1(n_230),
.B2(n_247),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_255),
.B(n_273),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_252),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_0),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_251),
.A3(n_274),
.B1(n_265),
.B2(n_267),
.C1(n_263),
.C2(n_271),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_258),
.C(n_24),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_278),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_24),
.B(n_1),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_305),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

AOI211xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_290),
.B(n_286),
.C(n_277),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_30),
.C(n_3),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_30),
.C(n_4),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_8),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_315),
.B(n_295),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_4),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_316),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_5),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_314),
.A2(n_8),
.B(n_9),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_11),
.B(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_5),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_6),
.B(n_7),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_318),
.B(n_7),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_297),
.C(n_306),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_321),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_293),
.A3(n_305),
.B1(n_8),
.B2(n_9),
.C1(n_6),
.C2(n_11),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_315),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_310),
.B(n_314),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_10),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_312),
.C(n_9),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_322),
.B(n_326),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_334),
.A2(n_335),
.B(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_330),
.C(n_331),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_331),
.B(n_328),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_10),
.Y(n_340)
);


endmodule