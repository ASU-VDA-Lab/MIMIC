module fake_jpeg_15830_n_130 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g15 ( 
.A(n_0),
.B(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_45),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_2),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_2),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_3),
.B(n_4),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_6),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_27),
.B(n_7),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_61),
.B(n_63),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_76),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_62),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_30),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_75),
.Y(n_92)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_27),
.B1(n_23),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_43),
.B1(n_40),
.B2(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_24),
.B1(n_23),
.B2(n_39),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_83),
.B1(n_86),
.B2(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_14),
.B(n_89),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_63),
.B1(n_54),
.B2(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_43),
.B1(n_19),
.B2(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

XOR2x2_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_14),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_88),
.B(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_70),
.B1(n_58),
.B2(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_9),
.B1(n_12),
.B2(n_42),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_95),
.B(n_52),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_14),
.B1(n_60),
.B2(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_51),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_107),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_86),
.C(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_79),
.C(n_91),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_111),
.B(n_114),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_107),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_98),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_81),
.B(n_14),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_100),
.B1(n_106),
.B2(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_109),
.B1(n_108),
.B2(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_110),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_122),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_123),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g128 ( 
.A(n_126),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_82),
.A3(n_94),
.B1(n_96),
.B2(n_116),
.C(n_127),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_116),
.Y(n_130)
);


endmodule