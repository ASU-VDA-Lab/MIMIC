module fake_jpeg_23127_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_50),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_25),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_60),
.Y(n_103)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_59),
.B(n_86),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_21),
.C(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_36),
.B1(n_17),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_66),
.B1(n_68),
.B2(n_80),
.Y(n_105)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_17),
.B1(n_36),
.B2(n_27),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_17),
.B1(n_36),
.B2(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_84),
.B1(n_85),
.B2(n_19),
.Y(n_110)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_22),
.B1(n_18),
.B2(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_41),
.A2(n_18),
.B1(n_22),
.B2(n_33),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_24),
.B1(n_37),
.B2(n_31),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_91),
.Y(n_142)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_19),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_44),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_92),
.A2(n_47),
.B(n_34),
.Y(n_130)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_33),
.B1(n_66),
.B2(n_45),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_94),
.A2(n_102),
.B1(n_121),
.B2(n_10),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_100),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_99),
.B(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_33),
.B1(n_21),
.B2(n_30),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_111),
.B1(n_29),
.B2(n_28),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_109),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_24),
.B1(n_37),
.B2(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_0),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_29),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_47),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_1),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_54),
.A2(n_47),
.B1(n_34),
.B2(n_32),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_61),
.B1(n_77),
.B2(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_67),
.B(n_25),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_92),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_125),
.A2(n_130),
.B(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_75),
.B1(n_70),
.B2(n_28),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_129),
.B1(n_155),
.B2(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_127),
.B(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_137),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_148),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_32),
.B1(n_26),
.B2(n_0),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_143),
.B1(n_147),
.B2(n_97),
.Y(n_179)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_120),
.A3(n_115),
.B1(n_106),
.B2(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_146),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_26),
.B1(n_8),
.B2(n_2),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_0),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_1),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_88),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_156),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_107),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_104),
.C(n_117),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_171),
.C(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_166),
.B1(n_172),
.B2(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_159),
.B1(n_155),
.B2(n_128),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_157),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_167),
.A2(n_158),
.B1(n_137),
.B2(n_140),
.Y(n_203)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_189),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_107),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_119),
.B1(n_93),
.B2(n_100),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_173),
.B(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_117),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_144),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_125),
.A2(n_141),
.B1(n_127),
.B2(n_129),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_184),
.B1(n_188),
.B2(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_104),
.C(n_97),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_5),
.B(n_6),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_182),
.A2(n_163),
.B(n_177),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_124),
.B1(n_118),
.B2(n_10),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_124),
.B1(n_7),
.B2(n_10),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_186),
.A2(n_15),
.B1(n_16),
.B2(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_129),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_136),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_145),
.B1(n_149),
.B2(n_156),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_203),
.B1(n_215),
.B2(n_224),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_133),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_201),
.B(n_204),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_158),
.B(n_144),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_202),
.A2(n_207),
.B(n_213),
.C(n_190),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_205),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_138),
.B(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_209),
.Y(n_230)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_151),
.B(n_15),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_176),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_218),
.C(n_167),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_16),
.C(n_174),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_161),
.B(n_16),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_219),
.B(n_189),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_202),
.B1(n_201),
.B2(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_178),
.A2(n_165),
.B1(n_166),
.B2(n_192),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_190),
.B1(n_198),
.B2(n_202),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_171),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_215),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_186),
.B(n_195),
.C(n_170),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_238),
.C(n_224),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_167),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_236),
.A2(n_243),
.B(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_169),
.C(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_246),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_202),
.B1(n_196),
.B2(n_221),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_207),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_216),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_220),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_198),
.B1(n_202),
.B2(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_237),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_255),
.C(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_243),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_278),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_265),
.B(n_260),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_259),
.B1(n_228),
.B2(n_264),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_243),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.C(n_284),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_227),
.C(n_241),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_227),
.C(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_235),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_275),
.C(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_295),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_273),
.B1(n_271),
.B2(n_276),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_263),
.B1(n_246),
.B2(n_256),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_257),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_300),
.C(n_283),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_277),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_299),
.B1(n_269),
.B2(n_252),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_257),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_309),
.B1(n_232),
.B2(n_244),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_308),
.C(n_290),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_282),
.C(n_274),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_279),
.B1(n_250),
.B2(n_228),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_287),
.CI(n_244),
.CON(n_310),
.SN(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_297),
.Y(n_312)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_301),
.B(n_294),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_244),
.B(n_289),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.C(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_300),
.C(n_288),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_288),
.B(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_305),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_303),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_321),
.B(n_320),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_301),
.B(n_303),
.Y(n_329)
);

OAI311xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_313),
.A3(n_327),
.B1(n_309),
.C1(n_307),
.Y(n_330)
);

AOI221xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_240),
.B1(n_304),
.B2(n_213),
.C(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_274),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_323),
.Y(n_333)
);


endmodule