module fake_jpeg_16926_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_42),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_0),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_64),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_21),
.Y(n_70)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_29),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_70),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_94),
.B1(n_102),
.B2(n_18),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_33),
.B(n_30),
.C(n_28),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_77),
.A2(n_79),
.B(n_20),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_87),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_4),
.B(n_5),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_92),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_34),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_100),
.C(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_22),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_34),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_18),
.B1(n_38),
.B2(n_37),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_17),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_60),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_106),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_5),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_109),
.A2(n_110),
.B1(n_125),
.B2(n_6),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_85),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_20),
.Y(n_155)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_119),
.Y(n_145)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_124),
.Y(n_157)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_22),
.B1(n_35),
.B2(n_33),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_101),
.B1(n_104),
.B2(n_67),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_130),
.B1(n_103),
.B2(n_39),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_131),
.Y(n_159)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_39),
.B1(n_35),
.B2(n_30),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_138),
.Y(n_166)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_68),
.Y(n_151)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_88),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_77),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_149),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_85),
.B(n_81),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_155),
.B1(n_9),
.B2(n_10),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_69),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_165),
.C(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_92),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_163),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_156),
.C(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_66),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_153),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_74),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_170),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_79),
.B(n_7),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_96),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_6),
.B(n_7),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_96),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_99),
.C(n_80),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_86),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_90),
.C(n_80),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_109),
.B(n_86),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_9),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_13),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_185),
.C(n_200),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_126),
.B1(n_124),
.B2(n_141),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_132),
.B1(n_113),
.B2(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_187),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

XNOR2x2_ASAP7_75t_SL g192 ( 
.A(n_144),
.B(n_13),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_201),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_14),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_157),
.B(n_159),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_149),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_155),
.A2(n_146),
.B1(n_174),
.B2(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_178),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_152),
.A3(n_146),
.B1(n_162),
.B2(n_155),
.C1(n_168),
.C2(n_142),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_209),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_169),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_215),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_222),
.B(n_223),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_143),
.A3(n_150),
.B1(n_160),
.B2(n_163),
.C1(n_173),
.C2(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_217),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_175),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_175),
.C(n_196),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_185),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_206),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_186),
.B1(n_173),
.B2(n_196),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_213),
.B1(n_214),
.B2(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_220),
.C(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_188),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_184),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_235),
.B(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_248),
.Y(n_258)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_207),
.C(n_223),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_238),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_208),
.C(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_250),
.C(n_249),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_211),
.B(n_218),
.C(n_206),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_225),
.B(n_233),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_186),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_229),
.C(n_219),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_180),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_237),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_232),
.B1(n_234),
.B2(n_239),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_243),
.B1(n_247),
.B2(n_224),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_254),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_228),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_262),
.B(n_264),
.Y(n_270)
);

O2A1O1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_259),
.B(n_247),
.C(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_255),
.C(n_253),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_266),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_259),
.B1(n_262),
.B2(n_247),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.C(n_270),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);


endmodule