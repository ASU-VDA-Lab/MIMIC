module fake_ariane_880_n_1694 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1694);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1694;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_94),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_60),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_35),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_80),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_48),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_48),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_51),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_57),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_109),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_46),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_69),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_85),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_65),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_53),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_56),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_53),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_79),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_36),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_106),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_46),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_100),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_90),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_91),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_30),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_5),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_23),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_35),
.Y(n_197)
);

INVxp33_ASAP7_75t_SL g198 ( 
.A(n_83),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_34),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_21),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_132),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_113),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_101),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_52),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_64),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_49),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_42),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_67),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_81),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_68),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_43),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_107),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_62),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_16),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_37),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_59),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_33),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_89),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_117),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_128),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_110),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_5),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_24),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_142),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_8),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_70),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_134),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_114),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_49),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_20),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_26),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_137),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_125),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_72),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_26),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_15),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_50),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_119),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_123),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_50),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_4),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_22),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_0),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_118),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_2),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_96),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_146),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_103),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_12),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_20),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_55),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_127),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_43),
.Y(n_276)
);

CKINVDCx11_ASAP7_75t_R g277 ( 
.A(n_121),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_115),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_17),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_108),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_40),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_61),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_148),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_54),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_33),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_124),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_27),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_13),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_38),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_55),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_111),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_14),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_66),
.Y(n_295)
);

INVxp33_ASAP7_75t_R g296 ( 
.A(n_47),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_1),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_R g299 ( 
.A(n_150),
.B(n_97),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_290),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_282),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_154),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_183),
.B(n_2),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_193),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_202),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_3),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_191),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_244),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_188),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_159),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_252),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_257),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_3),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_158),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_283),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_4),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_152),
.B(n_6),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_194),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_194),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_194),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_194),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_188),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_194),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_169),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_195),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_276),
.B(n_7),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_199),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_179),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_206),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_8),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_164),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_216),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_161),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_166),
.B(n_9),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_239),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_164),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_223),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_223),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_245),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_158),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_245),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_157),
.Y(n_356)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_169),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_186),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_171),
.B(n_9),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_157),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_163),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_265),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_196),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_197),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_214),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_214),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_224),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_201),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_180),
.Y(n_369)
);

BUFx2_ASAP7_75t_SL g370 ( 
.A(n_158),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_182),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_326),
.B(n_354),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_234),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_316),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_234),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_175),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_307),
.Y(n_382)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_205),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_205),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_370),
.A2(n_271),
.B1(n_274),
.B2(n_296),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_312),
.B(n_234),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

AND2x6_ASAP7_75t_L g397 ( 
.A(n_329),
.B(n_231),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_R g400 ( 
.A(n_338),
.B(n_357),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_326),
.B(n_354),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_334),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_178),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_287),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_330),
.B(n_198),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_337),
.Y(n_412)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_360),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_366),
.B(n_181),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_336),
.B(n_243),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_367),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_207),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_311),
.B(n_198),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_370),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_350),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_306),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_359),
.B(n_224),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_313),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_303),
.Y(n_433)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_308),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_287),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_380),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_376),
.B(n_250),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_250),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_372),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_342),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_426),
.B(n_358),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_440),
.A2(n_304),
.B1(n_298),
.B2(n_348),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_377),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_364),
.C(n_363),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_426),
.B(n_368),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_377),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_324),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_321),
.C(n_298),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_377),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_430),
.B1(n_411),
.B2(n_413),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_318),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_440),
.A2(n_430),
.B1(n_411),
.B2(n_413),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_301),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_373),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_347),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_376),
.B(n_327),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_376),
.B(n_150),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_438),
.B(n_323),
.Y(n_476)
);

INVx4_ASAP7_75t_SL g477 ( 
.A(n_397),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_429),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_382),
.B(n_300),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_397),
.B(n_156),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

AND2x2_ASAP7_75t_SL g484 ( 
.A(n_378),
.B(n_328),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_374),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_416),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_416),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_438),
.B(n_340),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_438),
.B(n_361),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_228),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_390),
.A2(n_420),
.B1(n_378),
.B2(n_400),
.Y(n_498)
);

AO22x2_ASAP7_75t_L g499 ( 
.A1(n_378),
.A2(n_225),
.B1(n_286),
.B2(n_261),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_418),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_418),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_378),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_390),
.B(n_151),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_373),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_439),
.B(n_369),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_373),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_379),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_433),
.B(n_302),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_439),
.B(n_258),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_439),
.B(n_309),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_400),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_399),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_413),
.A2(n_344),
.B1(n_260),
.B2(n_288),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_390),
.B(n_151),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_387),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_380),
.Y(n_531)
);

BUFx4f_ASAP7_75t_L g532 ( 
.A(n_397),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_413),
.A2(n_344),
.B1(n_291),
.B2(n_200),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_403),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_406),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_384),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_413),
.B(n_310),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_433),
.B(n_314),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_406),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_379),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_397),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_413),
.B(n_315),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_387),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_390),
.B(n_153),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_408),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_431),
.B(n_173),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_408),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

BUFx8_ASAP7_75t_SL g551 ( 
.A(n_433),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_380),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_408),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_388),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_379),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_420),
.B(n_213),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_395),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_420),
.B(n_230),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_420),
.Y(n_561)
);

AO22x1_ASAP7_75t_L g562 ( 
.A1(n_397),
.A2(n_254),
.B1(n_256),
.B2(n_262),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_408),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_395),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_434),
.B(n_212),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_431),
.B(n_173),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_380),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_395),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_414),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_412),
.Y(n_570)
);

CKINVDCx6p67_ASAP7_75t_R g571 ( 
.A(n_375),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_384),
.B(n_153),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_414),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_384),
.B(n_155),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_434),
.B(n_375),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_434),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_412),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_414),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_412),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_425),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_412),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_412),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_414),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_434),
.B(n_215),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_434),
.A2(n_247),
.B1(n_255),
.B2(n_294),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_434),
.B(n_219),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_532),
.B(n_380),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_451),
.A2(n_434),
.B1(n_253),
.B2(n_241),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_485),
.B(n_405),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_561),
.B(n_405),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_561),
.B(n_384),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_485),
.B(n_388),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_496),
.B(n_384),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_509),
.B(n_384),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_532),
.B(n_387),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_443),
.B(n_385),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_469),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_499),
.A2(n_397),
.B1(n_410),
.B2(n_415),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_468),
.B(n_388),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_443),
.B(n_385),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_523),
.B(n_299),
.C(n_381),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_508),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_532),
.B(n_387),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_484),
.A2(n_465),
.B1(n_462),
.B2(n_459),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_484),
.B(n_482),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_443),
.B(n_385),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_498),
.B(n_385),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_505),
.A2(n_449),
.B1(n_460),
.B2(n_527),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_468),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_511),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_472),
.B(n_385),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_443),
.B(n_385),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_442),
.B(n_387),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_513),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_452),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_441),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_514),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_443),
.B(n_410),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_443),
.B(n_446),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_446),
.B(n_410),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_576),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_446),
.B(n_410),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_514),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_472),
.B(n_477),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_499),
.A2(n_397),
.B1(n_410),
.B2(n_415),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_542),
.A2(n_381),
.B(n_391),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_529),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_452),
.Y(n_633)
);

AOI221xp5_ASAP7_75t_L g634 ( 
.A1(n_472),
.A2(n_262),
.B1(n_237),
.B2(n_241),
.C(n_246),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_542),
.A2(n_436),
.B(n_425),
.C(n_432),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_446),
.A2(n_397),
.B1(n_410),
.B2(n_172),
.Y(n_636)
);

NAND3x1_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_341),
.C(n_339),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_505),
.B(n_391),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_478),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_529),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_446),
.B(n_397),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_471),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_517),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_446),
.A2(n_397),
.B1(n_172),
.B2(n_168),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_442),
.B(n_391),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_442),
.B(n_391),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_520),
.B(n_391),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_575),
.B(n_391),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_535),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_507),
.A2(n_546),
.B1(n_475),
.B2(n_556),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_522),
.B(n_391),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_536),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_464),
.B(n_391),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_478),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_523),
.B(n_454),
.C(n_544),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_536),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_476),
.B(n_432),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_467),
.B(n_391),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_497),
.B(n_521),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_478),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_495),
.B(n_432),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_436),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_558),
.A2(n_165),
.B1(n_273),
.B2(n_162),
.Y(n_666)
);

AO221x1_ASAP7_75t_L g667 ( 
.A1(n_499),
.A2(n_292),
.B1(n_238),
.B2(n_249),
.C(n_156),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_520),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_479),
.B(n_409),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_483),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_520),
.B(n_392),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_450),
.B(n_392),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_464),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_558),
.B(n_436),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_540),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_565),
.B(n_415),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_488),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_488),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_455),
.B(n_392),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_491),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_584),
.B(n_415),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_531),
.B(n_392),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_541),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_474),
.B(n_392),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_586),
.B(n_419),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_479),
.B(n_419),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_531),
.B(n_552),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_531),
.B(n_392),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_548),
.A2(n_422),
.B1(n_256),
.B2(n_253),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_541),
.Y(n_690)
);

INVx8_ASAP7_75t_L g691 ( 
.A(n_457),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_555),
.A2(n_422),
.B(n_428),
.C(n_427),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_552),
.B(n_424),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_552),
.B(n_392),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_567),
.B(n_424),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_567),
.B(n_424),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_491),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_572),
.A2(n_177),
.B1(n_176),
.B2(n_174),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_557),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_477),
.B(n_424),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_567),
.B(n_427),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_557),
.B(n_427),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_463),
.B(n_254),
.C(n_264),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_564),
.B(n_427),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_492),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_564),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_492),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_574),
.B(n_392),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_506),
.Y(n_710)
);

AOI221xp5_ASAP7_75t_L g711 ( 
.A1(n_499),
.A2(n_264),
.B1(n_275),
.B2(n_227),
.C(n_220),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_537),
.B(n_392),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_568),
.A2(n_412),
.B(n_435),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_537),
.A2(n_162),
.B1(n_177),
.B2(n_176),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_477),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_571),
.B(n_394),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_568),
.B(n_428),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_516),
.B(n_343),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_453),
.A2(n_275),
.B1(n_204),
.B2(n_210),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_482),
.A2(n_435),
.B1(n_428),
.B2(n_417),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_510),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_394),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_512),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_512),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_490),
.B(n_394),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_SL g727 ( 
.A1(n_493),
.A2(n_435),
.B(n_428),
.C(n_401),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_500),
.B(n_435),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_524),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_501),
.B(n_394),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_548),
.B(n_346),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_444),
.A2(n_447),
.B(n_445),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_477),
.B(n_383),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_383),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_515),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_518),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_519),
.B(n_394),
.Y(n_737)
);

AOI22x1_ASAP7_75t_L g738 ( 
.A1(n_524),
.A2(n_394),
.B1(n_396),
.B2(n_404),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_559),
.B(n_394),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_560),
.A2(n_417),
.B1(n_437),
.B2(n_243),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_580),
.B(n_526),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_457),
.B(n_494),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_534),
.B(n_396),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_569),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_457),
.B(n_396),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_457),
.B(n_383),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_569),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_445),
.B(n_396),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_457),
.B(n_396),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_494),
.B(n_396),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_573),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_588),
.A2(n_448),
.B(n_447),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_661),
.B(n_566),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_675),
.B(n_562),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_719),
.Y(n_755)
);

AOI21x1_ASAP7_75t_L g756 ( 
.A1(n_596),
.A2(n_456),
.B(n_448),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_607),
.A2(n_486),
.B1(n_481),
.B2(n_504),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_621),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_607),
.A2(n_486),
.B1(n_481),
.B2(n_504),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_606),
.A2(n_487),
.B(n_480),
.C(n_470),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_588),
.A2(n_461),
.B(n_456),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_687),
.A2(n_685),
.B(n_695),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_591),
.B(n_516),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_695),
.A2(n_466),
.B(n_461),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_694),
.A2(n_470),
.B(n_466),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_628),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_609),
.B(n_566),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_609),
.B(n_562),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_696),
.A2(n_487),
.B(n_480),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_598),
.A2(n_549),
.B1(n_582),
.B2(n_581),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_689),
.B(n_612),
.C(n_611),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_591),
.B(n_573),
.Y(n_772)
);

INVx11_ASAP7_75t_L g773 ( 
.A(n_629),
.Y(n_773)
);

OAI21xp33_ASAP7_75t_L g774 ( 
.A1(n_666),
.A2(n_211),
.B(n_203),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_697),
.A2(n_525),
.B(n_582),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_623),
.B(n_673),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_620),
.Y(n_777)
);

AO21x1_ASAP7_75t_L g778 ( 
.A1(n_649),
.A2(n_583),
.B(n_578),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_632),
.A2(n_583),
.B(n_578),
.C(n_579),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_702),
.A2(n_581),
.B(n_579),
.Y(n_780)
);

OAI21xp33_ASAP7_75t_L g781 ( 
.A1(n_634),
.A2(n_229),
.B(n_285),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_525),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_640),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_665),
.B(n_530),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_645),
.A2(n_577),
.B(n_570),
.C(n_563),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_673),
.B(n_464),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_674),
.B(n_530),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_614),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_649),
.A2(n_577),
.B(n_570),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_650),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_614),
.B(n_533),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_653),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_730),
.A2(n_563),
.B(n_553),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_656),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_737),
.A2(n_739),
.B(n_663),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_658),
.A2(n_553),
.B(n_550),
.C(n_549),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_731),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_669),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_748),
.A2(n_533),
.B(n_550),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_617),
.A2(n_538),
.B(n_547),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_617),
.A2(n_538),
.B(n_547),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_646),
.A2(n_502),
.B(n_545),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_604),
.A2(n_473),
.B1(n_545),
.B2(n_464),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_646),
.A2(n_502),
.B(n_545),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_647),
.A2(n_502),
.B(n_545),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_600),
.B(n_349),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_659),
.B(n_473),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_631),
.A2(n_543),
.B(n_494),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_594),
.B(n_473),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_595),
.B(n_473),
.Y(n_810)
);

OAI21xp33_ASAP7_75t_L g811 ( 
.A1(n_589),
.A2(n_217),
.B(n_280),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_673),
.B(n_473),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_656),
.B(n_494),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_624),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_683),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_669),
.B(n_554),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_660),
.B(n_489),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_673),
.B(n_489),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_647),
.A2(n_545),
.B(n_528),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_657),
.B(n_554),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_648),
.A2(n_502),
.B(n_528),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_648),
.A2(n_502),
.B(n_528),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_624),
.B(n_489),
.Y(n_823)
);

CKINVDCx14_ASAP7_75t_R g824 ( 
.A(n_593),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_660),
.B(n_489),
.Y(n_825)
);

NAND2x1p5_ASAP7_75t_L g826 ( 
.A(n_716),
.B(n_494),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_652),
.B(n_489),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_671),
.A2(n_528),
.B(n_543),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_671),
.A2(n_528),
.B(n_543),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_599),
.A2(n_437),
.B1(n_417),
.B2(n_362),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_652),
.A2(n_222),
.B(n_281),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_682),
.A2(n_543),
.B(n_396),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_732),
.A2(n_543),
.B(n_401),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_669),
.B(n_437),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_686),
.B(n_735),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_682),
.A2(n_396),
.B(n_503),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_686),
.B(n_736),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_688),
.A2(n_396),
.B(n_503),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_633),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_686),
.B(n_437),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_596),
.A2(n_401),
.B(n_404),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_716),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_639),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_643),
.B(n_437),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_633),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_592),
.B(n_437),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_662),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_688),
.A2(n_458),
.B(n_503),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_626),
.B(n_417),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_651),
.B(n_437),
.Y(n_850)
);

INVx11_ASAP7_75t_L g851 ( 
.A(n_629),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_613),
.B(n_437),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_626),
.B(n_417),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_690),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_692),
.A2(n_437),
.B(n_233),
.C(n_295),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_605),
.A2(n_458),
.B(n_167),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_701),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_714),
.A2(n_404),
.B(n_401),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_618),
.B(n_417),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_700),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_629),
.Y(n_861)
);

OAI21xp33_ASAP7_75t_L g862 ( 
.A1(n_689),
.A2(n_218),
.B(n_232),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_707),
.B(n_417),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_587),
.B(n_601),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_590),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_610),
.B(n_417),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_629),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_616),
.B(n_417),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_655),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_605),
.A2(n_458),
.B(n_160),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_703),
.A2(n_718),
.B(n_705),
.Y(n_871)
);

AOI33xp33_ASAP7_75t_L g872 ( 
.A1(n_711),
.A2(n_699),
.A3(n_747),
.B1(n_744),
.B2(n_751),
.B3(n_630),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_629),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_726),
.A2(n_404),
.B(n_263),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_668),
.B(n_717),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_622),
.B(n_383),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_625),
.B(n_383),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_684),
.A2(n_160),
.B1(n_155),
.B2(n_165),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_635),
.A2(n_293),
.B(n_268),
.C(n_251),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_655),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_720),
.A2(n_289),
.B(n_551),
.C(n_14),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_717),
.B(n_383),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_723),
.B(n_383),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_684),
.B(n_551),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_672),
.A2(n_273),
.B(n_170),
.C(n_242),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_722),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_240),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_672),
.B(n_240),
.Y(n_888)
);

CKINVDCx6p67_ASAP7_75t_R g889 ( 
.A(n_627),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_724),
.Y(n_890)
);

NAND3x1_ASAP7_75t_L g891 ( 
.A(n_704),
.B(n_284),
.C(n_267),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_726),
.A2(n_242),
.B(n_149),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_679),
.B(n_243),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_679),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_701),
.B(n_407),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_676),
.A2(n_235),
.B(n_190),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_638),
.A2(n_407),
.B1(n_402),
.B2(n_398),
.Y(n_897)
);

AOI33xp33_ASAP7_75t_L g898 ( 
.A1(n_599),
.A2(n_10),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.B3(n_17),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_681),
.A2(n_236),
.B(n_192),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_654),
.A2(n_185),
.B(n_208),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_713),
.A2(n_278),
.B(n_221),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_284),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_638),
.A2(n_407),
.B1(n_402),
.B2(n_398),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_637),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_713),
.A2(n_184),
.B(n_226),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_715),
.B(n_267),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_597),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_630),
.B(n_267),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_602),
.B(n_284),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_740),
.B(n_10),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_725),
.B(n_187),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_729),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_733),
.B(n_407),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_728),
.A2(n_189),
.B(n_209),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_727),
.A2(n_407),
.B(n_402),
.C(n_398),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_709),
.A2(n_407),
.B(n_402),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_709),
.A2(n_402),
.B(n_398),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_727),
.A2(n_402),
.B(n_398),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_693),
.A2(n_407),
.B(n_402),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_664),
.Y(n_920)
);

AOI21xp33_ASAP7_75t_L g921 ( 
.A1(n_608),
.A2(n_407),
.B(n_402),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_670),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_678),
.B(n_19),
.Y(n_923)
);

CKINVDCx8_ASAP7_75t_R g924 ( 
.A(n_734),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_636),
.B(n_398),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_615),
.A2(n_398),
.B1(n_249),
.B2(n_238),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_691),
.A2(n_398),
.B(n_249),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_678),
.B(n_19),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_710),
.B(n_23),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_644),
.A2(n_398),
.B1(n_249),
.B2(n_238),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_817),
.A2(n_691),
.B(n_641),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_841),
.A2(n_738),
.B(n_712),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_773),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_825),
.A2(n_691),
.B(n_749),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_777),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_763),
.B(n_710),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_830),
.A2(n_734),
.B1(n_667),
.B2(n_642),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_758),
.Y(n_938)
);

AO32x1_ASAP7_75t_L g939 ( 
.A1(n_910),
.A2(n_712),
.A3(n_619),
.B1(n_677),
.B2(n_680),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_763),
.B(n_698),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_867),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_753),
.B(n_740),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_760),
.A2(n_706),
.B(n_708),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_767),
.A2(n_721),
.B1(n_743),
.B2(n_745),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_797),
.B(n_750),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_830),
.A2(n_721),
.B1(n_750),
.B2(n_745),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_867),
.B(n_733),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_766),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_847),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_794),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_SL g951 ( 
.A(n_867),
.B(n_746),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_749),
.B(n_742),
.C(n_746),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_768),
.A2(n_156),
.B1(n_238),
.B2(n_249),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_783),
.A2(n_156),
.B1(n_238),
.B2(n_28),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_843),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_754),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_906),
.A2(n_742),
.B(n_25),
.C(n_28),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_SL g958 ( 
.A(n_867),
.B(n_156),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_790),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_873),
.B(n_84),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_845),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_788),
.B(n_31),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_816),
.B(n_31),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_906),
.B(n_32),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_827),
.A2(n_86),
.B(n_147),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_884),
.B(n_32),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_884),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_788),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_762),
.A2(n_92),
.B(n_145),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_851),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_871),
.A2(n_88),
.B(n_133),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_807),
.A2(n_82),
.B(n_122),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_L g973 ( 
.A1(n_862),
.A2(n_44),
.B(n_45),
.Y(n_973)
);

BUFx4f_ASAP7_75t_L g974 ( 
.A(n_754),
.Y(n_974)
);

INVx6_ASAP7_75t_L g975 ( 
.A(n_755),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_861),
.B(n_44),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_904),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_809),
.A2(n_95),
.B(n_116),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_SL g979 ( 
.A1(n_806),
.A2(n_45),
.B1(n_47),
.B2(n_51),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_869),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_792),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_895),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_824),
.A2(n_820),
.B1(n_893),
.B2(n_781),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_888),
.A2(n_98),
.B(n_99),
.C(n_112),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_857),
.B(n_889),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_SL g987 ( 
.A(n_881),
.B(n_774),
.C(n_811),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_857),
.B(n_798),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_813),
.B(n_894),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_SL g990 ( 
.A1(n_823),
.A2(n_779),
.B(n_785),
.C(n_796),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_810),
.A2(n_875),
.B(n_795),
.Y(n_991)
);

INVx3_ASAP7_75t_SL g992 ( 
.A(n_754),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_893),
.A2(n_888),
.B1(n_909),
.B2(n_835),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_918),
.A2(n_756),
.B(n_915),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_SL g995 ( 
.A(n_885),
.B(n_837),
.C(n_854),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_SL g996 ( 
.A(n_924),
.B(n_861),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_815),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_860),
.A2(n_772),
.B1(n_784),
.B2(n_787),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_879),
.A2(n_782),
.B(n_872),
.C(n_909),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_920),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_885),
.A2(n_760),
.B(n_791),
.C(n_759),
.Y(n_1001)
);

AOI22x1_ASAP7_75t_L g1002 ( 
.A1(n_775),
.A2(n_780),
.B1(n_765),
.B2(n_769),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_842),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_813),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_757),
.A2(n_864),
.B(n_779),
.C(n_796),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_907),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_865),
.B(n_907),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_834),
.B(n_840),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_778),
.A2(n_831),
.B(n_919),
.C(n_823),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_785),
.A2(n_855),
.B(n_770),
.C(n_887),
.Y(n_1010)
);

AND2x2_ASAP7_75t_SL g1011 ( 
.A(n_898),
.B(n_908),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_898),
.B(n_878),
.C(n_855),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_764),
.A2(n_799),
.B(n_793),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_782),
.A2(n_850),
.B(n_902),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_890),
.A2(n_912),
.B1(n_844),
.B2(n_922),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_803),
.A2(n_786),
.B(n_818),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_895),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_913),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_786),
.A2(n_818),
.B(n_812),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_913),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_842),
.B(n_849),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_814),
.B(n_911),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_891),
.B(n_892),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_874),
.A2(n_929),
.B(n_928),
.C(n_923),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_852),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_859),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_826),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_846),
.B(n_789),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_812),
.A2(n_916),
.B(n_752),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_761),
.A2(n_804),
.B(n_819),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_849),
.A2(n_853),
.B(n_863),
.C(n_868),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_776),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_866),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_853),
.B(n_901),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_826),
.Y(n_1036)
);

CKINVDCx8_ASAP7_75t_R g1037 ( 
.A(n_905),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_930),
.A2(n_800),
.B(n_801),
.C(n_896),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_802),
.A2(n_805),
.B(n_821),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_899),
.A2(n_914),
.B(n_858),
.C(n_897),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_876),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_925),
.A2(n_917),
.B(n_882),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_822),
.A2(n_848),
.B(n_828),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_876),
.B(n_877),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_900),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_L g1046 ( 
.A(n_903),
.B(n_877),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_925),
.A2(n_856),
.B1(n_870),
.B2(n_838),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_921),
.B(n_836),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_927),
.B(n_832),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_829),
.A2(n_883),
.B(n_808),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_833),
.A2(n_825),
.B(n_817),
.Y(n_1051)
);

INVx5_ASAP7_75t_L g1052 ( 
.A(n_867),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_906),
.A2(n_888),
.B(n_763),
.C(n_767),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_839),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_767),
.A2(n_607),
.B1(n_606),
.B2(n_753),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_767),
.A2(n_607),
.B1(n_606),
.B2(n_753),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_763),
.B(n_523),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_763),
.B(n_426),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_867),
.B(n_794),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_SL g1060 ( 
.A1(n_919),
.A2(n_423),
.B(n_638),
.C(n_726),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_847),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_839),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_763),
.B(n_426),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_964),
.B(n_1057),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_998),
.A2(n_1051),
.B(n_1029),
.Y(n_1066)
);

AOI221x1_ASAP7_75t_L g1067 ( 
.A1(n_973),
.A2(n_954),
.B1(n_1012),
.B2(n_999),
.C(n_1014),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1050),
.A2(n_1025),
.B(n_1039),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_935),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1055),
.A2(n_1056),
.B1(n_993),
.B2(n_1011),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_963),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1009),
.A2(n_1056),
.B(n_1055),
.Y(n_1073)
);

AOI211x1_ASAP7_75t_L g1074 ( 
.A1(n_959),
.A2(n_954),
.B(n_966),
.C(n_962),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_968),
.B(n_979),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1013),
.A2(n_1031),
.B(n_1002),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1000),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1058),
.B(n_1063),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_945),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1017),
.A2(n_1046),
.B(n_1045),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1030),
.A2(n_1005),
.B(n_1048),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_953),
.A2(n_1047),
.A3(n_1038),
.B(n_944),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_938),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_948),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1001),
.A2(n_1010),
.B(n_1032),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_1036),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1006),
.B(n_940),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_957),
.A2(n_987),
.B(n_995),
.C(n_936),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_992),
.A2(n_967),
.B1(n_956),
.B2(n_1007),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1042),
.A2(n_1049),
.B(n_1020),
.Y(n_1090)
);

BUFx5_ASAP7_75t_L g1091 ( 
.A(n_1034),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1047),
.A2(n_943),
.B(n_931),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1023),
.A2(n_942),
.B(n_952),
.C(n_984),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_997),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_949),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_943),
.A2(n_969),
.B(n_971),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1040),
.A2(n_934),
.B(n_965),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_982),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_933),
.B(n_1004),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_SL g1101 ( 
.A1(n_1024),
.A2(n_1041),
.B(n_1033),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_974),
.A2(n_1018),
.B1(n_1054),
.B2(n_980),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1008),
.B(n_988),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_989),
.B(n_988),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_941),
.B(n_1052),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1059),
.B(n_996),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1059),
.B(n_996),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_990),
.A2(n_1060),
.B(n_958),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_985),
.A2(n_946),
.B(n_974),
.C(n_1026),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_972),
.A2(n_978),
.B(n_1035),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_975),
.B(n_950),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1022),
.A2(n_960),
.B(n_1016),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_949),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_961),
.A2(n_983),
.A3(n_1062),
.B(n_939),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_958),
.A2(n_1028),
.B(n_981),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1027),
.A2(n_981),
.B(n_1028),
.C(n_959),
.Y(n_1116)
);

CKINVDCx8_ASAP7_75t_R g1117 ( 
.A(n_941),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_977),
.B(n_1015),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_SL g1119 ( 
.A1(n_976),
.A2(n_960),
.B(n_947),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_941),
.B(n_1052),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_976),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_975),
.B(n_986),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_937),
.A2(n_947),
.B(n_1021),
.C(n_970),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1052),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_1061),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_939),
.A2(n_1044),
.A3(n_1037),
.B(n_1022),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_976),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_970),
.B(n_933),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1019),
.B(n_1003),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1019),
.B(n_1044),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1052),
.A2(n_1019),
.B(n_951),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_951),
.A2(n_1042),
.B(n_1043),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1057),
.B(n_753),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_935),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1057),
.B(n_753),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1000),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1000),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_935),
.B(n_468),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1025),
.A2(n_778),
.A3(n_953),
.B(n_831),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1057),
.B(n_753),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_935),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1057),
.B(n_753),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_949),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_935),
.B(n_468),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_964),
.B(n_523),
.C(n_540),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_938),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_938),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_1006),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_938),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_964),
.B(n_523),
.Y(n_1162)
);

CKINVDCx11_ASAP7_75t_R g1163 ( 
.A(n_955),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1165)
);

INVx3_ASAP7_75t_SL g1166 ( 
.A(n_975),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_964),
.B(n_523),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1025),
.A2(n_778),
.A3(n_953),
.B(n_831),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_935),
.B(n_612),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_964),
.A2(n_906),
.B1(n_992),
.B2(n_967),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_994),
.A2(n_932),
.B(n_1043),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1025),
.A2(n_778),
.A3(n_953),
.B(n_831),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_964),
.A2(n_1053),
.B(n_993),
.C(n_906),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1025),
.A2(n_778),
.A3(n_953),
.B(n_831),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_935),
.B(n_468),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_1004),
.B(n_941),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1053),
.A2(n_964),
.B1(n_767),
.B2(n_993),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_1053),
.A2(n_999),
.B(n_1060),
.C(n_964),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_933),
.B(n_1004),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_933),
.B(n_1004),
.Y(n_1182)
);

BUFx4_ASAP7_75t_SL g1183 ( 
.A(n_976),
.Y(n_1183)
);

AOI221x1_ASAP7_75t_L g1184 ( 
.A1(n_964),
.A2(n_1053),
.B1(n_973),
.B2(n_954),
.C(n_1012),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_935),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_964),
.A2(n_771),
.B1(n_767),
.B2(n_1053),
.Y(n_1186)
);

NOR2xp67_ASAP7_75t_SL g1187 ( 
.A(n_955),
.B(n_426),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1057),
.B(n_753),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_935),
.B(n_612),
.Y(n_1189)
);

AO21x1_ASAP7_75t_L g1190 ( 
.A1(n_993),
.A2(n_964),
.B(n_998),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1025),
.A2(n_778),
.A3(n_953),
.B(n_831),
.Y(n_1191)
);

AO32x2_ASAP7_75t_L g1192 ( 
.A1(n_1055),
.A2(n_1056),
.A3(n_998),
.B1(n_954),
.B2(n_953),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_964),
.A2(n_689),
.B1(n_451),
.B2(n_304),
.C(n_460),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_991),
.A2(n_998),
.B(n_1053),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1117),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1083),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1190),
.B(n_1178),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1166),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1065),
.A2(n_1195),
.B1(n_1162),
.B2(n_1167),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1105),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1146),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1084),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1077),
.Y(n_1205)
);

INVx3_ASAP7_75t_SL g1206 ( 
.A(n_1113),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1096),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1178),
.A2(n_1075),
.B1(n_1154),
.B2(n_1164),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1186),
.B(n_1071),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1153),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1171),
.A2(n_1186),
.B1(n_1156),
.B2(n_1071),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1139),
.B(n_1155),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1086),
.Y(n_1213)
);

CKINVDCx6p67_ASAP7_75t_R g1214 ( 
.A(n_1163),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1137),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1174),
.A2(n_1154),
.B1(n_1164),
.B2(n_1188),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1073),
.A2(n_1133),
.B1(n_1152),
.B2(n_1142),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1089),
.A2(n_1136),
.B1(n_1102),
.B2(n_1099),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1094),
.B(n_1087),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1088),
.A2(n_1074),
.B1(n_1116),
.B2(n_1073),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1138),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1095),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1157),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1158),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1170),
.Y(n_1225)
);

CKINVDCx11_ASAP7_75t_R g1226 ( 
.A(n_1141),
.Y(n_1226)
);

CKINVDCx6p67_ASAP7_75t_R g1227 ( 
.A(n_1125),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1092),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1072),
.A2(n_1176),
.B1(n_1078),
.B2(n_1127),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1086),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1189),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1069),
.A2(n_1135),
.B1(n_1185),
.B2(n_1103),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1161),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1069),
.A2(n_1135),
.B1(n_1185),
.B2(n_1159),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1092),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1184),
.A2(n_1064),
.B(n_1194),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1121),
.A2(n_1079),
.B1(n_1104),
.B2(n_1187),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1147),
.B(n_1148),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1183),
.A2(n_1085),
.B1(n_1115),
.B2(n_1165),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1111),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1100),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_1118),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1122),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1106),
.Y(n_1244)
);

BUFx8_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1114),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1085),
.A2(n_1091),
.B1(n_1107),
.B2(n_1193),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1181),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1067),
.A2(n_1196),
.B1(n_1179),
.B2(n_1169),
.Y(n_1249)
);

INVx6_ASAP7_75t_L g1250 ( 
.A(n_1181),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1128),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1114),
.Y(n_1252)
);

BUFx10_ASAP7_75t_L g1253 ( 
.A(n_1182),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1182),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1130),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1129),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1151),
.A2(n_1192),
.B1(n_1080),
.B2(n_1074),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1192),
.A2(n_1112),
.B1(n_1097),
.B2(n_1091),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1101),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1091),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1109),
.A2(n_1066),
.B1(n_1123),
.B2(n_1119),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1091),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1091),
.Y(n_1263)
);

NAND2x1p5_ASAP7_75t_L g1264 ( 
.A(n_1131),
.B(n_1124),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1177),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1120),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1081),
.B(n_1180),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1192),
.A2(n_1108),
.B1(n_1097),
.B2(n_1068),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1090),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1093),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_R g1271 ( 
.A1(n_1082),
.A2(n_1191),
.B1(n_1173),
.B2(n_1140),
.Y(n_1271)
);

BUFx4f_ASAP7_75t_SL g1272 ( 
.A(n_1132),
.Y(n_1272)
);

CKINVDCx6p67_ASAP7_75t_R g1273 ( 
.A(n_1140),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1082),
.A2(n_1191),
.B1(n_1173),
.B2(n_1140),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1126),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1110),
.Y(n_1276)
);

INVx5_ASAP7_75t_L g1277 ( 
.A(n_1082),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1168),
.Y(n_1278)
);

INVx5_ASAP7_75t_L g1279 ( 
.A(n_1098),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1168),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1173),
.A2(n_1191),
.B1(n_1175),
.B2(n_1076),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1175),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1175),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1070),
.A2(n_1134),
.B1(n_1143),
.B2(n_1144),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1145),
.A2(n_1149),
.B1(n_1150),
.B2(n_1160),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1172),
.A2(n_1065),
.B1(n_964),
.B2(n_1195),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1065),
.A2(n_964),
.B1(n_1178),
.B2(n_979),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1077),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1093),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1190),
.B(n_1178),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1065),
.A2(n_1174),
.B1(n_1071),
.B2(n_1186),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1163),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1077),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1083),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_1096),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1065),
.A2(n_1174),
.B1(n_1071),
.B2(n_1186),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1071),
.B1(n_1065),
.B2(n_1178),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1083),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_SL g1299 ( 
.A(n_1096),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1065),
.A2(n_964),
.B1(n_1178),
.B2(n_979),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_R g1301 ( 
.A1(n_1065),
.A2(n_298),
.B1(n_304),
.B2(n_423),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_SL g1302 ( 
.A(n_1153),
.Y(n_1302)
);

INVx4_ASAP7_75t_L g1303 ( 
.A(n_1113),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1163),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1083),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1065),
.A2(n_964),
.B1(n_1167),
.B2(n_1162),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1083),
.Y(n_1307)
);

BUFx12f_ASAP7_75t_L g1308 ( 
.A(n_1163),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1166),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1100),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1301),
.A2(n_1300),
.B1(n_1287),
.B2(n_1291),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1246),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1252),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1260),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1198),
.B(n_1204),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1283),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1283),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1235),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1212),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1203),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_SL g1321 ( 
.A(n_1292),
.B(n_1308),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1238),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1209),
.B(n_1199),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1222),
.B(n_1223),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1287),
.A2(n_1300),
.B1(n_1282),
.B2(n_1208),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1260),
.Y(n_1326)
);

BUFx8_ASAP7_75t_SL g1327 ( 
.A(n_1228),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1277),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1224),
.B(n_1233),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1238),
.Y(n_1330)
);

AO32x2_ASAP7_75t_L g1331 ( 
.A1(n_1274),
.A2(n_1291),
.A3(n_1296),
.B1(n_1220),
.B2(n_1216),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1306),
.A2(n_1201),
.B1(n_1297),
.B2(n_1296),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1277),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1294),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1262),
.B(n_1263),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1236),
.A2(n_1249),
.B(n_1274),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1236),
.A2(n_1281),
.B(n_1199),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1284),
.A2(n_1267),
.B(n_1270),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1240),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1298),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1305),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1208),
.A2(n_1209),
.B1(n_1297),
.B2(n_1275),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1307),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1249),
.A2(n_1290),
.B(n_1216),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1277),
.B(n_1259),
.Y(n_1345)
);

AOI222xp33_ASAP7_75t_L g1346 ( 
.A1(n_1220),
.A2(n_1219),
.B1(n_1290),
.B2(n_1211),
.C1(n_1261),
.C2(n_1218),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1261),
.A2(n_1257),
.B(n_1219),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1271),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1272),
.Y(n_1349)
);

INVx6_ASAP7_75t_SL g1350 ( 
.A(n_1241),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1273),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1280),
.Y(n_1352)
);

AOI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1217),
.A2(n_1286),
.B1(n_1257),
.B2(n_1268),
.C(n_1229),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1269),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1277),
.B(n_1258),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1289),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1289),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1234),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1225),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1205),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1217),
.A2(n_1239),
.B(n_1267),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1215),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1221),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1279),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1258),
.B(n_1247),
.Y(n_1365)
);

INVxp33_ASAP7_75t_L g1366 ( 
.A(n_1309),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1272),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1231),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1288),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1278),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1293),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_SL g1372 ( 
.A1(n_1265),
.A2(n_1266),
.B(n_1239),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1268),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1276),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1232),
.B(n_1244),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1276),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1264),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1264),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1242),
.A2(n_1243),
.B1(n_1256),
.B2(n_1251),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1237),
.A2(n_1279),
.B(n_1285),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1302),
.A2(n_1200),
.B1(n_1248),
.B2(n_1250),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1285),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1255),
.Y(n_1383)
);

OAI21xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1265),
.A2(n_1266),
.B(n_1197),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1202),
.A2(n_1197),
.B(n_1255),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1248),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1254),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1310),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1310),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1241),
.B(n_1253),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1344),
.A2(n_1230),
.B(n_1245),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1332),
.A2(n_1302),
.B1(n_1207),
.B2(n_1210),
.C(n_1213),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1320),
.B(n_1295),
.Y(n_1393)
);

INVx5_ASAP7_75t_L g1394 ( 
.A(n_1364),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1323),
.B(n_1213),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1334),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1361),
.A2(n_1245),
.B(n_1303),
.Y(n_1397)
);

AO32x2_ASAP7_75t_L g1398 ( 
.A1(n_1331),
.A2(n_1227),
.A3(n_1214),
.B1(n_1304),
.B2(n_1299),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_SL g1399 ( 
.A1(n_1383),
.A2(n_1299),
.B(n_1226),
.C(n_1206),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1327),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1318),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1319),
.B(n_1206),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1334),
.Y(n_1403)
);

NOR2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1348),
.B(n_1383),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1346),
.A2(n_1325),
.B(n_1347),
.C(n_1311),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1370),
.B(n_1351),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1370),
.B(n_1351),
.Y(n_1407)
);

AO32x2_ASAP7_75t_L g1408 ( 
.A1(n_1331),
.A2(n_1348),
.A3(n_1358),
.B1(n_1323),
.B2(n_1347),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1311),
.A2(n_1342),
.B1(n_1353),
.B2(n_1331),
.Y(n_1409)
);

AND2x2_ASAP7_75t_SL g1410 ( 
.A(n_1349),
.B(n_1367),
.Y(n_1410)
);

NOR4xp25_ASAP7_75t_SL g1411 ( 
.A(n_1349),
.B(n_1367),
.C(n_1374),
.D(n_1322),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1339),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1323),
.B(n_1330),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1323),
.A2(n_1365),
.B1(n_1336),
.B2(n_1381),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1323),
.A2(n_1365),
.B1(n_1336),
.B2(n_1381),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1359),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1328),
.B(n_1333),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1315),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1323),
.B(n_1373),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1321),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1323),
.A2(n_1368),
.B1(n_1375),
.B2(n_1337),
.Y(n_1421)
);

AO32x2_ASAP7_75t_L g1422 ( 
.A1(n_1331),
.A2(n_1337),
.A3(n_1329),
.B1(n_1324),
.B2(n_1352),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1379),
.A2(n_1331),
.B1(n_1382),
.B2(n_1366),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1382),
.A2(n_1340),
.B1(n_1341),
.B2(n_1343),
.C(n_1312),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_1356),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1387),
.B(n_1345),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_SL g1427 ( 
.A1(n_1341),
.A2(n_1343),
.B(n_1389),
.C(n_1388),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1337),
.A2(n_1350),
.B1(n_1356),
.B2(n_1357),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1380),
.A2(n_1384),
.B(n_1372),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1384),
.A2(n_1385),
.B(n_1338),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1390),
.B(n_1314),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1312),
.B(n_1313),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1380),
.B(n_1386),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1357),
.Y(n_1434)
);

AO32x2_ASAP7_75t_L g1435 ( 
.A1(n_1360),
.A2(n_1371),
.A3(n_1362),
.B1(n_1363),
.B2(n_1369),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1377),
.A2(n_1378),
.B1(n_1376),
.B2(n_1316),
.C(n_1317),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1413),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1434),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1432),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1432),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1418),
.B(n_1355),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1422),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1394),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1422),
.B(n_1355),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1422),
.B(n_1338),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1419),
.B(n_1414),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1419),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1396),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1421),
.B(n_1354),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1417),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1435),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1403),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1393),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1421),
.B(n_1415),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1409),
.A2(n_1350),
.B1(n_1314),
.B2(n_1326),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1425),
.B(n_1424),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_1335),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1408),
.B(n_1374),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1417),
.B(n_1430),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1428),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1428),
.Y(n_1461)
);

INVx3_ASAP7_75t_SL g1462 ( 
.A(n_1420),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1457),
.B(n_1398),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1451),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1462),
.B(n_1410),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1457),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1456),
.B(n_1404),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1444),
.B(n_1398),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1461),
.A2(n_1405),
.B1(n_1409),
.B2(n_1423),
.C(n_1429),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_SL g1470 ( 
.A(n_1443),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1444),
.B(n_1398),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1455),
.A2(n_1423),
.B1(n_1392),
.B2(n_1397),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1451),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1459),
.B(n_1426),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1461),
.A2(n_1402),
.B1(n_1431),
.B2(n_1395),
.C(n_1436),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_L g1477 ( 
.A(n_1460),
.B(n_1454),
.C(n_1449),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1455),
.A2(n_1397),
.B1(n_1391),
.B2(n_1406),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1453),
.B(n_1441),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1437),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1462),
.Y(n_1481)
);

NOR2x1_ASAP7_75t_SL g1482 ( 
.A(n_1450),
.B(n_1395),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1451),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1460),
.B(n_1454),
.C(n_1449),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1441),
.B(n_1426),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1448),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

AND4x1_ASAP7_75t_L g1488 ( 
.A(n_1462),
.B(n_1420),
.C(n_1458),
.D(n_1446),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1441),
.B(n_1411),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1454),
.A2(n_1391),
.B1(n_1406),
.B2(n_1407),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1442),
.A2(n_1407),
.B1(n_1433),
.B2(n_1427),
.C(n_1416),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1452),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1452),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1486),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1470),
.B(n_1468),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1464),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1439),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1463),
.B(n_1447),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1488),
.B(n_1459),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1486),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1477),
.B(n_1439),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1487),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1488),
.B(n_1450),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1464),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1467),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1468),
.B(n_1437),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1484),
.B(n_1439),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1487),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1510)
);

AND2x4_ASAP7_75t_SL g1511 ( 
.A(n_1475),
.B(n_1478),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1484),
.B(n_1440),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1476),
.B(n_1440),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1481),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1480),
.B(n_1440),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1481),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1438),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1489),
.B(n_1445),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1489),
.B(n_1446),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1471),
.B(n_1446),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1481),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1497),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1497),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1521),
.B(n_1471),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1504),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1498),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1502),
.B(n_1469),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1497),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1510),
.B(n_1485),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1505),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1502),
.B(n_1492),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1510),
.B(n_1512),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1505),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1508),
.B(n_1474),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1462),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1501),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1522),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1501),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1505),
.Y(n_1544)
);

INVx5_ASAP7_75t_L g1545 ( 
.A(n_1515),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1495),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1508),
.B(n_1493),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_1482),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1513),
.B(n_1493),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1513),
.B(n_1474),
.Y(n_1550)
);

NOR2x1p5_ASAP7_75t_SL g1551 ( 
.A(n_1505),
.B(n_1483),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1510),
.B(n_1485),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1483),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1495),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1503),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1503),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1504),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1494),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1509),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1496),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1511),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1532),
.B(n_1400),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1532),
.B(n_1542),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1546),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1546),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1537),
.B(n_1506),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1554),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1528),
.B(n_1522),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1558),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1531),
.B(n_1515),
.C(n_1517),
.Y(n_1570)
);

NAND4xp25_ASAP7_75t_L g1571 ( 
.A(n_1560),
.B(n_1496),
.C(n_1518),
.D(n_1491),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1528),
.B(n_1512),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1554),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1542),
.B(n_1507),
.Y(n_1574)
);

NAND3x1_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1520),
.C(n_1519),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1561),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1531),
.B(n_1528),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1555),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1553),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1401),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1529),
.B(n_1520),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1537),
.B(n_1518),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1537),
.B(n_1516),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1556),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1553),
.B(n_1516),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1540),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1540),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1561),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1561),
.B(n_1511),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1558),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1527),
.B(n_1520),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1556),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1527),
.B(n_1499),
.Y(n_1596)
);

AOI32xp33_ASAP7_75t_L g1597 ( 
.A1(n_1563),
.A2(n_1579),
.A3(n_1519),
.B1(n_1583),
.B2(n_1558),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1562),
.B(n_1560),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1564),
.Y(n_1599)
);

OAI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1563),
.A2(n_1539),
.B1(n_1525),
.B2(n_1550),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1562),
.A2(n_1500),
.B(n_1543),
.C(n_1541),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1589),
.B(n_1545),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1570),
.B(n_1576),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1592),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1589),
.A2(n_1500),
.B(n_1543),
.C(n_1541),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1592),
.B(n_1548),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1527),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1575),
.A2(n_1594),
.B1(n_1584),
.B2(n_1592),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1534),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1534),
.Y(n_1613)
);

OAI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1571),
.A2(n_1545),
.B(n_1530),
.C(n_1557),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1579),
.B(n_1534),
.Y(n_1615)
);

AOI211xp5_ASAP7_75t_L g1616 ( 
.A1(n_1577),
.A2(n_1530),
.B(n_1557),
.C(n_1548),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1552),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1575),
.A2(n_1473),
.B1(n_1519),
.B2(n_1490),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1590),
.A2(n_1574),
.B(n_1566),
.C(n_1595),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1573),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1593),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1601),
.A2(n_1557),
.B(n_1530),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1605),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1618),
.A2(n_1473),
.B1(n_1511),
.B2(n_1490),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1621),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1610),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1599),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1613),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1617),
.B(n_1593),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1602),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1600),
.B(n_1572),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1604),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1611),
.Y(n_1633)
);

AOI21xp33_ASAP7_75t_L g1634 ( 
.A1(n_1601),
.A2(n_1606),
.B(n_1619),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1614),
.A2(n_1557),
.B1(n_1530),
.B2(n_1478),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1598),
.A2(n_1557),
.B1(n_1582),
.B2(n_1581),
.Y(n_1636)
);

NOR2xp67_ASAP7_75t_SL g1637 ( 
.A(n_1607),
.B(n_1545),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1597),
.A2(n_1588),
.B(n_1596),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1606),
.A2(n_1580),
.B(n_1578),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1619),
.A2(n_1547),
.B(n_1536),
.Y(n_1640)
);

AOI21xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1634),
.A2(n_1609),
.B(n_1603),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1632),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1634),
.A2(n_1631),
.B1(n_1640),
.B2(n_1639),
.C(n_1625),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1628),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1631),
.Y(n_1645)
);

NOR3xp33_ASAP7_75t_L g1646 ( 
.A(n_1623),
.B(n_1615),
.C(n_1620),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1629),
.Y(n_1647)
);

O2A1O1Ixp5_ASAP7_75t_L g1648 ( 
.A1(n_1637),
.A2(n_1612),
.B(n_1608),
.C(n_1587),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1626),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1624),
.A2(n_1551),
.B(n_1616),
.C(n_1550),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1627),
.B(n_1586),
.Y(n_1651)
);

XNOR2xp5_ASAP7_75t_L g1652 ( 
.A(n_1636),
.B(n_1412),
.Y(n_1652)
);

OAI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1643),
.A2(n_1622),
.B(n_1638),
.C(n_1635),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1642),
.B(n_1630),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1652),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1649),
.Y(n_1656)
);

NAND3x1_ASAP7_75t_L g1657 ( 
.A(n_1646),
.B(n_1633),
.C(n_1552),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1645),
.B(n_1533),
.C(n_1526),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1644),
.B(n_1548),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1647),
.B(n_1552),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1641),
.B(n_1545),
.C(n_1585),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1651),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1651),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1648),
.Y(n_1664)
);

OAI21xp33_ASAP7_75t_L g1665 ( 
.A1(n_1653),
.A2(n_1650),
.B(n_1517),
.Y(n_1665)
);

NOR3xp33_ASAP7_75t_SL g1666 ( 
.A(n_1654),
.B(n_1465),
.C(n_1536),
.Y(n_1666)
);

AOI221x1_ASAP7_75t_L g1667 ( 
.A1(n_1658),
.A2(n_1526),
.B1(n_1533),
.B2(n_1535),
.C(n_1559),
.Y(n_1667)
);

NOR3xp33_ASAP7_75t_L g1668 ( 
.A(n_1663),
.B(n_1656),
.C(n_1661),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_L g1669 ( 
.A(n_1664),
.B(n_1660),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1665),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1666),
.A2(n_1659),
.B1(n_1525),
.B2(n_1550),
.C(n_1539),
.Y(n_1671)
);

OAI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1667),
.A2(n_1657),
.B(n_1545),
.C(n_1515),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1663),
.A2(n_1545),
.B1(n_1548),
.B2(n_1547),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1670),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1668),
.A2(n_1671),
.B1(n_1672),
.B2(n_1673),
.C(n_1669),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1669),
.A2(n_1545),
.B1(n_1549),
.B2(n_1539),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_L g1677 ( 
.A(n_1669),
.B(n_1548),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1670),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1674),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1678),
.B(n_1526),
.C(n_1533),
.Y(n_1680)
);

INVxp67_ASAP7_75t_SL g1681 ( 
.A(n_1677),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1681),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1682),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1679),
.B1(n_1675),
.B2(n_1676),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1683),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1685),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1684),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1687),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1686),
.A2(n_1680),
.B1(n_1538),
.B2(n_1524),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1688),
.A2(n_1538),
.B(n_1544),
.Y(n_1690)
);

OAI21xp33_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1689),
.B(n_1517),
.Y(n_1691)
);

XOR2xp5_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1399),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1524),
.B1(n_1523),
.B2(n_1544),
.C(n_1538),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1525),
.B(n_1523),
.C(n_1524),
.Y(n_1694)
);


endmodule