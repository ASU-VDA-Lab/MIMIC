module fake_jpeg_28171_n_68 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_55;
wire n_27;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_25;
wire n_56;
wire n_31;
wire n_67;
wire n_43;
wire n_37;
wire n_50;
wire n_29;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_2),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_44),
.B(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_13),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_25),
.C(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_50),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_54),
.B(n_20),
.Y(n_57)
);

OAI22x1_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_34),
.B1(n_26),
.B2(n_37),
.Y(n_58)
);

AOI322xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_59),
.A3(n_34),
.B1(n_39),
.B2(n_45),
.C1(n_49),
.C2(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_42),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_24),
.B1(n_40),
.B2(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_51),
.Y(n_63)
);

OA21x2_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_46),
.B(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_29),
.B(n_27),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_65),
.B(n_28),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_47),
.Y(n_68)
);


endmodule