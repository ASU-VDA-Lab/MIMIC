module real_aes_263_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_671;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_283;
wire n_314;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_0), .A2(n_210), .B1(n_377), .B2(n_378), .Y(n_376) );
AO222x2_ASAP7_75t_SL g517 ( .A1(n_1), .A2(n_33), .B1(n_146), .B2(n_485), .C1(n_518), .C2(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_2), .A2(n_214), .B1(n_392), .B2(n_393), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_3), .A2(n_230), .B1(n_343), .B2(n_347), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_4), .A2(n_25), .B1(n_302), .B2(n_523), .Y(n_522) );
AO22x2_ASAP7_75t_L g292 ( .A1(n_5), .A2(n_171), .B1(n_282), .B2(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g667 ( .A(n_5), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_6), .A2(n_52), .B1(n_630), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_7), .A2(n_113), .B1(n_343), .B2(n_349), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_8), .A2(n_208), .B1(n_343), .B2(n_347), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_9), .A2(n_65), .B1(n_424), .B2(n_426), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_10), .A2(n_238), .B1(n_450), .B2(n_453), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_11), .A2(n_235), .B1(n_336), .B2(n_633), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_12), .A2(n_157), .B1(n_333), .B2(n_389), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_13), .A2(n_67), .B1(n_393), .B2(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_14), .A2(n_101), .B1(n_325), .B2(n_518), .Y(n_622) );
OA22x2_ASAP7_75t_L g495 ( .A1(n_15), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_15), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_16), .A2(n_88), .B1(n_303), .B2(n_431), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_17), .A2(n_27), .B1(n_453), .B2(n_455), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_18), .A2(n_42), .B1(n_609), .B2(n_611), .Y(n_608) );
AO22x2_ASAP7_75t_L g289 ( .A1(n_19), .A2(n_68), .B1(n_282), .B2(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_19), .B(n_666), .Y(n_665) );
XOR2x2_ASAP7_75t_L g594 ( .A(n_20), .B(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_21), .A2(n_50), .B1(n_392), .B2(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_22), .A2(n_159), .B1(n_329), .B2(n_332), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_23), .A2(n_48), .B1(n_308), .B2(n_312), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_24), .A2(n_130), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_26), .A2(n_183), .B1(n_383), .B2(n_448), .Y(n_577) );
AO222x2_ASAP7_75t_SL g678 ( .A1(n_28), .A2(n_145), .B1(n_239), .B2(n_276), .C1(n_427), .C2(n_651), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_29), .A2(n_133), .B1(n_409), .B2(n_411), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g254 ( .A1(n_30), .A2(n_255), .B(n_263), .C(n_669), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_31), .A2(n_54), .B1(n_296), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_32), .A2(n_85), .B1(n_389), .B2(n_390), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_34), .A2(n_61), .B1(n_450), .B2(n_451), .Y(n_506) );
AOI222xp33_ASAP7_75t_L g500 ( .A1(n_35), .A2(n_211), .B1(n_245), .B2(n_367), .C1(n_377), .C2(n_462), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_36), .A2(n_188), .B1(n_383), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_37), .A2(n_252), .B1(n_392), .B2(n_393), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_38), .A2(n_241), .B1(n_411), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_39), .A2(n_198), .B1(n_389), .B2(n_407), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_40), .A2(n_221), .B1(n_343), .B2(n_347), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_41), .A2(n_116), .B1(n_392), .B2(n_393), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_43), .A2(n_175), .B1(n_385), .B2(n_393), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_44), .A2(n_234), .B1(n_392), .B2(n_393), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_45), .A2(n_165), .B1(n_374), .B2(n_375), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_46), .A2(n_237), .B1(n_352), .B2(n_356), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_47), .A2(n_182), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_49), .A2(n_142), .B1(n_421), .B2(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_51), .A2(n_181), .B1(n_563), .B2(n_564), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_53), .A2(n_248), .B1(n_370), .B2(n_504), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_55), .A2(n_89), .B1(n_295), .B2(n_302), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_56), .A2(n_131), .B1(n_523), .B2(n_621), .Y(n_709) );
AO222x2_ASAP7_75t_L g459 ( .A1(n_57), .A2(n_69), .B1(n_173), .B2(n_367), .C1(n_370), .C2(n_371), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_58), .A2(n_144), .B1(n_598), .B2(n_637), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_59), .B(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_60), .A2(n_186), .B1(n_358), .B2(n_392), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_62), .A2(n_98), .B1(n_424), .B2(n_426), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_63), .A2(n_121), .B1(n_336), .B2(n_451), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_64), .A2(n_176), .B1(n_451), .B2(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_66), .A2(n_111), .B1(n_378), .B2(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_70), .A2(n_151), .B1(n_374), .B2(n_375), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_71), .A2(n_75), .B1(n_444), .B2(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_72), .A2(n_231), .B1(n_370), .B2(n_371), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_73), .A2(n_247), .B1(n_383), .B2(n_448), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_74), .A2(n_141), .B1(n_425), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_76), .A2(n_99), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_77), .A2(n_156), .B1(n_451), .B2(n_471), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_78), .A2(n_206), .B1(n_386), .B2(n_528), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_79), .A2(n_122), .B1(n_406), .B2(n_407), .Y(n_599) );
INVx3_ASAP7_75t_L g282 ( .A(n_80), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_81), .A2(n_250), .B1(n_431), .B2(n_675), .Y(n_674) );
AO21x2_ASAP7_75t_L g694 ( .A1(n_82), .A2(n_695), .B(n_710), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_82), .B(n_697), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_82), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_83), .A2(n_87), .B1(n_424), .B2(n_426), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_84), .A2(n_218), .B1(n_413), .B2(n_607), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_86), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_90), .A2(n_163), .B1(n_450), .B2(n_451), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_91), .A2(n_105), .B1(n_421), .B2(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_92), .A2(n_168), .B1(n_453), .B2(n_455), .Y(n_472) );
OA22x2_ASAP7_75t_L g399 ( .A1(n_93), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_93), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_94), .B(n_417), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_95), .A2(n_117), .B1(n_406), .B2(n_407), .Y(n_405) );
INVx1_ASAP7_75t_SL g283 ( .A(n_96), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_96), .B(n_120), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_97), .A2(n_107), .B1(n_215), .B2(n_424), .C1(n_426), .C2(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g262 ( .A(n_100), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_102), .A2(n_671), .B1(n_689), .B2(n_690), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_102), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_103), .A2(n_205), .B1(n_309), .B2(n_427), .Y(n_487) );
XOR2x2_ASAP7_75t_L g641 ( .A(n_104), .B(n_642), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_106), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_108), .A2(n_123), .B1(n_523), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_109), .A2(n_253), .B1(n_389), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_110), .A2(n_127), .B1(n_409), .B2(n_633), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_112), .A2(n_224), .B1(n_374), .B2(n_375), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_114), .B(n_275), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_115), .A2(n_200), .B1(n_343), .B2(n_541), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_118), .A2(n_207), .B1(n_450), .B2(n_451), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_119), .B(n_367), .Y(n_441) );
AO22x2_ASAP7_75t_L g285 ( .A1(n_120), .A2(n_178), .B1(n_282), .B2(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_124), .B(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_125), .A2(n_150), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_126), .A2(n_236), .B1(n_604), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_128), .A2(n_199), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_129), .A2(n_143), .B1(n_611), .B2(n_685), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_132), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_134), .A2(n_219), .B1(n_336), .B2(n_339), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_135), .A2(n_140), .B1(n_383), .B2(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_136), .Y(n_368) );
INVx1_ASAP7_75t_L g284 ( .A(n_137), .Y(n_284) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_138), .A2(n_185), .B1(n_382), .B2(n_383), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_139), .A2(n_161), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_147), .A2(n_217), .B1(n_375), .B2(n_431), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_148), .A2(n_244), .B1(n_382), .B2(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_149), .B(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_152), .A2(n_216), .B1(n_519), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_153), .A2(n_203), .B1(n_358), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_154), .A2(n_242), .B1(n_374), .B2(n_375), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_155), .A2(n_169), .B1(n_383), .B2(n_448), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_158), .A2(n_201), .B1(n_627), .B2(n_630), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_160), .A2(n_222), .B1(n_429), .B2(n_433), .Y(n_428) );
XNOR2x1_ASAP7_75t_L g438 ( .A(n_162), .B(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_164), .A2(n_192), .B1(n_413), .B2(n_414), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_166), .A2(n_233), .B1(n_374), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_167), .A2(n_191), .B1(n_413), .B2(n_607), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_170), .A2(n_193), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_172), .A2(n_213), .B1(n_319), .B2(n_323), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_174), .A2(n_227), .B1(n_313), .B2(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_177), .B(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_179), .A2(n_187), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_180), .A2(n_226), .B1(n_370), .B2(n_504), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_184), .Y(n_529) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_189), .A2(n_515), .B(n_542), .Y(n_514) );
INVx1_ASAP7_75t_L g544 ( .A(n_189), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_190), .B(n_582), .Y(n_656) );
AO22x2_ASAP7_75t_L g573 ( .A1(n_194), .A2(n_574), .B1(n_586), .B2(n_587), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_194), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_195), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g663 ( .A(n_195), .Y(n_663) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_196), .B(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_197), .A2(n_228), .B1(n_377), .B2(n_462), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_202), .A2(n_212), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
AND2x2_ASAP7_75t_R g692 ( .A(n_204), .B(n_663), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_209), .A2(n_271), .B1(n_272), .B2(n_359), .Y(n_270) );
INVx1_ASAP7_75t_L g359 ( .A(n_209), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_220), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g394 ( .A(n_223), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_225), .A2(n_251), .B1(n_377), .B2(n_462), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_229), .A2(n_240), .B1(n_392), .B2(n_393), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_232), .B(n_485), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_243), .A2(n_246), .B1(n_444), .B2(n_462), .Y(n_584) );
OA22x2_ASAP7_75t_L g473 ( .A1(n_249), .A2(n_474), .B1(n_475), .B2(n_489), .Y(n_473) );
INVx1_ASAP7_75t_L g489 ( .A(n_249), .Y(n_489) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g716 ( .A(n_258), .B(n_260), .Y(n_716) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_259), .B(n_663), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_510), .B1(n_658), .B2(n_659), .C(n_660), .Y(n_263) );
INVx1_ASAP7_75t_L g659 ( .A(n_264), .Y(n_659) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_396), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI22x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B1(n_360), .B2(n_395), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_327), .Y(n_272) );
NAND4xp25_ASAP7_75t_SL g273 ( .A(n_274), .B(n_294), .C(n_307), .D(n_318), .Y(n_273) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx3_ASAP7_75t_SL g419 ( .A(n_277), .Y(n_419) );
INVx3_ASAP7_75t_L g485 ( .A(n_277), .Y(n_485) );
INVx4_ASAP7_75t_SL g582 ( .A(n_277), .Y(n_582) );
INVx4_ASAP7_75t_SL g613 ( .A(n_277), .Y(n_613) );
INVx6_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_287), .Y(n_278) );
AND2x4_ASAP7_75t_L g304 ( .A(n_279), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g325 ( .A(n_279), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g367 ( .A(n_279), .B(n_287), .Y(n_367) );
AND2x2_ASAP7_75t_L g375 ( .A(n_279), .B(n_305), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_279), .B(n_326), .Y(n_378) );
AND2x2_ASAP7_75t_L g462 ( .A(n_279), .B(n_326), .Y(n_462) );
AND2x2_ASAP7_75t_L g502 ( .A(n_279), .B(n_305), .Y(n_502) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_285), .Y(n_279) );
AND2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_280), .Y(n_317) );
INVx2_ASAP7_75t_L g322 ( .A(n_280), .Y(n_322) );
OAI22x1_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_283), .B2(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g286 ( .A(n_282), .Y(n_286) );
INVx2_ASAP7_75t_L g290 ( .A(n_282), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_282), .Y(n_293) );
INVx2_ASAP7_75t_L g301 ( .A(n_285), .Y(n_301) );
AND2x2_ASAP7_75t_L g321 ( .A(n_285), .B(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g350 ( .A(n_285), .Y(n_350) );
AND2x4_ASAP7_75t_L g331 ( .A(n_287), .B(n_300), .Y(n_331) );
AND2x4_ASAP7_75t_L g338 ( .A(n_287), .B(n_334), .Y(n_338) );
AND2x2_ASAP7_75t_L g355 ( .A(n_287), .B(n_321), .Y(n_355) );
AND2x6_ASAP7_75t_L g392 ( .A(n_287), .B(n_321), .Y(n_392) );
AND2x2_ASAP7_75t_L g450 ( .A(n_287), .B(n_300), .Y(n_450) );
AND2x2_ASAP7_75t_L g455 ( .A(n_287), .B(n_334), .Y(n_455) );
AND2x2_ASAP7_75t_L g471 ( .A(n_287), .B(n_300), .Y(n_471) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g299 ( .A(n_289), .Y(n_299) );
AND2x4_ASAP7_75t_L g311 ( .A(n_289), .B(n_291), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_292), .Y(n_316) );
INVxp67_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g298 ( .A(n_292), .B(n_299), .Y(n_298) );
BUFx6f_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx3_ASAP7_75t_L g432 ( .A(n_297), .Y(n_432) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_297), .Y(n_558) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
AND2x4_ASAP7_75t_L g341 ( .A(n_298), .B(n_334), .Y(n_341) );
AND2x2_ASAP7_75t_L g346 ( .A(n_298), .B(n_321), .Y(n_346) );
AND2x4_ASAP7_75t_L g374 ( .A(n_298), .B(n_300), .Y(n_374) );
AND2x6_ASAP7_75t_L g393 ( .A(n_298), .B(n_334), .Y(n_393) );
AND2x2_ASAP7_75t_L g448 ( .A(n_298), .B(n_321), .Y(n_448) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_298), .B(n_321), .Y(n_467) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
AND2x2_ASAP7_75t_L g310 ( .A(n_300), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g370 ( .A(n_300), .B(n_311), .Y(n_370) );
AND2x4_ASAP7_75t_L g334 ( .A(n_301), .B(n_322), .Y(n_334) );
BUFx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g435 ( .A(n_304), .Y(n_435) );
BUFx3_ASAP7_75t_L g559 ( .A(n_304), .Y(n_559) );
BUFx4f_ASAP7_75t_L g602 ( .A(n_304), .Y(n_602) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g425 ( .A(n_310), .Y(n_425) );
INVx2_ASAP7_75t_L g652 ( .A(n_310), .Y(n_652) );
AND2x4_ASAP7_75t_L g320 ( .A(n_311), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g358 ( .A(n_311), .B(n_334), .Y(n_358) );
AND2x2_ASAP7_75t_L g377 ( .A(n_311), .B(n_321), .Y(n_377) );
AND2x2_ASAP7_75t_L g444 ( .A(n_311), .B(n_321), .Y(n_444) );
AND2x2_ASAP7_75t_L g453 ( .A(n_311), .B(n_334), .Y(n_453) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g427 ( .A(n_314), .Y(n_427) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx12f_ASAP7_75t_L g552 ( .A(n_315), .Y(n_552) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x4_ASAP7_75t_L g333 ( .A(n_316), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g349 ( .A(n_316), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_316), .B(n_317), .Y(n_371) );
AND2x4_ASAP7_75t_L g383 ( .A(n_316), .B(n_350), .Y(n_383) );
AND2x4_ASAP7_75t_L g451 ( .A(n_316), .B(n_334), .Y(n_451) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_316), .B(n_317), .Y(n_504) );
BUFx4f_ASAP7_75t_SL g421 ( .A(n_319), .Y(n_421) );
BUFx2_ASAP7_75t_L g518 ( .A(n_319), .Y(n_518) );
BUFx2_ASAP7_75t_L g707 ( .A(n_319), .Y(n_707) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g555 ( .A(n_320), .Y(n_555) );
BUFx3_ASAP7_75t_L g677 ( .A(n_320), .Y(n_677) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g422 ( .A(n_324), .Y(n_422) );
INVx2_ASAP7_75t_L g519 ( .A(n_324), .Y(n_519) );
INVx2_ASAP7_75t_L g556 ( .A(n_324), .Y(n_556) );
INVx2_ASAP7_75t_SL g604 ( .A(n_324), .Y(n_604) );
INVx6_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_328), .B(n_335), .C(n_342), .D(n_351), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g406 ( .A(n_330), .Y(n_406) );
INVx1_ASAP7_75t_SL g636 ( .A(n_330), .Y(n_636) );
INVx2_ASAP7_75t_L g681 ( .A(n_330), .Y(n_681) );
INVx6_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g389 ( .A(n_331), .Y(n_389) );
BUFx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g390 ( .A(n_333), .Y(n_390) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_333), .Y(n_407) );
BUFx2_ASAP7_75t_SL g637 ( .A(n_333), .Y(n_637) );
INVx2_ASAP7_75t_L g410 ( .A(n_336), .Y(n_410) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_336), .Y(n_598) );
INVx4_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_SL g385 ( .A(n_337), .Y(n_385) );
INVx2_ASAP7_75t_L g528 ( .A(n_337), .Y(n_528) );
INVx3_ASAP7_75t_L g648 ( .A(n_337), .Y(n_648) );
INVx8_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g414 ( .A(n_340), .Y(n_414) );
INVx2_ASAP7_75t_SL g539 ( .A(n_340), .Y(n_539) );
INVx2_ASAP7_75t_L g567 ( .A(n_340), .Y(n_567) );
INVx1_ASAP7_75t_SL g607 ( .A(n_340), .Y(n_607) );
INVx2_ASAP7_75t_L g630 ( .A(n_340), .Y(n_630) );
INVx8_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g563 ( .A(n_345), .Y(n_563) );
INVx2_ASAP7_75t_L g610 ( .A(n_345), .Y(n_610) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g382 ( .A(n_346), .Y(n_382) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_346), .Y(n_685) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g541 ( .A(n_348), .Y(n_541) );
INVx2_ASAP7_75t_L g564 ( .A(n_348), .Y(n_564) );
INVx3_ASAP7_75t_L g611 ( .A(n_348), .Y(n_611) );
INVx5_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g481 ( .A(n_349), .Y(n_481) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_SL g413 ( .A(n_354), .Y(n_413) );
INVx3_ASAP7_75t_L g538 ( .A(n_354), .Y(n_538) );
INVx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g566 ( .A(n_355), .Y(n_566) );
BUFx2_ASAP7_75t_L g629 ( .A(n_355), .Y(n_629) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
BUFx3_ASAP7_75t_L g532 ( .A(n_358), .Y(n_532) );
INVx2_ASAP7_75t_L g683 ( .A(n_358), .Y(n_683) );
INVx1_ASAP7_75t_SL g395 ( .A(n_360), .Y(n_395) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
XOR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_394), .Y(n_362) );
NAND2x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_379), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_372), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_368), .B(n_369), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
NOR2x1_ASAP7_75t_L g379 ( .A(n_380), .B(n_387), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_386), .Y(n_411) );
INVx2_ASAP7_75t_L g634 ( .A(n_386), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_391), .Y(n_387) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_390), .Y(n_535) );
XOR2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_493), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_436), .B2(n_492), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_415), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .C(n_408), .D(n_412), .Y(n_403) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND4xp25_ASAP7_75t_SL g415 ( .A(n_416), .B(n_420), .C(n_423), .D(n_428), .Y(n_415) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp33_ASAP7_75t_SL g549 ( .A1(n_418), .A2(n_550), .B(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g524 ( .A(n_432), .Y(n_524) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g675 ( .A(n_435), .Y(n_675) );
INVx1_ASAP7_75t_L g492 ( .A(n_436), .Y(n_492) );
OA22x2_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_473), .B1(n_490), .B2(n_491), .Y(n_436) );
INVx1_ASAP7_75t_L g491 ( .A(n_437), .Y(n_491) );
XOR2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_456), .Y(n_437) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_446), .Y(n_439) );
NAND4xp25_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .C(n_443), .D(n_445), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g446 ( .A(n_447), .B(n_449), .C(n_452), .D(n_454), .Y(n_446) );
NAND2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_464), .Y(n_457) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g490 ( .A(n_473), .Y(n_490) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .C(n_482), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .C(n_487), .D(n_488), .Y(n_483) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .C(n_503), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .C(n_508), .D(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g658 ( .A(n_510), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_591), .B1(n_592), .B2(n_657), .Y(n_510) );
INVx1_ASAP7_75t_L g657 ( .A(n_511), .Y(n_657) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_545), .B1(n_589), .B2(n_590), .Y(n_513) );
INVx1_ASAP7_75t_L g589 ( .A(n_514), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .C(n_536), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .Y(n_516) );
NOR4xp25_ASAP7_75t_L g542 ( .A(n_517), .B(n_520), .C(n_526), .D(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
OAI221xp5_ASAP7_75t_SL g526 ( .A1(n_527), .A2(n_529), .B1(n_530), .B2(n_533), .C(n_534), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_536), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g590 ( .A(n_545), .Y(n_590) );
OAI22x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_572), .B1(n_573), .B2(n_588), .Y(n_545) );
INVx2_ASAP7_75t_L g588 ( .A(n_546), .Y(n_588) );
XNOR2x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_571), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_560), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
BUFx6f_ASAP7_75t_SL g621 ( .A(n_559), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_568), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
BUFx3_ASAP7_75t_L g701 ( .A(n_566), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g587 ( .A(n_574), .Y(n_587) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .C(n_578), .D(n_579), .Y(n_575) );
NAND4xp25_ASAP7_75t_SL g580 ( .A(n_581), .B(n_583), .C(n_584), .D(n_585), .Y(n_580) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_614), .B2(n_615), .Y(n_592) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND4xp75_ASAP7_75t_SL g595 ( .A(n_596), .B(n_600), .C(n_605), .D(n_612), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_617), .B1(n_638), .B2(n_639), .Y(n_615) );
INVx4_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2x1_ASAP7_75t_L g618 ( .A(n_619), .B(n_625), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .C(n_623), .D(n_624), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_631), .C(n_632), .D(n_635), .Y(n_625) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_649), .C(n_654), .Y(n_642) );
NAND4xp25_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .C(n_646), .D(n_647), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_662), .B(n_665), .Y(n_713) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OAI222xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_691), .B1(n_693), .B2(n_711), .C1(n_714), .C2(n_717), .Y(n_669) );
INVx1_ASAP7_75t_L g690 ( .A(n_671), .Y(n_690) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR4xp75_ASAP7_75t_L g672 ( .A(n_673), .B(n_678), .C(n_679), .D(n_686), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_704), .Y(n_697) );
NAND4xp25_ASAP7_75t_SL g698 ( .A(n_699), .B(n_700), .C(n_702), .D(n_703), .Y(n_698) );
NAND4xp25_ASAP7_75t_SL g704 ( .A(n_705), .B(n_706), .C(n_708), .D(n_709), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
CKINVDCx6p67_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
endmodule