module fake_jpeg_14960_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_57),
.B1(n_43),
.B2(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_48),
.Y(n_90)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_30),
.B1(n_26),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_100)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_30),
.B1(n_32),
.B2(n_20),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_33),
.B1(n_18),
.B2(n_26),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_26),
.B1(n_33),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_44),
.B1(n_39),
.B2(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

INVxp67_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_95),
.B(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_73),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_93),
.B1(n_51),
.B2(n_48),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_27),
.B(n_25),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_58),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_43),
.B1(n_21),
.B2(n_23),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_80),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_97),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_37),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_19),
.Y(n_120)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_43),
.B1(n_21),
.B2(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_27),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_91),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_35),
.B1(n_40),
.B2(n_17),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_16),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_16),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_102),
.B(n_40),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_103),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_35),
.B1(n_17),
.B2(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_59),
.B1(n_60),
.B2(n_48),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_31),
.B(n_1),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_78),
.B(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_117),
.B1(n_118),
.B2(n_94),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_127),
.B1(n_128),
.B2(n_0),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_35),
.B1(n_47),
.B2(n_31),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_124),
.B1(n_71),
.B2(n_99),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_35),
.B1(n_47),
.B2(n_11),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_82),
.B1(n_81),
.B2(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_102),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_19),
.C(n_22),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_126),
.C(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_47),
.B1(n_22),
.B2(n_16),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_22),
.C(n_40),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_93),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_135),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_79),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_141),
.B(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_74),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_144),
.Y(n_175)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_78),
.B(n_83),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_92),
.C(n_94),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_135),
.C(n_134),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_93),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_147),
.B(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_84),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_90),
.B1(n_96),
.B2(n_101),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_93),
.B1(n_101),
.B2(n_90),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_163),
.B(n_127),
.C(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_75),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_71),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_113),
.B(n_92),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_155),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_85),
.B1(n_87),
.B2(n_80),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_161),
.B1(n_119),
.B2(n_11),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_132),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_156),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_109),
.B(n_117),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_162),
.B1(n_128),
.B2(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_8),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_40),
.B1(n_1),
.B2(n_3),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_0),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_10),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_171),
.B(n_179),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_176),
.C(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_139),
.C(n_144),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_123),
.B(n_112),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_122),
.C(n_133),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_185),
.A2(n_186),
.B(n_187),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_143),
.B(n_138),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_114),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_143),
.A2(n_108),
.B(n_111),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_195),
.B(n_3),
.Y(n_212)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_124),
.C(n_131),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_12),
.C(n_13),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_131),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_196),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_154),
.B(n_163),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_131),
.A3(n_119),
.B1(n_5),
.B2(n_6),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_6),
.B1(n_7),
.B2(n_194),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_146),
.B1(n_163),
.B2(n_158),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_210),
.B1(n_220),
.B2(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_170),
.B(n_140),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_212),
.B(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_174),
.A2(n_40),
.B1(n_4),
.B2(n_5),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_217),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_185),
.B1(n_182),
.B2(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_215),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_171),
.B(n_5),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_191),
.B1(n_183),
.B2(n_179),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_7),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_170),
.B(n_7),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_180),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_168),
.A2(n_196),
.B1(n_195),
.B2(n_177),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_177),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_188),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_187),
.B1(n_190),
.B2(n_186),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_184),
.B1(n_172),
.B2(n_176),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_236),
.B1(n_238),
.B2(n_213),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_167),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_208),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_169),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_173),
.B1(n_191),
.B2(n_192),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_166),
.B1(n_212),
.B2(n_222),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_166),
.B(n_222),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_245),
.B(n_218),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_204),
.B(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_202),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_200),
.C(n_217),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_255),
.B1(n_243),
.B2(n_235),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_200),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_223),
.C(n_199),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_236),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_243),
.B(n_246),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_254),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_213),
.B1(n_208),
.B2(n_210),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_260),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_202),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_262),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_238),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_245),
.B1(n_264),
.B2(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_270),
.B(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_278),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_277),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_257),
.B1(n_264),
.B2(n_261),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_290),
.B1(n_265),
.B2(n_266),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_276),
.B1(n_273),
.B2(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_232),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_251),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_263),
.B1(n_235),
.B2(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_279),
.B1(n_283),
.B2(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_232),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_299),
.C(n_288),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_266),
.B(n_252),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_272),
.B(n_250),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_302),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_299),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_282),
.B(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_298),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_293),
.B(n_294),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_308),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_292),
.C(n_248),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_307),
.C(n_304),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_313),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_272),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_241),
.Y(n_316)
);


endmodule