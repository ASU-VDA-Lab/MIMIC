module real_jpeg_5459_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_1),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_1),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_1),
.A2(n_139),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_1),
.A2(n_48),
.B1(n_139),
.B2(n_278),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_1),
.A2(n_139),
.B1(n_300),
.B2(n_303),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_3),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_47),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_3),
.A2(n_47),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_126),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_263),
.B(n_265),
.C(n_269),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_3),
.B(n_290),
.C(n_292),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_77),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_3),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_3),
.B(n_61),
.Y(n_329)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_5),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_5),
.Y(n_317)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_6),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_6),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_8),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_8),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_9),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_38),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_38),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_10),
.A2(n_38),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_21),
.B1(n_193),
.B2(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_230),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_228),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_200),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_16),
.B(n_200),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.C(n_177),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_17),
.B(n_177),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_75),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_18),
.B(n_107),
.C(n_141),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_19),
.B(n_39),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B(n_35),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_20),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_31),
.B(n_36),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_31),
.A2(n_183),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_31),
.B(n_183),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_31),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_35),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_35),
.B(n_298),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_69),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_40),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_51),
.Y(n_40)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_41),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_45),
.Y(n_196)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_46),
.Y(n_198)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_47),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_138),
.B(n_159),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_47),
.A2(n_266),
.B(n_268),
.Y(n_265)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_51),
.B(n_70),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_51),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_51),
.B(n_277),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_61),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_61),
.B(n_277),
.Y(n_294)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_65),
.Y(n_303)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_68),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_68),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_69),
.A2(n_192),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_69),
.B(n_276),
.Y(n_305)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_107),
.B1(n_141),
.B2(n_142),
.Y(n_75)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_102),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_77),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_77),
.B(n_171),
.Y(n_252)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_169),
.Y(n_168)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_81),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_85),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_86),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_86),
.B(n_102),
.Y(n_217)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_87),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_94),
.Y(n_271)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_102),
.Y(n_169)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_136),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_126),
.Y(n_145)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_114),
.B(n_209),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_126),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_120),
.B2(n_124),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_126),
.B(n_209),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_134),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_136),
.B(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_143),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_166),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_144),
.B(n_166),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_147),
.B(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_148),
.B(n_152),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.A3(n_157),
.B1(n_158),
.B2(n_162),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_211),
.Y(n_237)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_190),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_186),
.Y(n_302)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_189),
.B(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B(n_199),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_191),
.A2(n_225),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_191),
.B(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_199),
.B(n_294),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_227),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_218),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_217),
.B(n_252),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_219),
.A2(n_226),
.B1(n_262),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_350),
.B(n_361),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_281),
.B(n_349),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_257),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_233),
.B(n_257),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_242),
.B2(n_243),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_236),
.B(n_242),
.C(n_244),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_240),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_241),
.B(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_245),
.B(n_248),
.C(n_254),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.C(n_272),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_258),
.B(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_261),
.A2(n_272),
.B1(n_273),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_261),
.Y(n_346)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_343),
.B(n_348),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_333),
.B(n_342),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_309),
.B(n_332),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_295),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_295),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_287),
.B1(n_293),
.B2(n_312),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_304),
.Y(n_295)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_307),
.C(n_335),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_318),
.B(n_331),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_313),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_327),
.B(n_330),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_326),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_336),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_347),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_358),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_353),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_353),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_359),
.Y(n_363)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_355),
.CI(n_356),
.CON(n_353),
.SN(n_353)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_358),
.A2(n_362),
.B(n_363),
.Y(n_361)
);


endmodule