module real_jpeg_24541_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_0),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_0),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_0),
.B(n_60),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_0),
.B(n_49),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_0),
.B(n_37),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_0),
.B(n_30),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_0),
.B(n_57),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_1),
.B(n_93),
.Y(n_311)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_3),
.B(n_17),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_3),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_3),
.B(n_93),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_60),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_3),
.B(n_49),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_3),
.B(n_37),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_3),
.B(n_30),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_86),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_93),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_4),
.B(n_37),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_4),
.B(n_30),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_4),
.B(n_24),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_7),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_86),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_7),
.B(n_93),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_7),
.B(n_49),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_7),
.B(n_37),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_10),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_49),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_10),
.B(n_37),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_30),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_10),
.B(n_24),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_12),
.B(n_86),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_12),
.B(n_93),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_60),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_12),
.B(n_49),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_12),
.B(n_37),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_12),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_12),
.B(n_57),
.Y(n_324)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_14),
.B(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_14),
.B(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_14),
.B(n_60),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_14),
.B(n_49),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_14),
.B(n_37),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_14),
.B(n_57),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_30),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_15),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_15),
.B(n_86),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_93),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_15),
.B(n_60),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_15),
.B(n_49),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_15),
.B(n_37),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_16),
.B(n_60),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_16),
.B(n_49),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_16),
.B(n_37),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_16),
.B(n_30),
.Y(n_167)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_17),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_41),
.B2(n_42),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_27),
.B(n_103),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_36),
.C(n_40),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_28),
.A2(n_34),
.B1(n_36),
.B2(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_29),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_29),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_29),
.B(n_243),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_32),
.B(n_109),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_32),
.B(n_231),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_62),
.C(n_63),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_43),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.C(n_54),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_44),
.B(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_47),
.A2(n_48),
.B1(n_58),
.B2(n_338),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_55),
.C(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.C(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_51),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_53),
.B(n_54),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_55),
.A2(n_56),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_58),
.A2(n_310),
.B1(n_311),
.B2(n_338),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_58),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_SL g368 ( 
.A(n_58),
.B(n_311),
.C(n_336),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_59),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_59),
.B(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_62),
.B(n_63),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_381),
.C(n_383),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_375),
.C(n_376),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_357),
.C(n_358),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_328),
.C(n_329),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_303),
.C(n_304),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_271),
.C(n_272),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_236),
.C(n_237),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_201),
.C(n_202),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_171),
.C(n_172),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_150),
.C(n_151),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_132),
.C(n_133),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_110),
.C(n_111),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_95),
.C(n_100),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_90),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_91),
.C(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_88),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_86),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.C(n_105),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_109),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_123),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_116),
.C(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_122),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_130),
.C(n_131),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.C(n_141),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_139),
.C(n_140),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_149),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_165),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_166),
.C(n_170),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_160),
.C(n_161),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_159),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_161),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.CI(n_164),
.CON(n_161),
.SN(n_161)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.CI(n_169),
.CON(n_166),
.SN(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_187),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_176),
.C(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_183),
.C(n_186),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_178),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.CI(n_181),
.CON(n_178),
.SN(n_178)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_194),
.C(n_199),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_199),
.B2(n_200),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_192),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_193),
.B(n_226),
.C(n_227),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_197),
.C(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_222),
.B2(n_235),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_223),
.C(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_207),
.C(n_215),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_211),
.C(n_214),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_213),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_220),
.C(n_221),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_219),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_269),
.B2(n_270),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_260),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_260),
.C(n_269),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_250),
.C(n_251),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_245),
.C(n_247),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_259),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_256),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_255),
.B(n_278),
.C(n_281),
.Y(n_326)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_275),
.C(n_302),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_289),
.B2(n_302),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_284),
.C(n_285),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_281),
.A2(n_282),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_SL g342 ( 
.A(n_281),
.B(n_308),
.C(n_311),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_285),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.CI(n_288),
.CON(n_285),
.SN(n_285)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_301),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_297),
.C(n_299),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_297),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_298),
.A2(n_299),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_325),
.C(n_326),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_327),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_318),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_318),
.C(n_327),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_313),
.C(n_314),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_314),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.CI(n_317),
.CON(n_314),
.SN(n_314)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_324),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_332),
.C(n_344),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_343),
.B2(n_344),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_339),
.B2(n_340),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_341),
.C(n_342),
.Y(n_360)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_347),
.C(n_350),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_353),
.C(n_356),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_354),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_355),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_358)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_361),
.C(n_374),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_367),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_368),
.C(n_369),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_377),
.C(n_379),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_365),
.CI(n_366),
.CON(n_363),
.SN(n_363)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_370),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);


endmodule