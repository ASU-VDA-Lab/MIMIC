module real_jpeg_21944_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_0),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_32),
.B1(n_58),
.B2(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_0),
.A2(n_32),
.B1(n_50),
.B2(n_51),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_67),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_2),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_53),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_5),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_91),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_91),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_6),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_151),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_151),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_151),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_186)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_64),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_10),
.A2(n_47),
.B(n_50),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_155),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_10),
.A2(n_80),
.B1(n_141),
.B2(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_10),
.B(n_42),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_10),
.A2(n_30),
.B(n_243),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_157),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_157),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_157),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_13),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_127),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_127),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_127),
.Y(n_246)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_14),
.A2(n_30),
.A3(n_39),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_92),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.C(n_77),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_23),
.A2(n_24),
.B1(n_71),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_24)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_43),
.C(n_54),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_30),
.A2(n_31),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_30),
.B(n_62),
.Y(n_169)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_35),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_31),
.A2(n_63),
.B1(n_154),
.B2(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_31),
.B(n_155),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_33),
.A2(n_40),
.B1(n_42),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_33),
.A2(n_42),
.B1(n_74),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_33),
.A2(n_42),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_34),
.A2(n_37),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_34),
.A2(n_37),
.B1(n_152),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_34),
.A2(n_37),
.B1(n_181),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_34),
.A2(n_37),
.B1(n_123),
.B2(n_165),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_35),
.B(n_38),
.Y(n_238)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_39),
.A2(n_48),
.B(n_155),
.C(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_44),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_49),
.B1(n_76),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_45),
.A2(n_49),
.B1(n_87),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_45),
.A2(n_49),
.B1(n_120),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_45),
.A2(n_49),
.B1(n_143),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_45),
.A2(n_49),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_45),
.A2(n_49),
.B1(n_208),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_45),
.A2(n_49),
.B1(n_228),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_45),
.A2(n_49),
.B1(n_147),
.B2(n_246),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

CKINVDCx9p33_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_49),
.B(n_155),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_51),
.B(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_70),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_66),
.B2(n_68),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_61),
.B1(n_64),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_62),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_58),
.B(n_155),
.CON(n_154),
.SN(n_154)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_66),
.B1(n_68),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_60),
.A2(n_68),
.B1(n_90),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_60),
.A2(n_68),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_60),
.A2(n_68),
.B1(n_126),
.B2(n_163),
.Y(n_284)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_64),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_78),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_88),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_88),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_79),
.A2(n_86),
.B1(n_112),
.B2(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_84),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_118),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_80),
.A2(n_82),
.B1(n_140),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_80),
.A2(n_81),
.B1(n_171),
.B2(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_80),
.A2(n_82),
.B1(n_197),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_80),
.A2(n_141),
.B1(n_200),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_80),
.A2(n_82),
.B1(n_186),
.B2(n_230),
.Y(n_236)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_86),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_103),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_132),
.B(n_308),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_128),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_108),
.B(n_128),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_114),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_109),
.B(n_113),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_114),
.A2(n_115),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_124),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_116),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_117),
.B(n_119),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_121),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_302),
.B(n_307),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_289),
.B(n_301),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_187),
.B(n_271),
.C(n_288),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_172),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_136),
.B(n_172),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_158),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_138),
.B(n_144),
.C(n_158),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_139),
.B(n_142),
.Y(n_281)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_155),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_166),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_160),
.B(n_166),
.C(n_167),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_170),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_173),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_184),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_179),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_270),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_265),
.B(n_269),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_251),
.B(n_264),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_232),
.B(n_250),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_220),
.B(n_231),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_209),
.B(n_219),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_201),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_214),
.B(n_218),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_222),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_240),
.B1(n_248),
.B2(n_249),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_237),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_261),
.C(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_260),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_273),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_287),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_280),
.C(n_287),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_283),
.C(n_286),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_285),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_300),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_298),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_298),
.C(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);


endmodule