module fake_jpeg_4316_n_300 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx4_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_48),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_64),
.Y(n_71)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2x1_ASAP7_75t_SL g109 ( 
.A(n_54),
.B(n_35),
.Y(n_109)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_61),
.Y(n_86)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_72),
.Y(n_121)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_45),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_9),
.B(n_1),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_27),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_83),
.Y(n_124)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_88),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_27),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_84),
.B(n_6),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_47),
.B1(n_22),
.B2(n_35),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_28),
.B1(n_34),
.B2(n_36),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_89),
.A2(n_92),
.B1(n_7),
.B2(n_11),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_32),
.B1(n_37),
.B2(n_36),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_97),
.B1(n_99),
.B2(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_34),
.B1(n_30),
.B2(n_38),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_95),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_37),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_96),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_38),
.B1(n_19),
.B2(n_31),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_35),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_47),
.B1(n_33),
.B2(n_20),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_112),
.B1(n_143),
.B2(n_84),
.Y(n_157)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_119),
.Y(n_145)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_131),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_130),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_74),
.B(n_22),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_1),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_35),
.B(n_3),
.C(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_132),
.B(n_13),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_2),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_139),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_85),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_144),
.B1(n_71),
.B2(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_140),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_4),
.C(n_5),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_83),
.C(n_104),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_85),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_87),
.B1(n_98),
.B2(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_150),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_155),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_84),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_164),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_111),
.B1(n_125),
.B2(n_117),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_166),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_108),
.B1(n_88),
.B2(n_80),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_132),
.A2(n_90),
.B1(n_70),
.B2(n_86),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_78),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_81),
.A3(n_72),
.B1(n_79),
.B2(n_68),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_67),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_141),
.C(n_15),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_115),
.B1(n_130),
.B2(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_138),
.B1(n_114),
.B2(n_111),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_176),
.Y(n_205)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_81),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_113),
.B(n_100),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_133),
.C(n_136),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_197),
.C(n_202),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_155),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_134),
.B(n_129),
.C(n_139),
.D(n_112),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_172),
.A3(n_164),
.B1(n_167),
.B2(n_147),
.C1(n_171),
.C2(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_185),
.A2(n_172),
.B1(n_153),
.B2(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_188),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_114),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_161),
.B1(n_160),
.B2(n_146),
.Y(n_216)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_154),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_117),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_198),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_157),
.B1(n_162),
.B2(n_177),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_67),
.B(n_93),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_200),
.B(n_180),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_67),
.B1(n_16),
.B2(n_14),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_93),
.C(n_94),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_113),
.B(n_145),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_151),
.C(n_158),
.Y(n_202)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_149),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_218),
.B1(n_203),
.B2(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_206),
.Y(n_243)
);

AOI221xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_204),
.B1(n_182),
.B2(n_189),
.C(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_178),
.A2(n_172),
.B1(n_173),
.B2(n_169),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_196),
.B(n_194),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_181),
.C(n_179),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_192),
.B(n_205),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_228),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_205),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_229),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_239),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_200),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_241),
.Y(n_256)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_227),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_194),
.Y(n_236)
);

BUFx12_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_240),
.C(n_219),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_184),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_184),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_206),
.B(n_203),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_248),
.B1(n_212),
.B2(n_233),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_234),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_183),
.B1(n_199),
.B2(n_190),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_253),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_254),
.C(n_260),
.Y(n_265)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_259),
.B(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_228),
.C(n_215),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_266),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_248),
.B1(n_242),
.B2(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_246),
.C(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_229),
.B1(n_233),
.B2(n_216),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_269),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_210),
.C(n_209),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_213),
.C(n_231),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_279),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_250),
.B(n_255),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_277),
.B(n_255),
.Y(n_283)
);

AOI21x1_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_250),
.B(n_221),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_187),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_265),
.B1(n_256),
.B2(n_232),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_275),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_287),
.B1(n_245),
.B2(n_274),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_271),
.B1(n_270),
.B2(n_208),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_265),
.C(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_255),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_288),
.C(n_280),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_224),
.Y(n_292)
);

NOR4xp25_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_221),
.C(n_287),
.D(n_220),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_295),
.B1(n_199),
.B2(n_187),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_293),
.A3(n_291),
.B1(n_290),
.B2(n_211),
.C1(n_221),
.C2(n_183),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_187),
.Y(n_300)
);


endmodule