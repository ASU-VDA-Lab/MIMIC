module real_jpeg_2332_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_197;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_293;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_70;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_1),
.A2(n_47),
.B1(n_51),
.B2(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_1),
.A2(n_37),
.B1(n_39),
.B2(n_58),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_3),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_37),
.B1(n_39),
.B2(n_133),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_133),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_3),
.A2(n_47),
.B1(n_51),
.B2(n_133),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_4),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_37),
.B1(n_39),
.B2(n_158),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_158),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_4),
.A2(n_47),
.B1(n_51),
.B2(n_158),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_178),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_178),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_6),
.A2(n_47),
.B1(n_51),
.B2(n_178),
.Y(n_257)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_8),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_8),
.A2(n_41),
.B1(n_47),
.B2(n_51),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_37),
.B1(n_39),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_71),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_9),
.A2(n_47),
.B1(n_51),
.B2(n_71),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_12),
.B(n_26),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_12),
.B(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_12),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_12),
.A2(n_26),
.B(n_168),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_12),
.B(n_65),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g236 ( 
.A1(n_12),
.A2(n_39),
.B(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_12),
.B(n_47),
.C(n_50),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_204),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_12),
.B(n_87),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_12),
.B(n_45),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_37),
.B1(n_39),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_14),
.A2(n_47),
.B1(n_51),
.B2(n_62),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_15),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_15),
.A2(n_37),
.B1(n_39),
.B2(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_96),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_15),
.A2(n_47),
.B1(n_51),
.B2(n_96),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_16),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_16),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_16),
.A2(n_29),
.B1(n_47),
.B2(n_51),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_97),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_21),
.B(n_97),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_80),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_22),
.A2(n_73),
.B1(n_74),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_22),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_23),
.A2(n_24),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_44),
.C(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_25),
.A2(n_30),
.B1(n_36),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_27),
.A2(n_35),
.A3(n_39),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_30),
.A2(n_36),
.B1(n_40),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_30),
.A2(n_36),
.B1(n_95),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_30),
.A2(n_36),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_30),
.A2(n_36),
.B1(n_177),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_31),
.A2(n_132),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_33),
.B(n_37),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_36),
.Y(n_159)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_39),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_37),
.B(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_39),
.A2(n_55),
.A3(n_66),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_43)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_72),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_52),
.B(n_57),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_52),
.B1(n_57),
.B2(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_52),
.B1(n_79),
.B2(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_45),
.A2(n_52),
.B1(n_92),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_45),
.A2(n_52),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_45),
.A2(n_52),
.B1(n_200),
.B2(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_45),
.A2(n_52),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_45),
.A2(n_52),
.B1(n_227),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_46),
.A2(n_126),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_46),
.A2(n_151),
.B1(n_199),
.B2(n_239),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_47),
.B(n_255),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_52),
.Y(n_151)
);

AO22x2_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_54),
.B(n_67),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_55),
.B(n_245),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_69),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_63),
.A2(n_65),
.B1(n_129),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_70),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_64),
.A2(n_77),
.B1(n_104),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_64),
.A2(n_104),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_64),
.A2(n_104),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_64),
.A2(n_104),
.B1(n_174),
.B2(n_190),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_64),
.A2(n_104),
.B1(n_189),
.B2(n_236),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_80),
.B(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_93),
.B(n_94),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_82),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_83),
.A2(n_93),
.B1(n_94),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_83),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_88),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_84),
.A2(n_86),
.B1(n_122),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_84),
.A2(n_86),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_84),
.A2(n_86),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_85),
.A2(n_87),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_85),
.A2(n_87),
.B1(n_171),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_85),
.A2(n_87),
.B1(n_208),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_85),
.A2(n_87),
.B1(n_204),
.B2(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_85),
.A2(n_87),
.B1(n_257),
.B2(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_294),
.B(n_299),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_160),
.B(n_293),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_142),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_115),
.B(n_142),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_134),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_116),
.B(n_136),
.C(n_141),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.C(n_130),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_118),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_130),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_141),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_147),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.C(n_156),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_149),
.B(n_152),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_156),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_183),
.B(n_292),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_181),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_162),
.B(n_181),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_180),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_163),
.B(n_180),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_165),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.C(n_176),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_166),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_170),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_173),
.B(n_176),
.Y(n_283)
);

AOI31xp33_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_277),
.A3(n_286),
.B(n_289),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_222),
.B(n_276),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_210),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_186),
.B(n_210),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.C(n_201),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_187),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_192),
.C(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_197),
.B(n_201),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_210),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_210),
.B(n_287),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.CI(n_213),
.CON(n_210),
.SN(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_214),
.B(n_217),
.C(n_221),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_271),
.B(n_275),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_240),
.B(n_270),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_232),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_229),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_235),
.C(n_238),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_251),
.B(n_269),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_263),
.B(n_268),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_258),
.B(n_262),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_267),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_281),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_298),
.Y(n_299)
);


endmodule