module fake_aes_10277_n_656 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_656);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_656;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_65), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_20), .Y(n_79) );
NOR2xp67_ASAP7_75t_L g80 ( .A(n_2), .B(n_38), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_32), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_59), .Y(n_82) );
CKINVDCx14_ASAP7_75t_R g83 ( .A(n_31), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_54), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_71), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_41), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_61), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_28), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_48), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_55), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_36), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_26), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_58), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_21), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_4), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_35), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_27), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_43), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_52), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_74), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_24), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_49), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_12), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_5), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_5), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_63), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_25), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_45), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_4), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_102), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_108), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_102), .B(n_0), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_105), .B(n_1), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_102), .B(n_3), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_78), .A2(n_37), .B(n_76), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
CKINVDCx8_ASAP7_75t_R g131 ( .A(n_91), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_113), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_82), .A2(n_90), .B(n_97), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
BUFx8_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_107), .B(n_33), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_113), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_79), .A2(n_3), .B1(n_6), .B2(n_7), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_90), .A2(n_40), .B(n_75), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_79), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
NOR2x1_ASAP7_75t_L g146 ( .A(n_80), .B(n_6), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_99), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g148 ( .A1(n_119), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_148) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_81), .A2(n_44), .B(n_73), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_103), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_87), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_88), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_99), .B(n_14), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_138), .B(n_110), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
BUFx8_ASAP7_75t_SL g158 ( .A(n_138), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_127), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_123), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
OR2x2_ASAP7_75t_L g165 ( .A(n_143), .B(n_119), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_129), .B(n_83), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_129), .B(n_107), .Y(n_170) );
INVxp33_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
INVx1_ASAP7_75t_SL g172 ( .A(n_125), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_131), .B(n_101), .Y(n_173) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_155), .B(n_117), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_131), .B(n_95), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_130), .B(n_81), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_130), .B(n_85), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
NAND2xp33_ASAP7_75t_L g179 ( .A(n_137), .B(n_86), .Y(n_179) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_155), .B(n_117), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_135), .B(n_112), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_127), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_135), .B(n_98), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_136), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_155), .A2(n_134), .B1(n_139), .B2(n_144), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_139), .B(n_115), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_144), .B(n_114), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_145), .B(n_96), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_145), .B(n_104), .Y(n_193) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_136), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_155), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_147), .B(n_104), .Y(n_196) );
NAND3xp33_ASAP7_75t_L g197 ( .A(n_134), .B(n_94), .C(n_116), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_147), .B(n_116), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_197), .A2(n_149), .B(n_134), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_169), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_168), .B(n_134), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_190), .B(n_100), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_184), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_174), .A2(n_154), .B1(n_152), .B2(n_140), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g209 ( .A1(n_172), .A2(n_140), .B1(n_154), .B2(n_152), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_190), .B(n_126), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_174), .A2(n_121), .B1(n_150), .B2(n_148), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_190), .B(n_186), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_186), .B(n_136), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_188), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_156), .B(n_171), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_174), .B(n_137), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_177), .B(n_147), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_180), .A2(n_137), .B1(n_111), .B2(n_103), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_181), .B(n_147), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_189), .B(n_146), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_188), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_165), .B(n_121), .Y(n_224) );
NAND3xp33_ASAP7_75t_SL g225 ( .A(n_165), .B(n_106), .C(n_111), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g226 ( .A1(n_162), .A2(n_97), .B(n_94), .C(n_118), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_191), .B(n_146), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_180), .A2(n_137), .B1(n_109), .B2(n_118), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_180), .A2(n_109), .B1(n_137), .B2(n_149), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_195), .B(n_162), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_183), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_161), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_185), .B(n_142), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_195), .B(n_128), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_163), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_164), .B(n_137), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_164), .B(n_137), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_164), .B(n_128), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_194), .B(n_93), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_164), .B(n_166), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_161), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_166), .B(n_128), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_158), .Y(n_243) );
AND3x1_ASAP7_75t_L g244 ( .A(n_198), .B(n_153), .C(n_141), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_166), .B(n_128), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_166), .B(n_142), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_163), .Y(n_247) );
BUFx12f_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_178), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_193), .A2(n_142), .B1(n_93), .B2(n_153), .Y(n_250) );
NAND2xp33_ASAP7_75t_L g251 ( .A(n_183), .B(n_151), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_225), .B(n_179), .Y(n_252) );
BUFx12f_ASAP7_75t_L g253 ( .A(n_224), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_248), .Y(n_254) );
AND2x6_ASAP7_75t_L g255 ( .A(n_234), .B(n_159), .Y(n_255) );
OAI22xp5_ASAP7_75t_SL g256 ( .A1(n_209), .A2(n_187), .B1(n_142), .B2(n_196), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_199), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_215), .B(n_192), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_175), .B1(n_173), .B2(n_170), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_230), .B(n_160), .Y(n_260) );
NAND3xp33_ASAP7_75t_SL g261 ( .A(n_211), .B(n_176), .C(n_157), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_240), .B(n_160), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_240), .B(n_159), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_200), .A2(n_157), .B(n_197), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_240), .B(n_183), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_240), .B(n_183), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_224), .B(n_15), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_221), .B(n_183), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_227), .B(n_16), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_208), .A2(n_182), .B(n_178), .C(n_153), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_223), .B(n_182), .Y(n_271) );
NOR3xp33_ASAP7_75t_L g272 ( .A(n_209), .B(n_141), .C(n_18), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_245), .B(n_242), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_223), .Y(n_274) );
CKINVDCx8_ASAP7_75t_R g275 ( .A(n_243), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_211), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g277 ( .A1(n_203), .A2(n_141), .B(n_151), .Y(n_277) );
OAI21xp33_ASAP7_75t_L g278 ( .A1(n_218), .A2(n_151), .B(n_133), .Y(n_278) );
BUFx12f_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_246), .A2(n_151), .B(n_133), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_235), .A2(n_151), .B1(n_133), .B2(n_124), .Y(n_282) );
BUFx4f_ASAP7_75t_L g283 ( .A(n_248), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_235), .B(n_17), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_247), .B(n_17), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_223), .Y(n_287) );
NOR3xp33_ASAP7_75t_SL g288 ( .A(n_204), .B(n_18), .C(n_19), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_201), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_220), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_247), .A2(n_151), .B(n_133), .C(n_124), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_220), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_201), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_217), .B(n_19), .Y(n_294) );
AOI22xp33_ASAP7_75t_SL g295 ( .A1(n_216), .A2(n_133), .B1(n_124), .B2(n_122), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_205), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_216), .A2(n_133), .B1(n_124), .B2(n_122), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_229), .B(n_124), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_259), .B(n_220), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_267), .B(n_219), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_SL g301 ( .A1(n_298), .A2(n_229), .B(n_250), .C(n_233), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
AO31x2_ASAP7_75t_L g303 ( .A1(n_273), .A2(n_202), .A3(n_206), .B(n_207), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_276), .B(n_228), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_270), .A2(n_226), .B(n_234), .C(n_206), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_261), .A2(n_210), .B(n_222), .C(n_207), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_280), .A2(n_200), .B(n_250), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_268), .A2(n_236), .B(n_237), .Y(n_308) );
AO31x2_ASAP7_75t_L g309 ( .A1(n_291), .A2(n_222), .A3(n_214), .B(n_205), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_298), .A2(n_213), .B(n_212), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_SL g311 ( .A1(n_291), .A2(n_239), .B(n_214), .C(n_241), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_253), .A2(n_244), .B1(n_249), .B2(n_232), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_272), .A2(n_249), .B(n_241), .C(n_232), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_256), .B1(n_281), .B2(n_255), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_286), .A2(n_244), .B(n_251), .C(n_124), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_279), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_269), .A2(n_122), .B(n_23), .C(n_29), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_253), .A2(n_231), .B1(n_122), .B2(n_42), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_294), .A2(n_122), .B(n_231), .C(n_46), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_263), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_279), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_258), .B(n_122), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_SL g324 ( .A1(n_257), .A2(n_22), .B(n_30), .C(n_47), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_287), .B(n_231), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_257), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_285), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_260), .A2(n_231), .B(n_51), .C(n_53), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_287), .B(n_231), .Y(n_330) );
AOI221xp5_ASAP7_75t_SL g331 ( .A1(n_278), .A2(n_50), .B1(n_56), .B2(n_60), .C(n_62), .Y(n_331) );
OAI21xp33_ASAP7_75t_L g332 ( .A1(n_314), .A2(n_252), .B(n_288), .Y(n_332) );
OA21x2_ASAP7_75t_L g333 ( .A1(n_331), .A2(n_277), .B(n_264), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_307), .A2(n_297), .B(n_282), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_304), .A2(n_252), .B1(n_255), .B2(n_292), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_326), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_320), .B(n_296), .Y(n_337) );
AND2x4_ASAP7_75t_SL g338 ( .A(n_316), .B(n_254), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_327), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_328), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_301), .A2(n_296), .B(n_293), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_314), .A2(n_293), .B1(n_289), .B2(n_295), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_305), .A2(n_289), .B(n_255), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_317), .A2(n_282), .B(n_271), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_299), .A2(n_290), .B1(n_292), .B2(n_274), .C(n_283), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_300), .A2(n_275), .B1(n_283), .B2(n_254), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_313), .B(n_254), .Y(n_350) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_315), .A2(n_266), .A3(n_255), .B(n_271), .Y(n_351) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_299), .A2(n_274), .B(n_290), .C(n_265), .Y(n_352) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_301), .A2(n_265), .B(n_255), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_308), .A2(n_254), .B(n_67), .Y(n_354) );
BUFx12f_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_64), .B(n_68), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_303), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_344), .B(n_302), .Y(n_359) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_341), .A2(n_329), .B(n_311), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_332), .A2(n_321), .B1(n_312), .B2(n_316), .Y(n_361) );
OA21x2_ASAP7_75t_L g362 ( .A1(n_344), .A2(n_310), .B(n_318), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_357), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_355), .Y(n_365) );
AOI21xp5_ASAP7_75t_SL g366 ( .A1(n_342), .A2(n_306), .B(n_330), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_357), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
OAI322xp33_ASAP7_75t_L g369 ( .A1(n_348), .A2(n_70), .A3(n_77), .B1(n_309), .B2(n_322), .C1(n_324), .C2(n_346), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_337), .A2(n_322), .B1(n_309), .B2(n_324), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_357), .A2(n_309), .B(n_334), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_346), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_349), .B(n_309), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_349), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_342), .B1(n_347), .B2(n_337), .C(n_335), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_336), .B(n_340), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_343), .A2(n_334), .B(n_345), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_338), .B(n_355), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_355), .B1(n_358), .B2(n_353), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_339), .B(n_340), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_339), .B(n_358), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_343), .A2(n_350), .B1(n_352), .B2(n_338), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_351), .B(n_353), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_353), .B(n_351), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_351), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_372), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_387), .B(n_351), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_374), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_387), .B(n_351), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_364), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_387), .B(n_351), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_379), .A2(n_350), .B1(n_356), .B2(n_333), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_374), .B(n_350), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_373), .B(n_350), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_367), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_367), .B(n_333), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_370), .A2(n_354), .B(n_345), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_388), .B(n_333), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_388), .B(n_333), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_380), .B(n_356), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_363), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_373), .B(n_350), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_380), .B(n_356), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_373), .B(n_356), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_359), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_359), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
INVx4_ASAP7_75t_L g423 ( .A(n_363), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_384), .B(n_386), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_359), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_386), .B(n_381), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_382), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_376), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_371), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_390), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_427), .B(n_386), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_427), .B(n_384), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
NOR3xp33_ASAP7_75t_SL g436 ( .A(n_401), .B(n_378), .C(n_369), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_419), .B(n_381), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_427), .B(n_371), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_419), .B(n_381), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_429), .B(n_371), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_429), .B(n_379), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_428), .B(n_377), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_389), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_394), .B(n_377), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_390), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_394), .B(n_377), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_394), .B(n_377), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_396), .B(n_377), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_396), .B(n_362), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_397), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_390), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_396), .B(n_362), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_428), .B(n_365), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_405), .B(n_365), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_398), .B(n_362), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_424), .B(n_360), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_391), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_400), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_397), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_420), .B(n_375), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_391), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_420), .B(n_361), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_400), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_393), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_416), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_398), .B(n_362), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_405), .B(n_385), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g476 ( .A(n_401), .B(n_375), .C(n_361), .D(n_366), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_398), .B(n_362), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_392), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_393), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_405), .B(n_385), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_425), .B(n_430), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_416), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_392), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_370), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_424), .B(n_360), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_421), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_424), .B(n_360), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_437), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_440), .B(n_424), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_433), .B(n_425), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
AOI21xp5_ASAP7_75t_SL g493 ( .A1(n_483), .A2(n_423), .B(n_392), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_470), .B(n_430), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_468), .B(n_426), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_468), .B(n_426), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_432), .Y(n_499) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_447), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_476), .A2(n_423), .B1(n_415), .B2(n_414), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_433), .B(n_395), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_435), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_481), .B(n_395), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_478), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_434), .B(n_415), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_435), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_481), .B(n_399), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_434), .B(n_415), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_462), .B(n_399), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_438), .B(n_418), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_440), .B(n_402), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_462), .B(n_402), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_472), .B(n_402), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_461), .B(n_411), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_438), .B(n_418), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_411), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_442), .B(n_406), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_450), .B(n_414), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_478), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_442), .B(n_418), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_439), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_439), .B(n_406), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_450), .B(n_412), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_458), .B(n_423), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_441), .B(n_410), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_476), .B(n_423), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_452), .B(n_421), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_441), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_443), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_452), .B(n_421), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_467), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_451), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_443), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_449), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_453), .B(n_422), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_453), .B(n_422), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_451), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_451), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_454), .B(n_412), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_454), .B(n_410), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_449), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_422), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_475), .B(n_423), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_455), .B(n_412), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_495), .B(n_445), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_490), .B(n_459), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_502), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_493), .A2(n_436), .B(n_445), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_490), .B(n_463), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_491), .B(n_463), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_527), .A2(n_484), .B1(n_459), .B2(n_477), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_497), .B(n_498), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_524), .B(n_455), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_527), .A2(n_436), .B(n_414), .C(n_484), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_524), .B(n_474), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_540), .B(n_474), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_540), .B(n_477), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_529), .Y(n_562) );
AO21x1_ASAP7_75t_L g563 ( .A1(n_500), .A2(n_479), .B(n_469), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_545), .B(n_446), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_530), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_545), .B(n_446), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_501), .A2(n_414), .B(n_480), .C(n_456), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_534), .Y(n_568) );
OAI21xp33_ASAP7_75t_SL g569 ( .A1(n_493), .A2(n_448), .B(n_456), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_535), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_512), .B(n_488), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_544), .A2(n_480), .B1(n_448), .B2(n_444), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_512), .B(n_488), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_542), .Y(n_574) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_519), .B(n_460), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_541), .B(n_444), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_525), .A2(n_509), .B1(n_506), .B2(n_511), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_518), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_496), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_500), .Y(n_581) );
AOI21xp33_ASAP7_75t_SL g582 ( .A1(n_525), .A2(n_479), .B(n_469), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_512), .B(n_486), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_505), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_532), .B(n_464), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_489), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_515), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_569), .A2(n_532), .B(n_520), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_554), .B(n_526), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_546), .B(n_510), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_579), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_580), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_552), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_558), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_575), .A2(n_486), .B1(n_516), .B2(n_521), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_549), .A2(n_464), .B1(n_513), .B2(n_514), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_546), .B(n_517), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_556), .A2(n_528), .B(n_531), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_560), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_562), .Y(n_601) );
OAI311xp33_ASAP7_75t_L g602 ( .A1(n_556), .A2(n_543), .A3(n_508), .B1(n_504), .C1(n_523), .Y(n_602) );
NAND3x2_ASAP7_75t_L g603 ( .A(n_576), .B(n_537), .C(n_536), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_567), .B(n_369), .C(n_465), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_584), .B(n_460), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_565), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_575), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_567), .A2(n_464), .B(n_465), .C(n_494), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_586), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_554), .B(n_539), .Y(n_610) );
OAI32xp33_ASAP7_75t_L g611 ( .A1(n_577), .A2(n_458), .A3(n_538), .B1(n_533), .B2(n_499), .Y(n_611) );
OAI22xp33_ASAP7_75t_SL g612 ( .A1(n_581), .A2(n_464), .B1(n_458), .B2(n_533), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_571), .B(n_539), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_563), .B(n_458), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g615 ( .A1(n_605), .A2(n_572), .A3(n_585), .B1(n_561), .B2(n_587), .Y(n_615) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_589), .A2(n_553), .B(n_559), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_602), .A2(n_572), .B1(n_548), .B2(n_578), .C(n_588), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_590), .B(n_581), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_599), .A2(n_566), .B(n_564), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_592), .B(n_568), .Y(n_620) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_607), .A2(n_585), .B(n_555), .Y(n_621) );
OAI21xp33_ASAP7_75t_SL g622 ( .A1(n_614), .A2(n_557), .B(n_547), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
AOI22xp5_ASAP7_75t_SL g624 ( .A1(n_612), .A2(n_585), .B1(n_550), .B2(n_551), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_614), .A2(n_582), .B(n_570), .Y(n_625) );
OAI322xp33_ASAP7_75t_SL g626 ( .A1(n_598), .A2(n_574), .A3(n_492), .B1(n_538), .B2(n_499), .C1(n_494), .C2(n_473), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_595), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_597), .A2(n_583), .B1(n_573), .B2(n_492), .C(n_466), .Y(n_628) );
AO22x1_ASAP7_75t_L g629 ( .A1(n_604), .A2(n_417), .B1(n_413), .B2(n_487), .Y(n_629) );
OAI31xp33_ASAP7_75t_L g630 ( .A1(n_608), .A2(n_417), .A3(n_413), .B(n_410), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g631 ( .A1(n_616), .A2(n_609), .B1(n_597), .B2(n_590), .C1(n_610), .C2(n_611), .Y(n_631) );
OAI221xp5_ASAP7_75t_SL g632 ( .A1(n_615), .A2(n_596), .B1(n_610), .B2(n_591), .C(n_603), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_SL g633 ( .A1(n_630), .A2(n_628), .B(n_625), .C(n_627), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_626), .A2(n_606), .B1(n_601), .B2(n_600), .C(n_593), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_622), .B(n_613), .Y(n_635) );
NOR2xp33_ASAP7_75t_R g636 ( .A(n_618), .B(n_417), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_624), .B(n_431), .C(n_487), .Y(n_637) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_623), .A2(n_466), .B1(n_485), .B2(n_482), .C1(n_473), .C2(n_471), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_620), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_631), .A2(n_621), .B(n_617), .C(n_619), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_632), .A2(n_629), .B1(n_620), .B2(n_471), .C(n_473), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_633), .A2(n_409), .B(n_413), .C(n_431), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_637), .A2(n_466), .B1(n_485), .B2(n_482), .C(n_471), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_635), .A2(n_457), .B1(n_485), .B2(n_482), .C(n_487), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_640), .B(n_639), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_642), .Y(n_646) );
NOR3xp33_ASAP7_75t_SL g647 ( .A(n_641), .B(n_638), .C(n_634), .Y(n_647) );
OR3x2_ASAP7_75t_L g648 ( .A(n_646), .B(n_644), .C(n_636), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_645), .B(n_457), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_649), .Y(n_650) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_648), .A2(n_643), .B(n_647), .Y(n_651) );
NOR2x1p5_ASAP7_75t_L g652 ( .A(n_651), .B(n_431), .Y(n_652) );
AOI21xp33_ASAP7_75t_SL g653 ( .A1(n_652), .A2(n_651), .B(n_650), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_457), .B1(n_408), .B2(n_409), .Y(n_654) );
AO221x2_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_360), .B1(n_408), .B2(n_409), .C(n_645), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_409), .B(n_408), .Y(n_656) );
endmodule