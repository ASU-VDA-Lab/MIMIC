module fake_jpeg_4280_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_60),
.Y(n_93)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_22),
.B1(n_28),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_19),
.B1(n_17),
.B2(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_82),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_95),
.B1(n_50),
.B2(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_84),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_41),
.C(n_27),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_31),
.C(n_48),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_31),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_20),
.B(n_24),
.C(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_54),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_24),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_31),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_84),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_21),
.B1(n_12),
.B2(n_11),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_59),
.B1(n_56),
.B2(n_15),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_31),
.B1(n_48),
.B2(n_32),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_71),
.B1(n_67),
.B2(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_110),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_66),
.B1(n_51),
.B2(n_55),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_101),
.Y(n_137)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_51),
.B1(n_55),
.B2(n_58),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_61),
.B1(n_45),
.B2(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_61),
.B1(n_45),
.B2(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_118),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_17),
.B1(n_19),
.B2(n_41),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_19),
.B1(n_68),
.B2(n_32),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_90),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_95),
.B(n_85),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_127),
.B(n_148),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_95),
.B1(n_118),
.B2(n_109),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_123),
.A2(n_114),
.B1(n_91),
.B2(n_86),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_95),
.B(n_90),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_98),
.B(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_147),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g136 ( 
.A(n_101),
.Y(n_136)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_90),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_146),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_94),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_117),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_76),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_112),
.C(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_72),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_82),
.B(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_100),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_168),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_160),
.C(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_159),
.Y(n_191)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_162),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_148),
.B(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_96),
.C(n_112),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_96),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_166),
.C(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_110),
.C(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_111),
.B(n_77),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_77),
.C(n_54),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_143),
.C(n_126),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_176),
.B1(n_123),
.B2(n_132),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_134),
.B1(n_138),
.B2(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_178),
.A2(n_194),
.B1(n_155),
.B2(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_138),
.B1(n_123),
.B2(n_122),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_188),
.B1(n_203),
.B2(n_162),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_0),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_123),
.B1(n_127),
.B2(n_132),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_14),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_130),
.C(n_133),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_199),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_142),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_195),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_123),
.B1(n_129),
.B2(n_133),
.Y(n_194)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_129),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_135),
.B(n_148),
.C(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_125),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_125),
.C(n_141),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_74),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_180),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_161),
.A2(n_114),
.B1(n_91),
.B2(n_86),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_158),
.B1(n_173),
.B2(n_177),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_216),
.B(n_218),
.C(n_228),
.Y(n_230)
);

NOR4xp25_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_151),
.C(n_165),
.D(n_153),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_222),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_157),
.B1(n_168),
.B2(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_170),
.B(n_171),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_212),
.A2(n_227),
.B(n_0),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_86),
.B1(n_150),
.B2(n_62),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_150),
.B1(n_74),
.B2(n_79),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_88),
.B1(n_79),
.B2(n_62),
.Y(n_224)
);

NAND4xp25_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_62),
.C(n_193),
.D(n_88),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_32),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_192),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_232),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_202),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_181),
.C(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_235),
.C(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_181),
.C(n_187),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_245),
.B1(n_210),
.B2(n_221),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_190),
.C(n_180),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_32),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_32),
.C(n_16),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_79),
.C(n_1),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_79),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_242),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_244),
.A2(n_215),
.B1(n_217),
.B2(n_223),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_254),
.B1(n_255),
.B2(n_259),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_236),
.A2(n_217),
.B1(n_224),
.B2(n_213),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_230),
.B1(n_233),
.B2(n_246),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_218),
.B1(n_204),
.B2(n_214),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_226),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_239),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_265),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_243),
.B1(n_230),
.B2(n_241),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_235),
.C(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_266),
.C(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_216),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_253),
.C(n_257),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_256),
.B(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_275),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_273),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_247),
.C(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_13),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_2),
.C(n_3),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_4),
.B(n_5),
.Y(n_276)
);

AOI21x1_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_7),
.B(n_8),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_275),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

AND2x4_ASAP7_75t_SL g281 ( 
.A(n_278),
.B(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_283),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_281),
.A2(n_270),
.B(n_277),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_9),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_289),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_288),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_10),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_9),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_296),
.A2(n_297),
.B(n_292),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_293),
.C(n_294),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);


endmodule