module real_aes_6183_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_726, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_726;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_713;
wire n_147;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g467 ( .A1(n_0), .A2(n_205), .B(n_468), .C(n_471), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_1), .B(n_462), .Y(n_472) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_2), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g240 ( .A(n_3), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_4), .B(n_157), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_5), .A2(n_457), .B(n_545), .Y(n_544) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_6), .A2(n_180), .B(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_7), .A2(n_38), .B1(n_150), .B2(n_174), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_8), .B(n_180), .Y(n_252) );
AND2x6_ASAP7_75t_L g165 ( .A(n_9), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_10), .A2(n_165), .B(n_448), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_11), .B(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_11), .B(n_39), .Y(n_127) );
INVx1_ASAP7_75t_L g146 ( .A(n_12), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_13), .B(n_155), .Y(n_188) );
INVx1_ASAP7_75t_L g232 ( .A(n_14), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_15), .A2(n_75), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_15), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_16), .B(n_157), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_17), .B(n_181), .Y(n_219) );
AO32x2_ASAP7_75t_L g202 ( .A1(n_18), .A2(n_179), .A3(n_180), .B1(n_203), .B2(n_207), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_19), .B(n_150), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_20), .B(n_181), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_21), .A2(n_55), .B1(n_150), .B2(n_174), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g177 ( .A1(n_22), .A2(n_82), .B1(n_150), .B2(n_155), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_23), .B(n_150), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_24), .A2(n_179), .B(n_448), .C(n_495), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_25), .A2(n_179), .B(n_448), .C(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_26), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_27), .B(n_142), .Y(n_261) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_28), .A2(n_93), .B1(n_703), .B2(n_704), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_28), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_29), .A2(n_701), .B1(n_702), .B2(n_705), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_29), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_30), .A2(n_457), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_31), .B(n_142), .Y(n_167) );
INVx2_ASAP7_75t_L g152 ( .A(n_32), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_33), .A2(n_454), .B(n_480), .C(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_34), .B(n_150), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_35), .B(n_142), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_36), .A2(n_43), .B1(n_438), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_36), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_37), .B(n_190), .Y(n_511) );
INVx1_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_40), .B(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_41), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_42), .B(n_157), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_43), .A2(n_133), .B1(n_438), .B2(n_439), .Y(n_132) );
INVx1_ASAP7_75t_L g438 ( .A(n_43), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_44), .B(n_457), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_45), .A2(n_454), .B(n_480), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_46), .B(n_150), .Y(n_247) );
INVx1_ASAP7_75t_L g469 ( .A(n_47), .Y(n_469) );
AOI22xp5_ASAP7_75t_SL g129 ( .A1(n_48), .A2(n_124), .B1(n_130), .B2(n_708), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_49), .A2(n_91), .B1(n_174), .B2(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g532 ( .A(n_50), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_51), .B(n_150), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_52), .B(n_150), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_53), .B(n_457), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_54), .B(n_238), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g223 ( .A1(n_56), .A2(n_60), .B1(n_150), .B2(n_155), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_57), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_58), .B(n_150), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_59), .B(n_150), .Y(n_260) );
INVx1_ASAP7_75t_L g166 ( .A(n_61), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_62), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_63), .B(n_462), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_64), .A2(n_235), .B(n_238), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_65), .B(n_150), .Y(n_241) );
INVx1_ASAP7_75t_L g145 ( .A(n_66), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_68), .B(n_157), .Y(n_485) );
AO32x2_ASAP7_75t_L g171 ( .A1(n_69), .A2(n_172), .A3(n_178), .B1(n_179), .B2(n_180), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_70), .B(n_158), .Y(n_522) );
INVx1_ASAP7_75t_L g259 ( .A(n_71), .Y(n_259) );
INVx1_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_73), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_74), .B(n_484), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_75), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_76), .A2(n_448), .B(n_450), .C(n_454), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_77), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_78), .B(n_155), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_79), .Y(n_546) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_81), .B(n_483), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_83), .B(n_174), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_84), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_85), .B(n_155), .Y(n_162) );
INVx2_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_87), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_88), .B(n_176), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_89), .B(n_155), .Y(n_248) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
OR2x2_ASAP7_75t_L g123 ( .A(n_90), .B(n_124), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_92), .A2(n_103), .B1(n_155), .B2(n_156), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_93), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_94), .B(n_457), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_95), .Y(n_482) );
INVxp67_ASAP7_75t_L g549 ( .A(n_96), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_97), .B(n_155), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_98), .A2(n_105), .B1(n_116), .B2(n_723), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g451 ( .A(n_100), .Y(n_451) );
INVx1_ASAP7_75t_L g518 ( .A(n_101), .Y(n_518) );
AND2x2_ASAP7_75t_L g534 ( .A(n_102), .B(n_142), .Y(n_534) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g724 ( .A(n_108), .Y(n_724) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AO22x2_ASAP7_75t_SL g131 ( .A1(n_112), .A2(n_132), .B1(n_440), .B2(n_699), .Y(n_131) );
INVx1_ASAP7_75t_L g699 ( .A(n_112), .Y(n_699) );
NOR2x2_ASAP7_75t_L g710 ( .A(n_112), .B(n_124), .Y(n_710) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AOI22x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_129), .B1(n_711), .B2(n_712), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g711 ( .A(n_119), .Y(n_711) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_121), .A2(n_713), .B(n_722), .Y(n_712) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_128), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g722 ( .A(n_123), .Y(n_722) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI22xp33_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_700), .B1(n_706), .B2(n_707), .Y(n_130) );
INVx1_ASAP7_75t_L g706 ( .A(n_131), .Y(n_706) );
INVx1_ASAP7_75t_L g439 ( .A(n_133), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_133), .A2(n_439), .B1(n_719), .B2(n_720), .Y(n_718) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_359), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_308), .C(n_350), .Y(n_134) );
AOI211xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_213), .B(n_262), .C(n_284), .Y(n_135) );
OAI211xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_168), .B(n_196), .C(n_208), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_138), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g371 ( .A(n_138), .B(n_288), .Y(n_371) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g273 ( .A(n_139), .B(n_199), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_139), .B(n_184), .Y(n_390) );
INVx1_ASAP7_75t_L g408 ( .A(n_139), .Y(n_408) );
AND2x2_ASAP7_75t_L g417 ( .A(n_139), .B(n_305), .Y(n_417) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g300 ( .A(n_140), .B(n_184), .Y(n_300) );
AND2x2_ASAP7_75t_L g358 ( .A(n_140), .B(n_305), .Y(n_358) );
INVx1_ASAP7_75t_L g402 ( .A(n_140), .Y(n_402) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g279 ( .A(n_141), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g287 ( .A(n_141), .Y(n_287) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_141), .Y(n_327) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_167), .Y(n_141) );
INVx2_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_142), .A2(n_185), .B(n_195), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_142), .A2(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g501 ( .A(n_142), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_142), .A2(n_529), .B(n_530), .Y(n_528) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_L g181 ( .A(n_143), .B(n_144), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_160), .B(n_165), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_153), .B(n_154), .C(n_157), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_150), .Y(n_453) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
AND2x6_ASAP7_75t_L g448 ( .A(n_151), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g156 ( .A(n_152), .Y(n_156) );
INVx1_ASAP7_75t_L g239 ( .A(n_152), .Y(n_239) );
INVx2_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_157), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_157), .A2(n_256), .B(n_257), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_157), .B(n_549), .Y(n_548) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g172 ( .A1(n_158), .A2(n_173), .B1(n_176), .B2(n_177), .Y(n_172) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_159), .Y(n_164) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
INVx1_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
INVx1_ASAP7_75t_L g449 ( .A(n_159), .Y(n_449) );
AND2x2_ASAP7_75t_L g458 ( .A(n_159), .B(n_239), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g235 ( .A(n_163), .Y(n_235) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g484 ( .A(n_164), .Y(n_484) );
BUFx3_ASAP7_75t_L g179 ( .A(n_165), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_165), .A2(n_186), .B(n_191), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_165), .A2(n_231), .B(n_236), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_165), .A2(n_246), .B(n_249), .Y(n_245) );
INVx4_ASAP7_75t_SL g455 ( .A(n_165), .Y(n_455) );
AND2x4_ASAP7_75t_L g457 ( .A(n_165), .B(n_458), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_165), .B(n_458), .Y(n_519) );
INVxp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
AND2x2_ASAP7_75t_L g266 ( .A(n_170), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g299 ( .A(n_170), .Y(n_299) );
OR2x2_ASAP7_75t_L g425 ( .A(n_170), .B(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_170), .B(n_184), .Y(n_429) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
INVx1_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
AND2x2_ASAP7_75t_L g288 ( .A(n_171), .B(n_201), .Y(n_288) );
AND2x2_ASAP7_75t_L g328 ( .A(n_171), .B(n_202), .Y(n_328) );
INVx2_ASAP7_75t_L g471 ( .A(n_175), .Y(n_471) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_175), .Y(n_486) );
INVx2_ASAP7_75t_L g194 ( .A(n_176), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_176), .A2(n_204), .B1(n_205), .B2(n_206), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_176), .A2(n_205), .B1(n_222), .B2(n_223), .Y(n_221) );
INVx4_ASAP7_75t_L g470 ( .A(n_176), .Y(n_470) );
INVx1_ASAP7_75t_L g498 ( .A(n_178), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g220 ( .A(n_179), .B(n_221), .C(n_224), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_179), .A2(n_255), .B(n_258), .Y(n_254) );
INVx4_ASAP7_75t_L g224 ( .A(n_180), .Y(n_224) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_180), .A2(n_245), .B(n_252), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_180), .A2(n_508), .B(n_509), .Y(n_507) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_180), .Y(n_543) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g207 ( .A(n_181), .Y(n_207) );
INVxp67_ASAP7_75t_L g370 ( .A(n_182), .Y(n_370) );
AND2x4_ASAP7_75t_L g395 ( .A(n_182), .B(n_288), .Y(n_395) );
BUFx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_SL g286 ( .A(n_183), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g200 ( .A(n_184), .B(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g274 ( .A(n_184), .B(n_202), .Y(n_274) );
INVx1_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
INVx2_ASAP7_75t_L g306 ( .A(n_184), .Y(n_306) );
AND2x2_ASAP7_75t_L g322 ( .A(n_184), .B(n_323), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
O2A1O1Ixp5_ASAP7_75t_L g258 ( .A1(n_194), .A2(n_237), .B(n_259), .C(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_197), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx2_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
AND2x2_ASAP7_75t_L g385 ( .A(n_199), .B(n_201), .Y(n_385) );
AND2x2_ASAP7_75t_L g302 ( .A(n_200), .B(n_287), .Y(n_302) );
AND2x2_ASAP7_75t_L g401 ( .A(n_200), .B(n_402), .Y(n_401) );
NOR2xp67_ASAP7_75t_L g323 ( .A(n_201), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g426 ( .A(n_201), .B(n_287), .Y(n_426) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g212 ( .A(n_202), .Y(n_212) );
AND2x2_ASAP7_75t_L g305 ( .A(n_202), .B(n_306), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_205), .A2(n_237), .B(n_240), .C(n_241), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_205), .A2(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g229 ( .A(n_207), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_207), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
AND2x2_ASAP7_75t_L g351 ( .A(n_210), .B(n_286), .Y(n_351) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_211), .B(n_287), .Y(n_336) );
INVx2_ASAP7_75t_L g335 ( .A(n_212), .Y(n_335) );
OAI222xp33_ASAP7_75t_L g339 ( .A1(n_212), .A2(n_279), .B1(n_340), .B2(n_342), .C1(n_343), .C2(n_346), .Y(n_339) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g264 ( .A(n_217), .Y(n_264) );
OR2x2_ASAP7_75t_L g375 ( .A(n_217), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g297 ( .A(n_218), .Y(n_297) );
NOR2x1_ASAP7_75t_L g348 ( .A(n_218), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g354 ( .A(n_218), .B(n_268), .Y(n_354) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_L g315 ( .A(n_219), .Y(n_315) );
AO21x1_ASAP7_75t_L g314 ( .A1(n_221), .A2(n_224), .B(n_315), .Y(n_314) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_224), .A2(n_446), .B(n_459), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_224), .B(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g462 ( .A(n_224), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_224), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_224), .A2(n_517), .B(n_524), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_225), .A2(n_318), .B1(n_357), .B2(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_243), .Y(n_225) );
INVx3_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
OR2x2_ASAP7_75t_L g423 ( .A(n_226), .B(n_299), .Y(n_423) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g296 ( .A(n_227), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_227), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_227), .B(n_268), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_227), .B(n_244), .Y(n_376) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g267 ( .A(n_228), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g271 ( .A(n_228), .B(n_244), .Y(n_271) );
AND2x2_ASAP7_75t_L g347 ( .A(n_228), .B(n_294), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_228), .B(n_253), .Y(n_387) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_242), .Y(n_228) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_229), .A2(n_254), .B(n_261), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .C(n_235), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_233), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_233), .A2(n_522), .B(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_235), .A2(n_451), .B(n_452), .C(n_453), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_237), .A2(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_243), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_243), .B(n_264), .Y(n_303) );
AND2x2_ASAP7_75t_L g307 ( .A(n_243), .B(n_297), .Y(n_307) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
INVx3_ASAP7_75t_L g268 ( .A(n_244), .Y(n_268) );
AND2x2_ASAP7_75t_L g293 ( .A(n_244), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g428 ( .A(n_244), .B(n_411), .Y(n_428) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_253), .Y(n_282) );
INVx2_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
AND2x2_ASAP7_75t_L g338 ( .A(n_253), .B(n_314), .Y(n_338) );
INVx1_ASAP7_75t_L g381 ( .A(n_253), .Y(n_381) );
OR2x2_ASAP7_75t_L g412 ( .A(n_253), .B(n_314), .Y(n_412) );
AND2x2_ASAP7_75t_L g432 ( .A(n_253), .B(n_268), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_269), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g270 ( .A(n_264), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_264), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
INVx2_ASAP7_75t_SL g283 ( .A(n_267), .Y(n_283) );
AND2x2_ASAP7_75t_L g403 ( .A(n_267), .B(n_297), .Y(n_403) );
INVx2_ASAP7_75t_L g349 ( .A(n_268), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_268), .B(n_381), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .B1(n_275), .B2(n_281), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_271), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g437 ( .A(n_271), .Y(n_437) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g362 ( .A(n_273), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_273), .B(n_305), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_274), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g378 ( .A(n_274), .B(n_327), .Y(n_378) );
INVx2_ASAP7_75t_L g434 ( .A(n_274), .Y(n_434) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_277), .B(n_322), .Y(n_355) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_279), .B(n_299), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g416 ( .A(n_282), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_283), .A2(n_367), .B(n_369), .C(n_372), .Y(n_366) );
OR2x2_ASAP7_75t_L g393 ( .A(n_283), .B(n_297), .Y(n_393) );
OAI221xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_289), .B1(n_291), .B2(n_298), .C(n_301), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_286), .B(n_335), .Y(n_342) );
AND2x2_ASAP7_75t_L g384 ( .A(n_286), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g420 ( .A(n_286), .Y(n_420) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
NOR2xp67_ASAP7_75t_L g344 ( .A(n_290), .B(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g398 ( .A(n_290), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_290), .B(n_338), .Y(n_414) );
INVx2_ASAP7_75t_L g400 ( .A(n_291), .Y(n_400) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g341 ( .A(n_293), .B(n_312), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_293), .A2(n_309), .B(n_351), .C(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g319 ( .A(n_294), .B(n_314), .Y(n_319) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_298), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g367 ( .A(n_299), .B(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_304), .B2(n_307), .Y(n_301) );
INVx1_ASAP7_75t_L g421 ( .A(n_303), .Y(n_421) );
INVx1_ASAP7_75t_L g368 ( .A(n_305), .Y(n_368) );
INVx1_ASAP7_75t_L g419 ( .A(n_307), .Y(n_419) );
AOI211xp5_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_312), .B(n_316), .C(n_339), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g331 ( .A(n_311), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g382 ( .A(n_312), .Y(n_382) );
AND2x2_ASAP7_75t_L g431 ( .A(n_312), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B(n_329), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g345 ( .A(n_319), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_319), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g337 ( .A(n_320), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g413 ( .A(n_320), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g424 ( .A1(n_320), .A2(n_372), .A3(n_379), .B1(n_420), .B2(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_SL g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_SL g392 ( .A(n_322), .Y(n_392) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g332 ( .A(n_328), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B(n_337), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_331), .A2(n_379), .B1(n_405), .B2(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_335), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g365 ( .A(n_349), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_356), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_358), .A2(n_400), .B1(n_401), .B2(n_403), .C(n_404), .Y(n_399) );
NAND5xp2_ASAP7_75t_L g359 ( .A(n_360), .B(n_383), .C(n_399), .D(n_409), .E(n_427), .Y(n_359) );
AOI211xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_363), .B(n_366), .C(n_373), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g430 ( .A(n_367), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_377), .B2(n_379), .Y(n_373) );
INVx1_ASAP7_75t_SL g406 ( .A(n_376), .Y(n_406) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI322xp33_ASAP7_75t_L g388 ( .A1(n_379), .A2(n_389), .A3(n_390), .B1(n_391), .B2(n_392), .C1(n_393), .C2(n_394), .Y(n_388) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g391 ( .A(n_381), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_381), .B(n_406), .Y(n_405) );
AOI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_388), .C(n_396), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_392), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_418) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_417), .B1(n_418), .B2(n_422), .C(n_424), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_413), .B(n_414), .C(n_415), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g436 ( .A(n_412), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_430), .B2(n_431), .C(n_433), .Y(n_427) );
AOI21xp33_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B(n_436), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_441), .B(n_642), .Y(n_440) );
AND4x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_582), .C(n_597), .D(n_622), .Y(n_441) );
NOR2xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_555), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_473), .B(n_535), .Y(n_443) );
AND2x2_ASAP7_75t_L g585 ( .A(n_444), .B(n_490), .Y(n_585) );
AND2x2_ASAP7_75t_L g598 ( .A(n_444), .B(n_489), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_444), .B(n_474), .Y(n_648) );
INVx1_ASAP7_75t_L g652 ( .A(n_444), .Y(n_652) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_461), .Y(n_444) );
INVx2_ASAP7_75t_L g569 ( .A(n_445), .Y(n_569) );
BUFx2_ASAP7_75t_L g596 ( .A(n_445), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_456), .Y(n_446) );
INVx5_ASAP7_75t_L g466 ( .A(n_448), .Y(n_466) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_455), .A2(n_465), .B(n_466), .C(n_467), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_455), .A2(n_466), .B(n_546), .C(n_547), .Y(n_545) );
BUFx2_ASAP7_75t_L g493 ( .A(n_457), .Y(n_493) );
AND2x2_ASAP7_75t_L g536 ( .A(n_461), .B(n_490), .Y(n_536) );
INVx2_ASAP7_75t_L g552 ( .A(n_461), .Y(n_552) );
AND2x2_ASAP7_75t_L g561 ( .A(n_461), .B(n_489), .Y(n_561) );
AND2x2_ASAP7_75t_L g640 ( .A(n_461), .B(n_569), .Y(n_640) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_472), .Y(n_461) );
INVx2_ASAP7_75t_L g480 ( .A(n_466), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_502), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_474), .B(n_567), .Y(n_605) );
INVx1_ASAP7_75t_L g693 ( .A(n_474), .Y(n_693) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_489), .Y(n_474) );
AND2x2_ASAP7_75t_L g551 ( .A(n_475), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g565 ( .A(n_475), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_475), .Y(n_594) );
OR2x2_ASAP7_75t_L g626 ( .A(n_475), .B(n_568), .Y(n_626) );
AND2x2_ASAP7_75t_L g634 ( .A(n_475), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g667 ( .A(n_475), .B(n_636), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_475), .B(n_536), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_475), .B(n_596), .Y(n_692) );
AND2x2_ASAP7_75t_L g698 ( .A(n_475), .B(n_585), .Y(n_698) );
INVx5_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g558 ( .A(n_476), .Y(n_558) );
AND2x2_ASAP7_75t_L g588 ( .A(n_476), .B(n_568), .Y(n_588) );
AND2x2_ASAP7_75t_L g621 ( .A(n_476), .B(n_581), .Y(n_621) );
AND2x2_ASAP7_75t_L g641 ( .A(n_476), .B(n_490), .Y(n_641) );
AND2x2_ASAP7_75t_L g675 ( .A(n_476), .B(n_541), .Y(n_675) );
OR2x6_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_485), .C(n_486), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_483), .A2(n_486), .B(n_532), .C(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g581 ( .A(n_489), .B(n_552), .Y(n_581) );
AND2x2_ASAP7_75t_L g592 ( .A(n_489), .B(n_588), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_489), .B(n_568), .Y(n_631) );
INVx2_ASAP7_75t_L g646 ( .A(n_489), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_489), .B(n_580), .Y(n_669) );
AND2x2_ASAP7_75t_L g688 ( .A(n_489), .B(n_640), .Y(n_688) );
INVx5_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
AND2x2_ASAP7_75t_L g595 ( .A(n_490), .B(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g636 ( .A(n_490), .B(n_552), .Y(n_636) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_499), .Y(n_490) );
AOI21xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_494), .B(n_498), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
AND2x2_ASAP7_75t_L g559 ( .A(n_504), .B(n_542), .Y(n_559) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_505), .B(n_516), .Y(n_539) );
OR2x2_ASAP7_75t_L g572 ( .A(n_505), .B(n_542), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_505), .B(n_542), .Y(n_577) );
AND2x2_ASAP7_75t_L g604 ( .A(n_505), .B(n_541), .Y(n_604) );
AND2x2_ASAP7_75t_L g656 ( .A(n_505), .B(n_515), .Y(n_656) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_506), .B(n_526), .Y(n_564) );
AND2x2_ASAP7_75t_L g600 ( .A(n_506), .B(n_516), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_513), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g590 ( .A(n_514), .B(n_572), .Y(n_590) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_526), .Y(n_514) );
OAI322xp33_ASAP7_75t_L g555 ( .A1(n_515), .A2(n_556), .A3(n_560), .B1(n_562), .B2(n_565), .C1(n_570), .C2(n_578), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_515), .B(n_541), .Y(n_563) );
OR2x2_ASAP7_75t_L g573 ( .A(n_515), .B(n_527), .Y(n_573) );
AND2x2_ASAP7_75t_L g575 ( .A(n_515), .B(n_527), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_515), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_515), .B(n_542), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_515), .B(n_671), .Y(n_670) );
INVx5_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_516), .B(n_559), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_526), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g553 ( .A(n_526), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_526), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g615 ( .A(n_526), .B(n_542), .Y(n_615) );
AOI211xp5_ASAP7_75t_SL g643 ( .A1(n_526), .A2(n_644), .B(n_647), .C(n_659), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_526), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g681 ( .A(n_526), .B(n_656), .Y(n_681) );
INVx5_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g609 ( .A(n_527), .B(n_542), .Y(n_609) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_527), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_527), .B(n_656), .Y(n_658) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_527), .B(n_559), .Y(n_689) );
AND2x2_ASAP7_75t_L g696 ( .A(n_527), .B(n_655), .Y(n_696) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B1(n_551), .B2(n_553), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_536), .B(n_558), .Y(n_606) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g554 ( .A(n_539), .Y(n_554) );
OR2x2_ASAP7_75t_L g614 ( .A(n_539), .B(n_615), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g662 ( .A1(n_539), .A2(n_663), .B1(n_665), .B2(n_666), .C(n_668), .Y(n_662) );
INVx2_ASAP7_75t_L g601 ( .A(n_540), .Y(n_601) );
AND2x2_ASAP7_75t_L g574 ( .A(n_541), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g664 ( .A(n_541), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_541), .B(n_656), .Y(n_677) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVxp67_ASAP7_75t_L g619 ( .A(n_542), .Y(n_619) );
AND2x2_ASAP7_75t_L g655 ( .A(n_542), .B(n_656), .Y(n_655) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_550), .Y(n_542) );
AND2x2_ASAP7_75t_L g657 ( .A(n_551), .B(n_596), .Y(n_657) );
AND2x2_ASAP7_75t_L g567 ( .A(n_552), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_552), .B(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_SL g638 ( .A(n_554), .B(n_601), .Y(n_638) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g644 ( .A(n_557), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OR2x2_ASAP7_75t_L g630 ( .A(n_558), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g695 ( .A(n_558), .B(n_640), .Y(n_695) );
INVx2_ASAP7_75t_L g628 ( .A(n_559), .Y(n_628) );
NAND4xp25_ASAP7_75t_SL g691 ( .A(n_560), .B(n_692), .C(n_693), .D(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_561), .B(n_625), .Y(n_660) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_SL g697 ( .A(n_564), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_565), .A2(n_628), .B(n_632), .C(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g654 ( .A(n_567), .B(n_646), .Y(n_654) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_568), .Y(n_580) );
INVx1_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_569), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B(n_574), .C(n_576), .Y(n_570) );
AND2x2_ASAP7_75t_L g591 ( .A(n_571), .B(n_575), .Y(n_591) );
OAI322xp33_ASAP7_75t_SL g629 ( .A1(n_571), .A2(n_630), .A3(n_632), .B1(n_633), .B2(n_637), .C1(n_638), .C2(n_639), .Y(n_629) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g651 ( .A(n_573), .B(n_577), .Y(n_651) );
INVx1_ASAP7_75t_L g632 ( .A(n_575), .Y(n_632) );
INVx1_ASAP7_75t_SL g650 ( .A(n_577), .Y(n_650) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI222xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_589), .B1(n_591), .B2(n_592), .C1(n_593), .C2(n_726), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_584), .B(n_586), .Y(n_583) );
OAI322xp33_ASAP7_75t_L g672 ( .A1(n_584), .A2(n_646), .A3(n_651), .B1(n_673), .B2(n_674), .C1(n_676), .C2(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_585), .A2(n_599), .B1(n_623), .B2(n_627), .C(n_629), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OAI222xp33_ASAP7_75t_L g602 ( .A1(n_590), .A2(n_603), .B1(n_605), .B2(n_606), .C1(n_607), .C2(n_610), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_592), .A2(n_599), .B1(n_669), .B2(n_670), .Y(n_668) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_602), .C(n_613), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_599), .A2(n_636), .B(n_679), .C(n_682), .Y(n_678) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g608 ( .A(n_600), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g671 ( .A(n_604), .Y(n_671) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_611), .B(n_636), .Y(n_665) );
BUFx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_620), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g682 ( .A1(n_614), .A2(n_683), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_682) );
INVxp33_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_618), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_625), .B(n_636), .Y(n_676) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g687 ( .A(n_640), .B(n_646), .Y(n_687) );
AND4x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_661), .C(n_678), .D(n_690), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI221xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B1(n_651), .B2(n_652), .C(n_653), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_657), .B2(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g683 ( .A(n_654), .Y(n_683) );
INVx1_ASAP7_75t_SL g673 ( .A(n_658), .Y(n_673) );
NOR2xp33_ASAP7_75t_SL g661 ( .A(n_662), .B(n_672), .Y(n_661) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_674), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_681), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g707 ( .A(n_700), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx3_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
XNOR2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
endmodule