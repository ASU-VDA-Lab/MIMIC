module fake_jpeg_20844_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_8),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_19),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_31),
.B1(n_15),
.B2(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_27),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_10),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_21),
.B(n_20),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_41),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_18),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_43),
.C(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_20),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_51),
.B1(n_50),
.B2(n_45),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_38),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_17),
.B1(n_14),
.B2(n_11),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_35),
.B(n_43),
.Y(n_52)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_11),
.B(n_17),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_56),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_49),
.B1(n_39),
.B2(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_32),
.C(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_57),
.Y(n_61)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_1),
.C(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_58),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_2),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

AOI221xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_69),
.B1(n_70),
.B2(n_6),
.C(n_4),
.Y(n_72)
);


endmodule