module fake_ariane_2325_n_108 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_108);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_108;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_81;
wire n_87;
wire n_43;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_1),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_R g46 ( 
.A(n_28),
.B(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_27),
.B1(n_30),
.B2(n_25),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_36),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_46),
.B1(n_26),
.B2(n_29),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_32),
.B(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_54),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_55),
.B(n_34),
.C(n_48),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_60),
.B1(n_52),
.B2(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

AND3x1_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_49),
.C(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_67),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_77),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_73),
.C(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_72),
.Y(n_86)
);

NAND2x1p5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_3),
.Y(n_89)
);

AOI33xp33_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_23),
.A3(n_21),
.B1(n_49),
.B2(n_45),
.B3(n_3),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_36),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.C(n_93),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_84),
.B(n_87),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_45),
.B(n_52),
.Y(n_99)
);

AOI311xp33_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_4),
.A3(n_5),
.B(n_50),
.C(n_52),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_99),
.C(n_80),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_5),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NAND5xp2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_103),
.C(n_43),
.D(n_13),
.E(n_14),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_43),
.B1(n_80),
.B2(n_70),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_59),
.B(n_66),
.Y(n_108)
);


endmodule