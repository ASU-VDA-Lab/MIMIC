module fake_jpeg_2639_n_196 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_3),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_17),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_0),
.Y(n_89)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_61),
.B1(n_60),
.B2(n_55),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_84),
.B1(n_71),
.B2(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_65),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_55),
.B1(n_57),
.B2(n_64),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_102),
.B1(n_20),
.B2(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_57),
.B1(n_47),
.B2(n_52),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_99),
.B(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_54),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_72),
.B1(n_85),
.B2(n_47),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_54),
.B1(n_59),
.B2(n_68),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_62),
.B1(n_56),
.B2(n_78),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_46),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_62),
.B1(n_56),
.B2(n_76),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_23),
.B1(n_36),
.B2(n_33),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_126),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_121),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_63),
.B1(n_53),
.B2(n_86),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_120),
.B1(n_131),
.B2(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_86),
.B(n_90),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_109),
.B1(n_95),
.B2(n_92),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_103),
.B(n_99),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_1),
.B(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_18),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_21),
.B1(n_42),
.B2(n_41),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_117),
.C(n_120),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_142),
.C(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_16),
.C(n_31),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_5),
.Y(n_144)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_9),
.CI(n_10),
.CON(n_146),
.SN(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_9),
.Y(n_147)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_151),
.A2(n_133),
.B(n_137),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_24),
.C(n_30),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_165),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_149),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_152),
.B1(n_142),
.B2(n_146),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_11),
.B(n_12),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_14),
.B(n_15),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_25),
.C(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_173),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_170),
.B(n_163),
.Y(n_181)
);

AOI22x1_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_146),
.B1(n_150),
.B2(n_145),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_140),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_156),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_155),
.C(n_153),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_181),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_180),
.C(n_160),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_155),
.C(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_187),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_186),
.B1(n_188),
.B2(n_178),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_193),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_194),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_177),
.Y(n_196)
);


endmodule