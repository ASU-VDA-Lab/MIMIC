module real_jpeg_13068_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_35),
.B1(n_38),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_4),
.A2(n_35),
.B1(n_38),
.B2(n_69),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_42),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_8),
.B(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_62),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_9),
.A2(n_35),
.B1(n_38),
.B2(n_62),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_35),
.B1(n_38),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_12),
.A2(n_35),
.B1(n_38),
.B2(n_54),
.Y(n_106)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_89),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_83),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_83),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_58),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_45),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_21),
.B(n_33),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_26),
.C(n_30),
.Y(n_21)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OA22x2_ASAP7_75t_SL g65 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_23),
.B(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_31),
.C(n_32),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_27),
.A2(n_61),
.B1(n_64),
.B2(n_86),
.Y(n_85)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_29),
.CON(n_27),
.SN(n_27)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_28),
.A2(n_31),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_29),
.B(n_38),
.C(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_29),
.B(n_42),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_29),
.B(n_51),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B(n_41),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_34),
.B(n_40),
.Y(n_123)
);

CKINVDCx6p67_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_39),
.B(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_39),
.A2(n_40),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_79),
.B(n_81),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_42),
.A2(n_104),
.B1(n_112),
.B2(n_113),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_52),
.B(n_55),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_53),
.B1(n_56),
.B2(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_56),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_47),
.A2(n_56),
.B1(n_88),
.B2(n_99),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.C(n_87),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_87),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_130),
.B(n_134),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_119),
.B(n_129),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_107),
.B(n_118),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_100),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_113),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_114),
.B(n_117),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_121),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_125),
.C(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_133),
.Y(n_134)
);


endmodule