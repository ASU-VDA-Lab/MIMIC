module fake_jpeg_18466_n_252 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_11),
.B1(n_14),
.B2(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_33),
.B(n_26),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_41),
.B1(n_22),
.B2(n_16),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_52),
.B1(n_38),
.B2(n_41),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_16),
.B1(n_22),
.B2(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_43),
.B1(n_42),
.B2(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_75),
.B1(n_56),
.B2(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_67),
.B1(n_71),
.B2(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_69),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_37),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_48),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_43),
.B1(n_31),
.B2(n_27),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_54),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_70),
.C(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_44),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_86),
.B1(n_89),
.B2(n_66),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_73),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_66),
.B(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_47),
.B1(n_52),
.B2(n_40),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_79),
.A3(n_85),
.B1(n_75),
.B2(n_70),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_111),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_98),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_110),
.B1(n_92),
.B2(n_76),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_69),
.B1(n_74),
.B2(n_72),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_74),
.B1(n_58),
.B2(n_65),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_57),
.C(n_58),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_34),
.B(n_11),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_30),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_81),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_29),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_93),
.B1(n_84),
.B2(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_28),
.B1(n_87),
.B2(n_29),
.Y(n_148)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_60),
.B1(n_76),
.B2(n_17),
.Y(n_123)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_138),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_45),
.A3(n_27),
.B1(n_30),
.B2(n_26),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_53),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_111),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_160),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_144),
.B1(n_21),
.B2(n_19),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_99),
.B1(n_57),
.B2(n_45),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_21),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_114),
.B1(n_129),
.B2(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_122),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_53),
.C(n_12),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_12),
.C(n_14),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_12),
.C(n_23),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_12),
.C(n_23),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_120),
.C(n_124),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_23),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_163),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_115),
.B(n_17),
.CI(n_12),
.CON(n_163),
.SN(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_125),
.B(n_121),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_168),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_161),
.A2(n_125),
.B(n_133),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_132),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_173),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_124),
.B(n_138),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_174),
.A2(n_178),
.B1(n_181),
.B2(n_163),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_145),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_160),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_158),
.B1(n_147),
.B2(n_142),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_146),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_163),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_191),
.B1(n_19),
.B2(n_6),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_142),
.B(n_141),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_189),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_190),
.B(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_152),
.B1(n_159),
.B2(n_144),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_157),
.C(n_155),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_196),
.C(n_164),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_174),
.B1(n_176),
.B2(n_169),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_8),
.B(n_10),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_12),
.C(n_23),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_7),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_171),
.B(n_172),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_203),
.B(n_208),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_186),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_178),
.B(n_173),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_181),
.B1(n_164),
.B2(n_21),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_209),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_187),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_193),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_6),
.B(n_10),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_19),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_5),
.B(n_8),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_218),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_206),
.C(n_200),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_188),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_194),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_202),
.B1(n_6),
.B2(n_4),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_4),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_4),
.B(n_7),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_9),
.B(n_1),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_218),
.B1(n_212),
.B2(n_7),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_9),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_9),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_9),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_238),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_0),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_227),
.C(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_242),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_232),
.B(n_227),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_241),
.B(n_1),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_243),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_1),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_246),
.B(n_3),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_3),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_3),
.Y(n_252)
);


endmodule