module fake_netlist_1_9355_n_37 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
NOR2x1_ASAP7_75t_L g15 ( .A(n_10), .B(n_8), .Y(n_15) );
OA21x2_ASAP7_75t_L g16 ( .A1(n_7), .A2(n_6), .B(n_9), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_1), .B(n_11), .Y(n_17) );
INVx4_ASAP7_75t_L g18 ( .A(n_3), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_4), .B(n_2), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
INVxp67_ASAP7_75t_SL g21 ( .A(n_19), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_17), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_21), .B(n_18), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_20), .B1(n_22), .B2(n_19), .C(n_14), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AOI22xp33_ASAP7_75t_SL g30 ( .A1(n_28), .A2(n_24), .B1(n_22), .B2(n_17), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVxp33_ASAP7_75t_SL g32 ( .A(n_30), .Y(n_32) );
NAND5xp2_ASAP7_75t_L g33 ( .A(n_31), .B(n_29), .C(n_15), .D(n_2), .E(n_0), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
OAI22xp5_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_16), .B1(n_22), .B2(n_1), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_22), .B1(n_16), .B2(n_13), .Y(n_36) );
AOI22x1_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_34), .B1(n_16), .B2(n_12), .Y(n_37) );
endmodule