module fake_jpeg_18085_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_21),
.B(n_18),
.C(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_34),
.B(n_15),
.Y(n_38)
);

NOR2x1p5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_21),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_38),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_19),
.B(n_4),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_3),
.B(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_19),
.B1(n_14),
.B2(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_36),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_37),
.C(n_40),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_11),
.C(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_50),
.B1(n_38),
.B2(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_47),
.B1(n_49),
.B2(n_13),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_11),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_52),
.C1(n_45),
.C2(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);


endmodule