module fake_jpeg_11941_n_186 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_1),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_30),
.B(n_23),
.Y(n_65)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_10),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_68),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_2),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_65),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_17),
.B1(n_30),
.B2(n_19),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_66),
.B1(n_40),
.B2(n_43),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_15),
.B1(n_19),
.B2(n_18),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_20),
.B(n_16),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_44),
.C(n_33),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_9),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_92),
.B1(n_33),
.B2(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_39),
.B1(n_41),
.B2(n_54),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_59),
.A3(n_62),
.B1(n_4),
.B2(n_50),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_105),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_61),
.B1(n_81),
.B2(n_55),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_119),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_99),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_122),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_75),
.C(n_58),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_55),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_4),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_93),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_112),
.C(n_124),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_97),
.B(n_87),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_134),
.B(n_108),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_94),
.B(n_103),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_84),
.B(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_45),
.B1(n_75),
.B2(n_39),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_69),
.B1(n_100),
.B2(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_69),
.B1(n_102),
.B2(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_145),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_118),
.B(n_126),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_134),
.B(n_129),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_125),
.C(n_121),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_141),
.C(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_159),
.C(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_164),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_130),
.B1(n_135),
.B2(n_140),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_155),
.B1(n_143),
.B2(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_132),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_150),
.B1(n_147),
.B2(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_161),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_130),
.B1(n_152),
.B2(n_135),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_159),
.B1(n_160),
.B2(n_156),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.C(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_175),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_169),
.C(n_165),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_180),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_168),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_146),
.B1(n_151),
.B2(n_121),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_177),
.B1(n_125),
.B2(n_126),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_182),
.C(n_179),
.Y(n_184)
);

AOI21x1_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_182),
.B(n_93),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_185),
.Y(n_186)
);


endmodule