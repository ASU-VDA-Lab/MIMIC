module fake_netlist_1_7317_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
AO21x2_ASAP7_75t_L g12 ( .A1(n_0), .A2(n_4), .B(n_5), .Y(n_12) );
NAND3xp33_ASAP7_75t_L g13 ( .A(n_3), .B(n_1), .C(n_2), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
AOI21x1_ASAP7_75t_L g16 ( .A1(n_4), .A2(n_7), .B(n_0), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_10), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_6), .Y(n_19) );
AOI221x1_ASAP7_75t_L g20 ( .A1(n_10), .A2(n_9), .B1(n_15), .B2(n_14), .C(n_11), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_15), .Y(n_21) );
OAI22xp5_ASAP7_75t_L g22 ( .A1(n_11), .A2(n_14), .B1(n_13), .B2(n_17), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_12), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_23), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
OAI22xp33_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_18), .B1(n_22), .B2(n_16), .Y(n_27) );
O2A1O1Ixp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B(n_18), .C(n_16), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_28), .B(n_25), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_24), .Y(n_30) );
AOI22xp5_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_17), .B1(n_12), .B2(n_20), .Y(n_31) );
AOI211xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_12), .B(n_17), .C(n_22), .Y(n_32) );
OAI21xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_17), .B(n_31), .Y(n_33) );
endmodule