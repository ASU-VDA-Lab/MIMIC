module fake_aes_7371_n_18 (n_1, n_2, n_4, n_3, n_5, n_0, n_18);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_17;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
AND2x2_ASAP7_75t_L g6 ( .A(n_2), .B(n_4), .Y(n_6) );
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_4), .B(n_1), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_0), .Y(n_9) );
INVx2_ASAP7_75t_SL g10 ( .A(n_8), .Y(n_10) );
OAI21xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_0), .B(n_1), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_9), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_10), .B(n_6), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
OAI221xp5_ASAP7_75t_SL g15 ( .A1(n_14), .A2(n_12), .B1(n_13), .B2(n_6), .C(n_11), .Y(n_15) );
INVx1_ASAP7_75t_SL g16 ( .A(n_15), .Y(n_16) );
NAND3xp33_ASAP7_75t_L g17 ( .A(n_15), .B(n_7), .C(n_3), .Y(n_17) );
AOI31xp33_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_2), .A3(n_5), .B(n_17), .Y(n_18) );
endmodule