module fake_jpeg_4058_n_302 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_46)
);

AOI22x1_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_40),
.B1(n_26),
.B2(n_17),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_42),
.B1(n_41),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_60),
.B1(n_62),
.B2(n_19),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_64),
.Y(n_80)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_18),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_23),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_23),
.Y(n_87)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_67),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_37),
.A3(n_43),
.B1(n_21),
.B2(n_42),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_60),
.C(n_34),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx11_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_89),
.B1(n_92),
.B2(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_81),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_95),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_93),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_12),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_94),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_19),
.B1(n_27),
.B2(n_43),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_43),
.Y(n_92)
);

BUFx16f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_21),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_10),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_99),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_11),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_121),
.Y(n_133)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_117),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_44),
.B1(n_64),
.B2(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_98),
.B1(n_108),
.B2(n_113),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_44),
.C(n_45),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_79),
.C(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_69),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_84),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_123),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_58),
.B1(n_45),
.B2(n_32),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_82),
.B1(n_65),
.B2(n_76),
.Y(n_129)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_45),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_20),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_20),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_78),
.B(n_68),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_147),
.B(n_32),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_113),
.B1(n_118),
.B2(n_98),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_129),
.B1(n_136),
.B2(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_153),
.C(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_138),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_96),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_88),
.B1(n_93),
.B2(n_28),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_95),
.B(n_93),
.C(n_20),
.D(n_34),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_9),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_34),
.B(n_20),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_10),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_20),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_106),
.B1(n_100),
.B2(n_110),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_100),
.B1(n_111),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_160),
.B1(n_172),
.B2(n_141),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_163),
.C(n_171),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_111),
.B1(n_105),
.B2(n_114),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_77),
.C(n_101),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_179),
.B(n_3),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_136),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_101),
.C(n_67),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_32),
.B1(n_28),
.B2(n_34),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_28),
.C(n_1),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_126),
.C(n_139),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_184),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_5),
.B1(n_13),
.B2(n_9),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_4),
.B1(n_8),
.B2(n_6),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_131),
.B(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_189),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_200),
.B(n_159),
.Y(n_229)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_206),
.B1(n_185),
.B2(n_162),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_149),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_192),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_201),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_155),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_209),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_211),
.Y(n_230)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_159),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_222),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_166),
.B(n_175),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_155),
.B1(n_175),
.B2(n_183),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_200),
.B1(n_206),
.B2(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_156),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_186),
.B(n_196),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_165),
.B1(n_181),
.B2(n_179),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_203),
.B1(n_211),
.B2(n_187),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_194),
.B1(n_210),
.B2(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_202),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_239),
.B(n_243),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_198),
.C(n_193),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_191),
.B(n_195),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_245),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_200),
.B1(n_195),
.B2(n_208),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_199),
.C(n_205),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_227),
.C(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_248),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_203),
.B1(n_165),
.B2(n_168),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_170),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_214),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_257),
.B(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_167),
.Y(n_256)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_220),
.C(n_215),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_221),
.C(n_213),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_262),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_241),
.A2(n_230),
.B(n_212),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_237),
.B(n_250),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_221),
.C(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_242),
.B(n_244),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_269),
.B(n_274),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_178),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_247),
.C(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_251),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_248),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_259),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_283),
.B(n_285),
.Y(n_288)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_284),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_257),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_242),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_255),
.C(n_270),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.C(n_4),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_293),
.B(n_4),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_269),
.C(n_265),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_234),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_281),
.A3(n_267),
.B1(n_251),
.B2(n_231),
.C1(n_167),
.C2(n_178),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_295),
.A3(n_288),
.B1(n_291),
.B2(n_5),
.C1(n_8),
.C2(n_16),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_3),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_297),
.B(n_5),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.C(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_1),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_2),
.C(n_300),
.Y(n_302)
);


endmodule