module fake_jpeg_26916_n_62 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_11),
.B1(n_21),
.B2(n_20),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_27),
.B1(n_25),
.B2(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_4),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_24),
.B(n_27),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_5),
.C(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_12),
.B(n_19),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_8),
.C(n_14),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_54),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_52),
.B(n_57),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_50),
.B1(n_39),
.B2(n_37),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_37),
.C(n_15),
.Y(n_62)
);


endmodule