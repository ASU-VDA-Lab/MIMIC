module fake_netlist_5_1826_n_75 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_75);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_75;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_70;
wire n_38;
wire n_71;
wire n_61;
wire n_68;
wire n_72;
wire n_35;
wire n_41;
wire n_32;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_74;
wire n_73;
wire n_19;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_52;
wire n_49;
wire n_60;
wire n_20;
wire n_39;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_1),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

OR2x6_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

OAI221xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.C(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_40),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.C(n_45),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_42),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_20),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_44),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

NAND2xp67_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_47),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_48),
.B1(n_56),
.B2(n_21),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_47),
.B(n_22),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_48),
.B(n_28),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_26),
.B(n_32),
.Y(n_64)
);

AOI321xp33_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OAI211xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_26),
.B(n_25),
.C(n_19),
.Y(n_67)
);

NAND4xp75_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.C(n_4),
.D(n_3),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_63),
.B(n_66),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NOR2xp67_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_69),
.B1(n_19),
.B2(n_18),
.Y(n_73)
);

AOI22x1_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_19),
.B1(n_10),
.B2(n_11),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_19),
.B1(n_72),
.B2(n_74),
.Y(n_75)
);


endmodule