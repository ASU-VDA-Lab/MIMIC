module fake_jpeg_30849_n_252 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_14),
.B(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_6),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_51),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_18),
.A2(n_8),
.B1(n_11),
.B2(n_2),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_8),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_65),
.B(n_91),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_28),
.C(n_23),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_76),
.C(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_77),
.B1(n_92),
.B2(n_97),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_29),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_20),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_29),
.B(n_28),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_9),
.Y(n_121)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_43),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_93),
.Y(n_119)
);

AOI31xp33_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_27),
.A3(n_26),
.B(n_24),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_20),
.B1(n_15),
.B2(n_23),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_24),
.C(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_21),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_41),
.A2(n_20),
.B1(n_16),
.B2(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_44),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_2),
.B1(n_5),
.B2(n_9),
.Y(n_118)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

BUFx6f_ASAP7_75t_SL g101 ( 
.A(n_35),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_125),
.Y(n_139)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_76),
.B1(n_62),
.B2(n_101),
.Y(n_130)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_122),
.Y(n_147)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_86),
.B1(n_62),
.B2(n_64),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_124),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_1),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_69),
.C(n_58),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_67),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_63),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_66),
.B(n_1),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_73),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_135),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_66),
.B1(n_85),
.B2(n_79),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_137),
.B1(n_146),
.B2(n_104),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_75),
.B1(n_96),
.B2(n_67),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_138),
.B1(n_143),
.B2(n_144),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_71),
.B(n_86),
.C(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_145),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_61),
.C(n_78),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_142),
.C(n_104),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_100),
.B1(n_79),
.B2(n_89),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_78),
.B(n_87),
.C(n_64),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_89),
.B1(n_87),
.B2(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_73),
.B1(n_70),
.B2(n_84),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_70),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_10),
.B(n_128),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_115),
.B(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_122),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_155),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_126),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_113),
.A2(n_102),
.B1(n_114),
.B2(n_109),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_157),
.A2(n_102),
.B(n_109),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_154),
.B(n_133),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_110),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_174),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_165),
.Y(n_184)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_148),
.A3(n_132),
.B1(n_143),
.B2(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_177),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_117),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_117),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_147),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_144),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_197),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_138),
.B1(n_153),
.B2(n_156),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_195),
.B1(n_199),
.B2(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_181),
.C(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_104),
.B1(n_133),
.B2(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_203),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_172),
.B(n_166),
.C(n_171),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_162),
.C(n_173),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_174),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_173),
.C(n_159),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_212),
.C(n_188),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_161),
.Y(n_212)
);

NOR4xp25_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_170),
.C(n_167),
.D(n_168),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_199),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_164),
.C(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_212),
.C(n_205),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_192),
.C(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_224),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_211),
.B(n_210),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_184),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_203),
.C(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_229),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_207),
.B(n_195),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_211),
.B(n_187),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_216),
.C(n_205),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_182),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_216),
.C(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_238),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_182),
.C(n_198),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_239),
.B(n_194),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_183),
.Y(n_240)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_244),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_238),
.B(n_237),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_233),
.B(n_187),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_240),
.B(n_198),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.C(n_245),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_164),
.B1(n_186),
.B2(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_186),
.Y(n_252)
);


endmodule