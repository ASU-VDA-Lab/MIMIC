module fake_jpeg_9949_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_1),
.B(n_5),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_1),
.B(n_0),
.Y(n_8)
);

CKINVDCx14_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_15),
.A2(n_17),
.B1(n_13),
.B2(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_3),
.B1(n_4),
.B2(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_20),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2x1p5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_9),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_12),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_10),
.C(n_9),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_26),
.C(n_28),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_7),
.B(n_11),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_17),
.B(n_21),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_12),
.C(n_13),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_13),
.B1(n_21),
.B2(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_32),
.B(n_33),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_35),
.B1(n_25),
.B2(n_22),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.C(n_32),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_40),
.C(n_37),
.Y(n_42)
);


endmodule