module real_aes_1621_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_835, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_836, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_835;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_836;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g180 ( .A(n_0), .B(n_154), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_1), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_2), .B(n_114), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_3), .Y(n_832) );
INVx1_ASAP7_75t_L g145 ( .A(n_4), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_5), .B(n_138), .Y(n_207) );
NAND2xp33_ASAP7_75t_SL g250 ( .A(n_6), .B(n_144), .Y(n_250) );
INVx1_ASAP7_75t_L g242 ( .A(n_7), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_8), .B(n_212), .Y(n_499) );
INVx1_ASAP7_75t_L g480 ( .A(n_9), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_10), .Y(n_114) );
AND2x2_ASAP7_75t_L g205 ( .A(n_11), .B(n_162), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_12), .Y(n_563) );
INVx2_ASAP7_75t_L g160 ( .A(n_13), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_14), .Y(n_116) );
INVx1_ASAP7_75t_L g507 ( .A(n_15), .Y(n_507) );
AOI221x1_ASAP7_75t_L g245 ( .A1(n_16), .A2(n_147), .B1(n_246), .B2(n_248), .C(n_249), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_17), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_19), .Y(n_799) );
INVx1_ASAP7_75t_L g505 ( .A(n_20), .Y(n_505) );
INVx1_ASAP7_75t_SL g517 ( .A(n_21), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_22), .B(n_139), .Y(n_495) );
AOI221xp5_ASAP7_75t_SL g169 ( .A1(n_23), .A2(n_44), .B1(n_138), .B2(n_147), .C(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_24), .A2(n_147), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_25), .B(n_154), .Y(n_210) );
AOI33xp33_ASAP7_75t_L g472 ( .A1(n_26), .A2(n_56), .A3(n_193), .B1(n_200), .B2(n_473), .B3(n_474), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_27), .A2(n_42), .B1(n_824), .B2(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_27), .Y(n_825) );
INVx1_ASAP7_75t_L g557 ( .A(n_28), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_29), .A2(n_120), .B1(n_121), .B2(n_127), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_29), .Y(n_127) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_30), .A2(n_93), .B(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g163 ( .A(n_30), .B(n_93), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_31), .B(n_156), .Y(n_155) );
INVxp67_ASAP7_75t_L g244 ( .A(n_32), .Y(n_244) );
AND2x2_ASAP7_75t_L g231 ( .A(n_33), .B(n_168), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_34), .B(n_191), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_35), .A2(n_147), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_36), .B(n_660), .Y(n_659) );
CKINVDCx16_ASAP7_75t_R g783 ( .A(n_36), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_37), .B(n_156), .Y(n_171) );
AND2x2_ASAP7_75t_L g144 ( .A(n_38), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g148 ( .A(n_38), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g199 ( .A(n_38), .Y(n_199) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_39), .B(n_113), .C(n_115), .Y(n_112) );
OR2x6_ASAP7_75t_L g787 ( .A(n_39), .B(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_40), .A2(n_73), .B1(n_820), .B2(n_821), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_40), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_41), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_42), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_43), .B(n_191), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_45), .A2(n_122), .B1(n_123), .B2(n_124), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_45), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_46), .A2(n_176), .B1(n_212), .B2(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_47), .A2(n_85), .B1(n_147), .B2(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_48), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_49), .B(n_139), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_50), .B(n_154), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_51), .B(n_158), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_52), .B(n_139), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_53), .Y(n_492) );
AND2x2_ASAP7_75t_L g183 ( .A(n_54), .B(n_168), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_55), .B(n_168), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_57), .B(n_139), .Y(n_463) );
INVx1_ASAP7_75t_L g141 ( .A(n_58), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_58), .Y(n_151) );
AND2x2_ASAP7_75t_L g464 ( .A(n_59), .B(n_168), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_60), .A2(n_78), .B1(n_191), .B2(n_197), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_61), .B(n_191), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_62), .B(n_138), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_63), .B(n_176), .Y(n_565) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_64), .A2(n_197), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g222 ( .A(n_65), .B(n_168), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_66), .B(n_156), .Y(n_181) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_67), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_68), .B(n_154), .Y(n_219) );
INVx1_ASAP7_75t_L g502 ( .A(n_69), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_70), .A2(n_147), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g461 ( .A(n_71), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_72), .B(n_156), .Y(n_211) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_73), .B(n_158), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_73), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_74), .A2(n_197), .B(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_75), .A2(n_97), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_75), .Y(n_125) );
INVx1_ASAP7_75t_L g143 ( .A(n_76), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_76), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_77), .B(n_191), .Y(n_475) );
AND2x2_ASAP7_75t_L g519 ( .A(n_79), .B(n_248), .Y(n_519) );
INVx1_ASAP7_75t_L g503 ( .A(n_80), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_81), .A2(n_197), .B(n_516), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_82), .A2(n_188), .B(n_197), .C(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_83), .A2(n_88), .B1(n_138), .B2(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_84), .B(n_138), .Y(n_220) );
INVx1_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_87), .B(n_248), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_89), .A2(n_197), .B1(n_470), .B2(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_90), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_91), .B(n_154), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_92), .A2(n_147), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g527 ( .A(n_94), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_95), .B(n_156), .Y(n_218) );
AND2x2_ASAP7_75t_L g476 ( .A(n_96), .B(n_248), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_97), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_98), .A2(n_555), .B(n_556), .C(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_99), .B(n_138), .Y(n_182) );
INVxp67_ASAP7_75t_L g247 ( .A(n_100), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_101), .B(n_156), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_102), .A2(n_147), .B(n_152), .Y(n_146) );
BUFx2_ASAP7_75t_L g810 ( .A(n_103), .Y(n_810) );
BUFx2_ASAP7_75t_SL g830 ( .A(n_103), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_104), .B(n_139), .Y(n_528) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_117), .B(n_831), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_107), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_SL g108 ( .A(n_109), .B(n_112), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_110), .B(n_111), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_115), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_116), .B(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_SL g793 ( .A(n_116), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_116), .B(n_794), .Y(n_804) );
OR2x2_ASAP7_75t_L g808 ( .A(n_116), .B(n_787), .Y(n_808) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_811), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_128), .B(n_785), .C(n_789), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_119), .A2(n_786), .B(n_787), .Y(n_785) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_119), .Y(n_796) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
OAI21xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_444), .B(n_445), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_SL g795 ( .A(n_130), .Y(n_795) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_336), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_264), .C(n_314), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_184), .B(n_232), .C(n_253), .Y(n_132) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_164), .Y(n_133) );
AND2x2_ASAP7_75t_L g263 ( .A(n_134), .B(n_165), .Y(n_263) );
INVx1_ASAP7_75t_L g394 ( .A(n_134), .Y(n_394) );
NOR2x1p5_ASAP7_75t_L g426 ( .A(n_134), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g237 ( .A(n_135), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g285 ( .A(n_135), .Y(n_285) );
OR2x2_ASAP7_75t_L g289 ( .A(n_135), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_135), .B(n_167), .Y(n_301) );
OR2x2_ASAP7_75t_L g323 ( .A(n_135), .B(n_167), .Y(n_323) );
AND2x4_ASAP7_75t_L g329 ( .A(n_135), .B(n_293), .Y(n_329) );
OR2x2_ASAP7_75t_L g346 ( .A(n_135), .B(n_239), .Y(n_346) );
INVx1_ASAP7_75t_L g381 ( .A(n_135), .Y(n_381) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_135), .Y(n_403) );
OR2x2_ASAP7_75t_L g417 ( .A(n_135), .B(n_350), .Y(n_417) );
AND2x4_ASAP7_75t_SL g421 ( .A(n_135), .B(n_239), .Y(n_421) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_161), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_158), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g251 ( .A(n_139), .Y(n_251) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x6_ASAP7_75t_L g154 ( .A(n_140), .B(n_149), .Y(n_154) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g156 ( .A(n_142), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_144), .Y(n_558) );
AND2x2_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
INVx2_ASAP7_75t_L g201 ( .A(n_149), .Y(n_201) );
AND2x4_ASAP7_75t_L g197 ( .A(n_150), .B(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
INVxp67_ASAP7_75t_L g506 ( .A(n_154), .Y(n_506) );
INVxp67_ASAP7_75t_L g508 ( .A(n_156), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_157), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_157), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_157), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_157), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_157), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_157), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g470 ( .A(n_157), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_157), .A2(n_462), .B(n_480), .C(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_157), .A2(n_495), .B(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_157), .B(n_212), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_157), .A2(n_462), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_157), .A2(n_462), .B(n_527), .C(n_528), .Y(n_526) );
INVx2_ASAP7_75t_SL g188 ( .A(n_158), .Y(n_188) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_158), .A2(n_478), .B(n_482), .Y(n_477) );
BUFx4f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_160), .B(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g212 ( .A(n_160), .B(n_163), .Y(n_212) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_162), .Y(n_168) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g373 ( .A(n_165), .B(n_329), .Y(n_373) );
AND2x2_ASAP7_75t_L g420 ( .A(n_165), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_174), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
AND2x2_ASAP7_75t_L g283 ( .A(n_167), .B(n_174), .Y(n_283) );
INVx2_ASAP7_75t_L g290 ( .A(n_167), .Y(n_290) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_167), .Y(n_411) );
BUFx3_ASAP7_75t_L g427 ( .A(n_167), .Y(n_427) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_173), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_168), .Y(n_221) );
INVx2_ASAP7_75t_L g252 ( .A(n_174), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_174), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g350 ( .A(n_174), .B(n_290), .Y(n_350) );
INVx1_ASAP7_75t_L g368 ( .A(n_174), .Y(n_368) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_174), .Y(n_384) );
INVx1_ASAP7_75t_L g406 ( .A(n_174), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_174), .B(n_285), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_174), .B(n_239), .Y(n_443) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21x1_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_183), .Y(n_175) );
INVx4_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_176), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_182), .Y(n_177) );
INVx1_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_203), .Y(n_185) );
AND2x4_ASAP7_75t_L g257 ( .A(n_186), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g268 ( .A(n_186), .Y(n_268) );
AND2x2_ASAP7_75t_L g273 ( .A(n_186), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g308 ( .A(n_186), .B(n_213), .Y(n_308) );
AND2x2_ASAP7_75t_L g318 ( .A(n_186), .B(n_214), .Y(n_318) );
OR2x2_ASAP7_75t_L g398 ( .A(n_186), .B(n_313), .Y(n_398) );
OAI322xp33_ASAP7_75t_L g428 ( .A1(n_186), .A2(n_341), .A3(n_380), .B1(n_413), .B2(n_429), .C1(n_430), .C2(n_431), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_186), .B(n_411), .Y(n_429) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
AOI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_202), .Y(n_187) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_188), .A2(n_468), .B(n_476), .Y(n_467) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_188), .A2(n_468), .B(n_476), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_196), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_191), .A2(n_197), .B1(n_241), .B2(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g566 ( .A(n_191), .Y(n_566) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_195), .Y(n_191) );
INVx1_ASAP7_75t_L g490 ( .A(n_192), .Y(n_490) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
OR2x6_ASAP7_75t_L g462 ( .A(n_193), .B(n_201), .Y(n_462) );
INVxp33_ASAP7_75t_L g473 ( .A(n_193), .Y(n_473) );
INVx1_ASAP7_75t_L g491 ( .A(n_195), .Y(n_491) );
INVxp67_ASAP7_75t_L g564 ( .A(n_197), .Y(n_564) );
NOR2x1p5_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g474 ( .A(n_200), .Y(n_474) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_203), .A2(n_375), .B1(n_379), .B2(n_382), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g434 ( .A1(n_203), .A2(n_435), .B(n_436), .C(n_439), .Y(n_434) );
AND2x4_ASAP7_75t_SL g203 ( .A(n_204), .B(n_213), .Y(n_203) );
AND2x4_ASAP7_75t_L g256 ( .A(n_204), .B(n_224), .Y(n_256) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_204), .Y(n_260) );
INVx5_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
INVx2_ASAP7_75t_L g281 ( .A(n_204), .Y(n_281) );
AND2x2_ASAP7_75t_L g304 ( .A(n_204), .B(n_214), .Y(n_304) );
AND2x2_ASAP7_75t_L g333 ( .A(n_204), .B(n_223), .Y(n_333) );
OR2x2_ASAP7_75t_L g342 ( .A(n_204), .B(n_262), .Y(n_342) );
OR2x2_ASAP7_75t_L g357 ( .A(n_204), .B(n_271), .Y(n_357) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_212), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_212), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_212), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_212), .B(n_247), .Y(n_246) );
NOR3xp33_ASAP7_75t_L g249 ( .A(n_212), .B(n_250), .C(n_251), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_212), .A2(n_525), .B(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_213), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_SL g341 ( .A(n_213), .Y(n_341) );
AND2x2_ASAP7_75t_L g364 ( .A(n_213), .B(n_272), .Y(n_364) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
INVx2_ASAP7_75t_L g258 ( .A(n_214), .Y(n_258) );
AND2x2_ASAP7_75t_L g261 ( .A(n_214), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g275 ( .A(n_214), .B(n_224), .Y(n_275) );
INVx1_ASAP7_75t_L g279 ( .A(n_214), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_214), .B(n_224), .Y(n_313) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_214), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_214), .B(n_272), .Y(n_388) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_221), .B(n_222), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_221), .A2(n_225), .B(n_231), .Y(n_224) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_221), .A2(n_225), .B(n_231), .Y(n_271) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_221), .A2(n_513), .B(n_519), .Y(n_512) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_224), .Y(n_294) );
AND2x2_ASAP7_75t_L g378 ( .A(n_224), .B(n_262), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_230), .Y(n_225) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_234), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x6_ASAP7_75t_SL g442 ( .A(n_235), .B(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_236), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_236), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g390 ( .A(n_236), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_237), .A2(n_299), .B1(n_302), .B2(n_309), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_238), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_238), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_238), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_238), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_252), .Y(n_238) );
AND2x2_ASAP7_75t_L g284 ( .A(n_239), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g293 ( .A(n_239), .Y(n_293) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_239), .A2(n_300), .B1(n_352), .B2(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g359 ( .A(n_239), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_239), .B(n_353), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_239), .B(n_283), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_239), .B(n_290), .Y(n_432) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_245), .Y(n_239) );
INVx3_ASAP7_75t_L g456 ( .A(n_248), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_248), .A2(n_456), .B1(n_554), .B2(n_559), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_251), .A2(n_462), .B1(n_502), .B2(n_503), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_251), .B(n_557), .Y(n_556) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_259), .B(n_263), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NAND4xp25_ASAP7_75t_SL g302 ( .A(n_255), .B(n_303), .C(n_305), .D(n_307), .Y(n_302) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_256), .B(n_363), .Y(n_392) );
AND2x2_ASAP7_75t_L g419 ( .A(n_256), .B(n_257), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_256), .B(n_279), .Y(n_430) );
INVx1_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_257), .A2(n_320), .B1(n_331), .B2(n_334), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g352 ( .A(n_257), .B(n_270), .C(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_257), .B(n_272), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_257), .B(n_280), .Y(n_423) );
AND2x2_ASAP7_75t_L g355 ( .A(n_258), .B(n_262), .Y(n_355) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_258), .Y(n_416) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
INVx1_ASAP7_75t_L g401 ( .A(n_261), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_261), .B(n_272), .Y(n_408) );
BUFx2_ASAP7_75t_L g363 ( .A(n_262), .Y(n_363) );
NAND3xp33_ASAP7_75t_SL g264 ( .A(n_265), .B(n_286), .C(n_298), .Y(n_264) );
OAI31xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_273), .A3(n_276), .B(n_282), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_266), .A2(n_320), .B1(n_324), .B2(n_325), .Y(n_319) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OR2x2_ASAP7_75t_L g305 ( .A(n_268), .B(n_306), .Y(n_305) );
NOR2x1_ASAP7_75t_L g331 ( .A(n_268), .B(n_332), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_269), .A2(n_371), .B(n_401), .C(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_270), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_271), .B(n_279), .Y(n_306) );
AND2x2_ASAP7_75t_L g324 ( .A(n_271), .B(n_304), .Y(n_324) );
AND2x2_ASAP7_75t_L g441 ( .A(n_274), .B(n_363), .Y(n_441) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g297 ( .A(n_275), .B(n_281), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_280), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g372 ( .A(n_280), .B(n_355), .Y(n_372) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_281), .B(n_355), .Y(n_361) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g353 ( .A(n_283), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_284), .B(n_384), .Y(n_383) );
AOI32xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_294), .A3(n_295), .B1(n_296), .B2(n_835), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_287), .A2(n_372), .B1(n_408), .B2(n_409), .C(n_412), .Y(n_407) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g300 ( .A(n_292), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g405 ( .A(n_293), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_294), .B(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_296), .A2(n_339), .B1(n_343), .B2(n_347), .C(n_351), .Y(n_338) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI211xp5_ASAP7_75t_L g314 ( .A1(n_301), .A2(n_315), .B(n_319), .C(n_330), .Y(n_314) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI322xp33_ASAP7_75t_L g412 ( .A1(n_307), .A2(n_317), .A3(n_366), .B1(n_413), .B2(n_414), .C1(n_415), .C2(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_310), .A2(n_440), .B(n_442), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_316), .A2(n_397), .B(n_399), .C(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g438 ( .A(n_323), .B(n_404), .Y(n_438) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_329), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g413 ( .A(n_329), .Y(n_413) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI31xp33_ASAP7_75t_L g369 ( .A1(n_333), .A2(n_370), .A3(n_372), .B(n_373), .Y(n_369) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_395), .Y(n_336) );
NAND5xp2_ASAP7_75t_L g337 ( .A(n_338), .B(n_358), .C(n_369), .D(n_374), .E(n_385), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_341), .A2(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g409 ( .A(n_345), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B(n_362), .C(n_365), .Y(n_358) );
INVxp33_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g387 ( .A(n_363), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_366), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g437 ( .A(n_378), .Y(n_437) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_387), .A2(n_392), .B(n_393), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_396), .B(n_407), .C(n_418), .D(n_434), .Y(n_395) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_405), .B(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g435 ( .A(n_417), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_428), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g786 ( .A(n_445), .Y(n_786) );
INVx2_ASAP7_75t_L g817 ( .A(n_446), .Y(n_817) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_780), .Y(n_446) );
NOR4xp25_ASAP7_75t_L g447 ( .A(n_448), .B(n_659), .C(n_683), .D(n_749), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_448), .A2(n_683), .B1(n_783), .B2(n_836), .Y(n_784) );
NAND3x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_611), .C(n_645), .Y(n_448) );
NOR3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_570), .C(n_590), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_545), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_483), .B1(n_534), .B2(n_542), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_465), .Y(n_452) );
AND2x2_ASAP7_75t_L g709 ( .A(n_453), .B(n_639), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_453), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_453), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_453), .B(n_579), .Y(n_768) );
OR2x2_ASAP7_75t_L g778 ( .A(n_453), .B(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_454), .B(n_536), .Y(n_599) );
AND2x4_ASAP7_75t_L g627 ( .A(n_454), .B(n_541), .Y(n_627) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g575 ( .A(n_455), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_455), .B(n_467), .Y(n_665) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_455), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_455), .B(n_552), .Y(n_702) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B(n_464), .Y(n_455) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_456), .A2(n_457), .B(n_464), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g497 ( .A(n_462), .Y(n_497) );
INVxp67_ASAP7_75t_L g555 ( .A(n_462), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_465), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g773 ( .A(n_465), .B(n_610), .Y(n_773) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g763 ( .A(n_466), .B(n_702), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
INVx2_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g537 ( .A(n_477), .Y(n_537) );
INVx2_ASAP7_75t_L g551 ( .A(n_477), .Y(n_551) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_477), .Y(n_576) );
INVx1_ASAP7_75t_L g589 ( .A(n_477), .Y(n_589) );
INVxp67_ASAP7_75t_L g608 ( .A(n_477), .Y(n_608) );
AND2x4_ASAP7_75t_L g639 ( .A(n_477), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_520), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_510), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g681 ( .A(n_486), .B(n_668), .Y(n_681) );
AND2x2_ASAP7_75t_L g705 ( .A(n_486), .B(n_521), .Y(n_705) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
INVx2_ASAP7_75t_L g533 ( .A(n_487), .Y(n_533) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
INVx1_ASAP7_75t_L g605 ( .A(n_487), .Y(n_605) );
AND2x4_ASAP7_75t_L g614 ( .A(n_487), .B(n_532), .Y(n_614) );
AND2x2_ASAP7_75t_L g670 ( .A(n_487), .B(n_522), .Y(n_670) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_493), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .C(n_492), .Y(n_489) );
INVx3_ASAP7_75t_L g532 ( .A(n_498), .Y(n_532) );
AND2x2_ASAP7_75t_L g544 ( .A(n_498), .B(n_512), .Y(n_544) );
INVx2_ASAP7_75t_L g583 ( .A(n_498), .Y(n_583) );
NOR2x1_ASAP7_75t_SL g596 ( .A(n_498), .B(n_522), .Y(n_596) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B(n_509), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_504) );
INVx1_ASAP7_75t_L g698 ( .A(n_510), .Y(n_698) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_512), .Y(n_579) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_512), .Y(n_595) );
AND2x2_ASAP7_75t_L g603 ( .A(n_512), .B(n_532), .Y(n_603) );
INVx1_ASAP7_75t_L g643 ( .A(n_512), .Y(n_643) );
INVx1_ASAP7_75t_L g668 ( .A(n_512), .Y(n_668) );
OR2x2_ASAP7_75t_L g729 ( .A(n_512), .B(n_522), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OA211x2_ASAP7_75t_L g750 ( .A1(n_520), .A2(n_751), .B(n_753), .C(n_760), .Y(n_750) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_544), .Y(n_671) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_521), .B(n_531), .Y(n_689) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g543 ( .A(n_522), .Y(n_543) );
INVx2_ASAP7_75t_L g585 ( .A(n_522), .Y(n_585) );
AND2x4_ASAP7_75t_L g648 ( .A(n_522), .B(n_605), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_522), .B(n_644), .Y(n_699) );
AND2x2_ASAP7_75t_L g742 ( .A(n_522), .B(n_583), .Y(n_742) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_531), .B(n_643), .Y(n_736) );
AND2x2_ASAP7_75t_L g756 ( .A(n_531), .B(n_579), .Y(n_756) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g644 ( .A(n_532), .Y(n_644) );
INVx1_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
NOR2xp67_ASAP7_75t_SL g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g712 ( .A(n_535), .Y(n_712) );
NOR2xp67_ASAP7_75t_L g759 ( .A(n_535), .B(n_713), .Y(n_759) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g732 ( .A(n_537), .B(n_574), .Y(n_732) );
OAI211xp5_ASAP7_75t_L g720 ( .A1(n_538), .A2(n_721), .B(n_724), .C(n_733), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g764 ( .A1(n_538), .A2(n_758), .B(n_765), .C(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g649 ( .A(n_539), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g568 ( .A(n_540), .Y(n_568) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_540), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g624 ( .A(n_540), .B(n_574), .Y(n_624) );
NOR2xp67_ASAP7_75t_L g734 ( .A(n_540), .B(n_574), .Y(n_734) );
AND2x2_ASAP7_75t_L g607 ( .A(n_541), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g658 ( .A(n_541), .Y(n_658) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x4_ASAP7_75t_SL g547 ( .A(n_543), .B(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g604 ( .A(n_543), .B(n_605), .Y(n_604) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_543), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g652 ( .A(n_543), .B(n_653), .Y(n_652) );
NOR2xp67_ASAP7_75t_SL g735 ( .A(n_543), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_544), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_SL g775 ( .A(n_544), .B(n_617), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx2_ASAP7_75t_SL g743 ( .A(n_549), .Y(n_743) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_567), .Y(n_549) );
INVx3_ASAP7_75t_L g666 ( .A(n_550), .Y(n_666) );
AND2x2_ASAP7_75t_L g687 ( .A(n_550), .B(n_678), .Y(n_687) );
AND2x2_ASAP7_75t_L g745 ( .A(n_550), .B(n_627), .Y(n_745) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g574 ( .A(n_552), .Y(n_574) );
INVx1_ASAP7_75t_L g610 ( .A(n_552), .Y(n_610) );
INVx1_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_560), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVxp67_ASAP7_75t_L g713 ( .A(n_567), .Y(n_713) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g573 ( .A(n_569), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g640 ( .A(n_569), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_577), .B1(n_580), .B2(n_586), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g587 ( .A(n_573), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g598 ( .A(n_573), .Y(n_598) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g647 ( .A(n_578), .B(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g667 ( .A(n_582), .B(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g675 ( .A(n_583), .Y(n_675) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g723 ( .A(n_585), .B(n_614), .Y(n_723) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_587), .A2(n_681), .B(n_682), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_597), .B(n_600), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g646 ( .A(n_596), .B(n_620), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_597), .A2(n_704), .B1(n_706), .B2(n_708), .Y(n_703) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_606), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_SL g653 ( .A(n_603), .Y(n_653) );
AND2x2_ASAP7_75t_L g682 ( .A(n_604), .B(n_620), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_604), .B(n_642), .Y(n_714) );
AND2x2_ASAP7_75t_L g718 ( .A(n_604), .B(n_675), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_606), .A2(n_663), .B(n_667), .Y(n_662) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
AND2x2_ASAP7_75t_L g623 ( .A(n_607), .B(n_624), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_607), .B(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g692 ( .A(n_610), .Y(n_692) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_635), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_622), .B1(n_625), .B2(n_631), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx4_ASAP7_75t_L g634 ( .A(n_614), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_614), .B(n_620), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_614), .B(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_617), .A2(n_641), .B(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g740 ( .A(n_617), .B(n_642), .Y(n_740) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g722 ( .A(n_619), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g758 ( .A(n_620), .B(n_742), .Y(n_758) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g638 ( .A(n_624), .B(n_639), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_624), .B(n_658), .Y(n_657) );
OAI22xp5_ASAP7_75t_SL g635 ( .A1(n_625), .A2(n_636), .B1(n_637), .B2(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g752 ( .A(n_629), .B(n_639), .Y(n_752) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g650 ( .A(n_630), .Y(n_650) );
AND2x2_ASAP7_75t_L g676 ( .A(n_630), .B(n_639), .Y(n_676) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_632), .B(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_633), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g727 ( .A(n_634), .Y(n_727) );
INVx1_ASAP7_75t_L g739 ( .A(n_636), .Y(n_739) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_638), .A2(n_682), .B1(n_761), .B2(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g677 ( .A(n_639), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g748 ( .A(n_639), .B(n_701), .Y(n_748) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g651 ( .A1(n_642), .A2(n_652), .B(n_654), .C(n_655), .Y(n_651) );
AND2x2_ASAP7_75t_SL g761 ( .A(n_642), .B(n_648), .Y(n_761) );
AND2x4_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_643), .Y(n_695) );
O2A1O1Ixp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_649), .C(n_651), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_673) );
INVx2_ASAP7_75t_L g654 ( .A(n_648), .Y(n_654) );
AND2x2_ASAP7_75t_L g674 ( .A(n_648), .B(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_648), .Y(n_741) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g782 ( .A(n_660), .Y(n_782) );
NOR2x1_ASAP7_75t_SL g660 ( .A(n_661), .B(n_672), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_669), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_663), .A2(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
INVx1_ASAP7_75t_L g769 ( .A(n_666), .Y(n_769) );
AND2x2_ASAP7_75t_L g707 ( .A(n_670), .B(n_695), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_671), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_680), .Y(n_672) );
AND2x2_ASAP7_75t_L g774 ( .A(n_676), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2x1_ASAP7_75t_L g683 ( .A(n_684), .B(n_719), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_703), .C(n_710), .Y(n_684) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_690), .B2(n_694), .C1(n_696), .C2(n_700), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g746 ( .A(n_705), .Y(n_746) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp67_ASAP7_75t_SL g719 ( .A(n_720), .B(n_737), .Y(n_719) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_730), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_727), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g779 ( .A(n_732), .Y(n_779) );
NAND2xp33_ASAP7_75t_SL g733 ( .A(n_734), .B(n_735), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_743), .B1(n_744), .B2(n_746), .C(n_747), .Y(n_737) );
NOR4xp25_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .C(n_741), .D(n_742), .Y(n_738) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_749), .A2(n_782), .B(n_783), .Y(n_781) );
NAND4xp75_ASAP7_75t_L g749 ( .A(n_750), .B(n_764), .C(n_770), .D(n_776), .Y(n_749) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_759), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_771), .B(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_787), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_796), .B(n_797), .Y(n_789) );
INVxp33_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2x1_ASAP7_75t_SL g791 ( .A(n_792), .B(n_795), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
OR3x1_ASAP7_75t_L g797 ( .A(n_798), .B(n_805), .C(n_809), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_798), .A2(n_813), .B(n_816), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_R g815 ( .A(n_804), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_827), .Y(n_811) );
INVx1_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_822), .B1(n_823), .B2(n_826), .Y(n_818) );
INVx1_ASAP7_75t_L g826 ( .A(n_819), .Y(n_826) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
CKINVDCx11_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
CKINVDCx8_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
endmodule