module fake_ariane_611_n_1106 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_122, n_268, n_257, n_266, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1106);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1106;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_1016;
wire n_346;
wire n_940;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_597;
wire n_1018;
wire n_816;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_1099;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_449;
wire n_333;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_20),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_180),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_39),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_68),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_31),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_2),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_213),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_170),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_67),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_45),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_215),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_126),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_164),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_139),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_169),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_138),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_125),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_42),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_121),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_187),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_56),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_74),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_192),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_104),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_233),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_168),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_23),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_136),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_7),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_265),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_35),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_166),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_153),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_97),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_30),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_244),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_149),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_134),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_61),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_9),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_113),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_177),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_144),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_29),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_47),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_24),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_42),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_124),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_76),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_120),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_48),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_280),
.B(n_0),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_302),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_0),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_302),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_304),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_280),
.B(n_1),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_278),
.B(n_1),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_304),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_330),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_273),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_283),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_281),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_277),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_283),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_293),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_328),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_287),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_295),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_2),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_300),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_312),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_314),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_3),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_318),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_322),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_325),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_315),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_R g379 ( 
.A(n_274),
.B(n_46),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_341),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_315),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_341),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

CKINVDCx8_ASAP7_75t_R g389 ( 
.A(n_343),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_347),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_316),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_368),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_316),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_344),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_344),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_332),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_323),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_352),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_352),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_366),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_290),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_348),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_353),
.B(n_324),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_R g424 ( 
.A(n_365),
.B(n_275),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_365),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_348),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_357),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_428),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_359),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_424),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_327),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_411),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_373),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_334),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_416),
.A2(n_370),
.B1(n_336),
.B2(n_368),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_375),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_394),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_425),
.B(n_377),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_336),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_370),
.Y(n_449)
);

INVx4_ASAP7_75t_SL g450 ( 
.A(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_301),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_394),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_426),
.A2(n_328),
.B1(n_335),
.B2(n_279),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_426),
.A2(n_416),
.B1(n_422),
.B2(n_419),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_393),
.B(n_285),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_394),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_276),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_3),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_422),
.B(n_284),
.C(n_282),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_396),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_L g471 ( 
.A(n_408),
.B(n_379),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_421),
.B(n_288),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_421),
.B(n_289),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_383),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_399),
.A2(n_285),
.B1(n_292),
.B2(n_291),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_407),
.B(n_296),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_285),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g480 ( 
.A(n_408),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_413),
.B(n_285),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_398),
.B(n_4),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_412),
.B(n_4),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_397),
.B(n_5),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_299),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_420),
.B(n_305),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_382),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_382),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_412),
.A2(n_308),
.B1(n_311),
.B2(n_306),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_452),
.B(n_395),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_470),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_435),
.A2(n_440),
.B(n_475),
.C(n_451),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_456),
.A2(n_387),
.B1(n_400),
.B2(n_386),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_395),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_442),
.A2(n_415),
.B1(n_414),
.B2(n_393),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_439),
.B(n_402),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_453),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_414),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_445),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_461),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_415),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_475),
.B(n_313),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_454),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_462),
.B(n_317),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_458),
.B(n_406),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_464),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_463),
.B(n_389),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_442),
.A2(n_409),
.B(n_423),
.C(n_320),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_462),
.B(n_319),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_466),
.A2(n_423),
.B1(n_403),
.B2(n_427),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_457),
.B(n_389),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_477),
.C(n_455),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_468),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_434),
.B(n_326),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_463),
.B(n_5),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_6),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_446),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_333),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_458),
.B(n_392),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_474),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_487),
.B(n_418),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_6),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_403),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_7),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_457),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_459),
.B(n_8),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_435),
.B(n_8),
.Y(n_537)
);

BUFx6f_ASAP7_75t_SL g538 ( 
.A(n_432),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_440),
.B(n_9),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_459),
.B(n_10),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_485),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_480),
.B(n_10),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_476),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_448),
.B(n_11),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_480),
.B(n_11),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_436),
.B(n_12),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_487),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_432),
.B(n_13),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_444),
.B(n_15),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_447),
.B(n_15),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_481),
.B(n_16),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_469),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_486),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_448),
.B(n_16),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_481),
.B(n_17),
.Y(n_559)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_471),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_491),
.B(n_18),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_472),
.B(n_19),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_486),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_483),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_477),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_436),
.B(n_21),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_495),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_507),
.B(n_488),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_498),
.A2(n_490),
.B(n_479),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_502),
.B(n_494),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_504),
.B(n_496),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_521),
.B(n_479),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_504),
.B(n_450),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_500),
.B(n_450),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_497),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_503),
.A2(n_484),
.B(n_491),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_L g578 ( 
.A1(n_562),
.A2(n_473),
.B(n_484),
.C(n_467),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_505),
.Y(n_579)
);

BUFx8_ASAP7_75t_SL g580 ( 
.A(n_506),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_516),
.B(n_450),
.Y(n_581)
);

AO21x1_ASAP7_75t_L g582 ( 
.A1(n_554),
.A2(n_478),
.B(n_482),
.Y(n_582)
);

AO21x1_ASAP7_75t_L g583 ( 
.A1(n_554),
.A2(n_491),
.B(n_50),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_499),
.B(n_22),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_509),
.A2(n_51),
.B(n_49),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_512),
.A2(n_518),
.B(n_526),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_527),
.A2(n_53),
.B(n_52),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_516),
.B(n_23),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_530),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_510),
.B(n_24),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_559),
.A2(n_55),
.B(n_54),
.Y(n_591)
);

NOR3xp33_ASAP7_75t_L g592 ( 
.A(n_549),
.B(n_25),
.C(n_26),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_520),
.B(n_25),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_531),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_540),
.A2(n_58),
.B(n_57),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_520),
.B(n_26),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_545),
.A2(n_558),
.B(n_539),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_515),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_537),
.A2(n_27),
.B(n_28),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_522),
.B(n_27),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_557),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_529),
.B(n_31),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_535),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_538),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_563),
.Y(n_605)
);

NAND2x1p5_ASAP7_75t_L g606 ( 
.A(n_534),
.B(n_59),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_501),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_566),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_508),
.B(n_36),
.Y(n_609)
);

NOR2x1_ASAP7_75t_L g610 ( 
.A(n_520),
.B(n_36),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_511),
.A2(n_62),
.B(n_60),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_552),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_552),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_566),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_553),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_567),
.B(n_44),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_541),
.Y(n_621)
);

NOR2x1p5_ASAP7_75t_SL g622 ( 
.A(n_542),
.B(n_63),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_567),
.B(n_45),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_525),
.B(n_64),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_514),
.A2(n_65),
.B(n_66),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_514),
.A2(n_536),
.B(n_544),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_530),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_536),
.A2(n_69),
.B(n_70),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_513),
.A2(n_71),
.B(n_72),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_553),
.A2(n_73),
.B(n_75),
.C(n_77),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_525),
.B(n_524),
.Y(n_631)
);

AO31x2_ASAP7_75t_L g632 ( 
.A1(n_582),
.A2(n_524),
.A3(n_517),
.B(n_547),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_572),
.B(n_501),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_588),
.B(n_564),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_571),
.B(n_551),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_631),
.B(n_523),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_568),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_584),
.A2(n_519),
.B(n_560),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_586),
.A2(n_546),
.B(n_543),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_579),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_612),
.A2(n_561),
.B(n_546),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_627),
.B(n_528),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_624),
.A2(n_543),
.B(n_561),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_597),
.A2(n_548),
.B(n_565),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_574),
.A2(n_538),
.B(n_532),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_598),
.B(n_519),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_603),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_577),
.A2(n_570),
.B(n_626),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_591),
.A2(n_78),
.B(n_79),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_569),
.B(n_80),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_578),
.A2(n_81),
.B(n_82),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_610),
.B(n_83),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_609),
.A2(n_84),
.B(n_85),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_614),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_583),
.A2(n_86),
.B(n_87),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_621),
.B(n_88),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_581),
.A2(n_89),
.B(n_90),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_589),
.B(n_91),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_576),
.B(n_92),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_576),
.B(n_93),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_620),
.B(n_94),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_595),
.A2(n_95),
.B(n_96),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_575),
.A2(n_98),
.B(n_99),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_573),
.A2(n_100),
.B(n_101),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_573),
.A2(n_102),
.B(n_103),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_589),
.B(n_105),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_590),
.A2(n_106),
.B(n_107),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_587),
.A2(n_108),
.B(n_109),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_585),
.A2(n_625),
.B(n_628),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_623),
.B(n_110),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_600),
.A2(n_111),
.B(n_112),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_594),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_608),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_629),
.A2(n_117),
.B(n_118),
.Y(n_675)
);

AOI21xp33_ASAP7_75t_L g676 ( 
.A1(n_605),
.A2(n_119),
.B(n_122),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_594),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_615),
.Y(n_678)
);

AO31x2_ASAP7_75t_L g679 ( 
.A1(n_608),
.A2(n_123),
.A3(n_127),
.B(n_128),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_593),
.B(n_129),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_580),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_606),
.A2(n_130),
.B(n_131),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_132),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_619),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_606),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_602),
.A2(n_133),
.B(n_135),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_596),
.B(n_137),
.Y(n_687)
);

AO31x2_ASAP7_75t_L g688 ( 
.A1(n_617),
.A2(n_140),
.A3(n_141),
.B(n_142),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_604),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_611),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_599),
.A2(n_143),
.B(n_145),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_617),
.A2(n_146),
.A3(n_147),
.B(n_150),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_637),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_633),
.A2(n_607),
.B1(n_618),
.B2(n_599),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_646),
.B(n_635),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_640),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_647),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_643),
.A2(n_630),
.A3(n_616),
.B(n_613),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_654),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_638),
.A2(n_601),
.B1(n_611),
.B2(n_592),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_680),
.B(n_151),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_SL g702 ( 
.A1(n_639),
.A2(n_622),
.B(n_154),
.C(n_155),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_634),
.A2(n_152),
.B(n_156),
.C(n_157),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_647),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_636),
.A2(n_158),
.B(n_159),
.C(n_160),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_678),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_680),
.B(n_161),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_678),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_681),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_690),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_642),
.B(n_272),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_657),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_670),
.A2(n_162),
.B(n_163),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_642),
.A2(n_165),
.B1(n_167),
.B2(n_171),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_657),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_657),
.B(n_172),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_662),
.A2(n_173),
.B(n_174),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_650),
.B(n_175),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_673),
.B(n_271),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_684),
.B(n_176),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_673),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_645),
.B(n_673),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_671),
.A2(n_178),
.B(n_179),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_685),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_677),
.B(n_181),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_651),
.A2(n_182),
.B(n_183),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_677),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_644),
.A2(n_184),
.B(n_185),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_677),
.B(n_186),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_685),
.B(n_270),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_687),
.B(n_188),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_667),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_656),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_660),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_661),
.B(n_189),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_689),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_648),
.A2(n_190),
.B(n_191),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_632),
.B(n_193),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_652),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_683),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_652),
.B(n_194),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_659),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_693),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_697),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_696),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_700),
.A2(n_674),
.B1(n_672),
.B2(n_668),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_738),
.A2(n_641),
.B(n_691),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_694),
.A2(n_739),
.B1(n_695),
.B2(n_714),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_736),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_SL g750 ( 
.A1(n_694),
.A2(n_652),
.B1(n_653),
.B2(n_666),
.Y(n_750)
);

AO21x1_ASAP7_75t_L g751 ( 
.A1(n_718),
.A2(n_665),
.B(n_676),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_707),
.A2(n_658),
.B1(n_655),
.B2(n_664),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_704),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_706),
.Y(n_754)
);

OA21x2_ASAP7_75t_L g755 ( 
.A1(n_738),
.A2(n_686),
.B(n_669),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_708),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_710),
.B(n_652),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_732),
.A2(n_682),
.B1(n_688),
.B2(n_692),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_709),
.Y(n_760)
);

INVxp33_ASAP7_75t_SL g761 ( 
.A(n_701),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_727),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_710),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_722),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_739),
.A2(n_692),
.B1(n_688),
.B2(n_679),
.Y(n_765)
);

CKINVDCx8_ASAP7_75t_R g766 ( 
.A(n_715),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_722),
.B(n_679),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_721),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_712),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_722),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_715),
.B(n_679),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_711),
.A2(n_663),
.B1(n_649),
.B2(n_675),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_741),
.A2(n_692),
.B1(n_688),
.B2(n_197),
.Y(n_773)
);

AO21x1_ASAP7_75t_SL g774 ( 
.A1(n_741),
.A2(n_195),
.B(n_196),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_715),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_716),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_716),
.Y(n_777)
);

INVx6_ASAP7_75t_L g778 ( 
.A(n_730),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_724),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_733),
.A2(n_269),
.B1(n_200),
.B2(n_201),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_724),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_725),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_698),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_713),
.A2(n_198),
.B(n_202),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_728),
.A2(n_203),
.B(n_204),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_740),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_730),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_720),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_742),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_719),
.B(n_208),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_734),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_734),
.A2(n_268),
.B1(n_214),
.B2(n_216),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_719),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_742),
.A2(n_212),
.B1(n_217),
.B2(n_218),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_731),
.A2(n_266),
.B1(n_220),
.B2(n_221),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_729),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_729),
.Y(n_797)
);

CKINVDCx11_ASAP7_75t_R g798 ( 
.A(n_702),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_698),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_698),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_735),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_703),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_717),
.B(n_219),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_705),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_776),
.B(n_723),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_800),
.B(n_737),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_768),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_744),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_783),
.B(n_726),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_762),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_753),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_770),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_799),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_764),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_764),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_746),
.A2(n_222),
.B(n_223),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_747),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_747),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_745),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_804),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_767),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_767),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_771),
.B(n_224),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_767),
.B(n_225),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_747),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_754),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_765),
.A2(n_226),
.B(n_227),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_756),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_777),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_755),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_779),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_779),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_755),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_758),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_797),
.B(n_228),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_755),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_786),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_787),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_786),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_781),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_769),
.B(n_229),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_765),
.B(n_230),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_788),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_759),
.A2(n_231),
.B(n_232),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_784),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_748),
.B(n_234),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_784),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_773),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_793),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_759),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_782),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_796),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_757),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_812),
.B(n_750),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_823),
.B(n_824),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_807),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_812),
.B(n_763),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_808),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_818),
.B(n_763),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_818),
.B(n_821),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

OAI221xp5_ASAP7_75t_L g864 ( 
.A1(n_850),
.A2(n_802),
.B1(n_787),
.B2(n_780),
.C(n_792),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_808),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_823),
.B(n_824),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_831),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_853),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_810),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_821),
.B(n_749),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_855),
.B(n_749),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_835),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_855),
.B(n_801),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_842),
.B(n_774),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_831),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_848),
.B(n_795),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_842),
.B(n_797),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

INVx3_ASAP7_75t_SL g879 ( 
.A(n_822),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_839),
.Y(n_880)
);

AOI221x1_ASAP7_75t_L g881 ( 
.A1(n_817),
.A2(n_752),
.B1(n_803),
.B2(n_790),
.C(n_751),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_845),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_842),
.B(n_775),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_845),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_839),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_840),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_828),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_852),
.B(n_802),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_853),
.B(n_761),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_817),
.B(n_780),
.C(n_792),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_852),
.B(n_811),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_833),
.B(n_772),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_820),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_841),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_848),
.A2(n_791),
.B(n_795),
.C(n_761),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_833),
.B(n_834),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_814),
.B(n_834),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_814),
.B(n_815),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_828),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_814),
.B(n_791),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_841),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_840),
.B(n_778),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_836),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_841),
.Y(n_904)
);

OAI221xp5_ASAP7_75t_L g905 ( 
.A1(n_850),
.A2(n_778),
.B1(n_766),
.B2(n_785),
.C(n_798),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_820),
.B(n_778),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_854),
.B(n_766),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_R g908 ( 
.A(n_843),
.B(n_760),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_805),
.B(n_794),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_876),
.B(n_805),
.C(n_844),
.Y(n_910)
);

OA21x2_ASAP7_75t_L g911 ( 
.A1(n_881),
.A2(n_838),
.B(n_835),
.Y(n_911)
);

NAND4xp25_ASAP7_75t_SL g912 ( 
.A(n_895),
.B(n_844),
.C(n_843),
.D(n_826),
.Y(n_912)
);

AOI221xp5_ASAP7_75t_L g913 ( 
.A1(n_888),
.A2(n_864),
.B1(n_890),
.B2(n_856),
.C(n_891),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_858),
.B(n_854),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_822),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_890),
.A2(n_846),
.B1(n_809),
.B2(n_837),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_909),
.A2(n_856),
.B1(n_889),
.B2(n_888),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_891),
.B(n_822),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_909),
.B(n_789),
.C(n_849),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_886),
.A2(n_846),
.B1(n_809),
.B2(n_837),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_886),
.B(n_859),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_875),
.B(n_822),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_867),
.B(n_830),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_862),
.B(n_830),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_886),
.A2(n_846),
.B1(n_837),
.B2(n_826),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_900),
.A2(n_846),
.B1(n_829),
.B2(n_798),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_902),
.A2(n_846),
.B1(n_837),
.B2(n_806),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_900),
.A2(n_829),
.B1(n_836),
.B2(n_851),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_859),
.B(n_861),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_862),
.B(n_830),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_857),
.B(n_820),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_861),
.B(n_851),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_892),
.A2(n_832),
.B(n_820),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_857),
.B(n_832),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_870),
.B(n_760),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_870),
.B(n_813),
.Y(n_936)
);

OAI221xp5_ASAP7_75t_SL g937 ( 
.A1(n_905),
.A2(n_832),
.B1(n_806),
.B2(n_825),
.C(n_838),
.Y(n_937)
);

OAI221xp5_ASAP7_75t_SL g938 ( 
.A1(n_892),
.A2(n_832),
.B1(n_825),
.B2(n_835),
.C(n_838),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_871),
.B(n_813),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_871),
.A2(n_849),
.B1(n_847),
.B2(n_813),
.Y(n_940)
);

OAI221xp5_ASAP7_75t_L g941 ( 
.A1(n_907),
.A2(n_851),
.B1(n_819),
.B2(n_827),
.C(n_849),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_882),
.B(n_819),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_882),
.B(n_819),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_884),
.B(n_827),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_879),
.A2(n_849),
.B1(n_847),
.B2(n_827),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_884),
.B(n_815),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_857),
.B(n_847),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_931),
.B(n_906),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_931),
.B(n_906),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_942),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_911),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_923),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_924),
.B(n_930),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_934),
.B(n_866),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_914),
.B(n_897),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_943),
.Y(n_956)
);

NAND2x1p5_ASAP7_75t_L g957 ( 
.A(n_911),
.B(n_829),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_934),
.B(n_921),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_932),
.B(n_897),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_944),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_917),
.B(n_873),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_946),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_911),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_922),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_947),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_929),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_941),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_857),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_938),
.B(n_866),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_910),
.B(n_873),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_936),
.B(n_874),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_939),
.B(n_866),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_935),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_918),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_915),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_913),
.B(n_883),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_971),
.Y(n_977)
);

NOR2x1p5_ASAP7_75t_L g978 ( 
.A(n_973),
.B(n_893),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_973),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_955),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_952),
.B(n_919),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_955),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_935),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_956),
.B(n_887),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_953),
.B(n_916),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_954),
.B(n_965),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_962),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_971),
.B(n_933),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_953),
.B(n_866),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_954),
.B(n_879),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_962),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_959),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_979),
.B(n_981),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_978),
.B(n_965),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_983),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_986),
.B(n_965),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_986),
.B(n_958),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_980),
.B(n_967),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_983),
.B(n_958),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_990),
.B(n_968),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_990),
.B(n_968),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_982),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_992),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_985),
.B(n_970),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_984),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_993),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1002),
.B(n_987),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_1004),
.A2(n_967),
.B1(n_926),
.B2(n_957),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_998),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_993),
.B(n_991),
.Y(n_1012)
);

AND2x4_ASAP7_75t_SL g1013 ( 
.A(n_995),
.B(n_986),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_SL g1014 ( 
.A1(n_1006),
.A2(n_995),
.B(n_994),
.Y(n_1014)
);

AOI21xp33_ASAP7_75t_SL g1015 ( 
.A1(n_1012),
.A2(n_994),
.B(n_977),
.Y(n_1015)
);

AOI32xp33_ASAP7_75t_L g1016 ( 
.A1(n_1009),
.A2(n_963),
.A3(n_951),
.B1(n_920),
.B2(n_925),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1007),
.A2(n_969),
.B1(n_997),
.B2(n_999),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1011),
.B(n_997),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1018),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_1014),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1017),
.B(n_1007),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_1015),
.B(n_1013),
.Y(n_1022)
);

AOI222xp33_ASAP7_75t_L g1023 ( 
.A1(n_1016),
.A2(n_951),
.B1(n_963),
.B2(n_1010),
.C1(n_976),
.C2(n_926),
.Y(n_1023)
);

AOI211xp5_ASAP7_75t_L g1024 ( 
.A1(n_1021),
.A2(n_1008),
.B(n_927),
.C(n_912),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1023),
.A2(n_957),
.B1(n_988),
.B2(n_977),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_1020),
.B(n_996),
.Y(n_1026)
);

AOI22x1_ASAP7_75t_L g1027 ( 
.A1(n_1020),
.A2(n_996),
.B1(n_988),
.B2(n_1000),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1019),
.B(n_1022),
.Y(n_1028)
);

OAI211xp5_ASAP7_75t_L g1029 ( 
.A1(n_1020),
.A2(n_881),
.B(n_908),
.C(n_1001),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_L g1030 ( 
.A(n_1020),
.B(n_937),
.C(n_969),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_1024),
.A2(n_1029),
.B1(n_1030),
.B2(n_1026),
.Y(n_1031)
);

AOI211xp5_ASAP7_75t_L g1032 ( 
.A1(n_1028),
.A2(n_961),
.B(n_940),
.C(n_945),
.Y(n_1032)
);

NAND4xp25_ASAP7_75t_L g1033 ( 
.A(n_1025),
.B(n_975),
.C(n_964),
.D(n_974),
.Y(n_1033)
);

NOR4xp25_ASAP7_75t_L g1034 ( 
.A(n_1027),
.B(n_975),
.C(n_964),
.D(n_960),
.Y(n_1034)
);

AND3x1_ASAP7_75t_L g1035 ( 
.A(n_1026),
.B(n_974),
.C(n_972),
.Y(n_1035)
);

AOI211xp5_ASAP7_75t_L g1036 ( 
.A1(n_1029),
.A2(n_874),
.B(n_879),
.C(n_989),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_SL g1037 ( 
.A(n_1034),
.B(n_957),
.C(n_966),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_950),
.C(n_960),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_L g1039 ( 
.A(n_1033),
.B(n_950),
.C(n_887),
.Y(n_1039)
);

XNOR2xp5_ASAP7_75t_L g1040 ( 
.A(n_1035),
.B(n_928),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_1036),
.B(n_899),
.C(n_903),
.Y(n_1041)
);

NAND4xp25_ASAP7_75t_SL g1042 ( 
.A(n_1032),
.B(n_949),
.C(n_948),
.D(n_972),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1034),
.B(n_959),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_L g1044 ( 
.A(n_1031),
.B(n_954),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1040),
.A2(n_928),
.B1(n_948),
.B2(n_949),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_1044),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_1043),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1037),
.A2(n_903),
.B1(n_899),
.B2(n_847),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1038),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1041),
.A2(n_883),
.B1(n_877),
.B2(n_872),
.Y(n_1050)
);

AO22x1_ASAP7_75t_L g1051 ( 
.A1(n_1039),
.A2(n_877),
.B1(n_860),
.B2(n_865),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1042),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_878),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1044),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1044),
.B(n_878),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_1040),
.A2(n_872),
.B1(n_860),
.B2(n_869),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1044),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1044),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1044),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1049),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_1054),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1057),
.Y(n_1062)
);

OAI211xp5_ASAP7_75t_L g1063 ( 
.A1(n_1058),
.A2(n_869),
.B(n_865),
.C(n_872),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_1059),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1047),
.Y(n_1065)
);

OAI21xp33_ASAP7_75t_SL g1066 ( 
.A1(n_1046),
.A2(n_896),
.B(n_898),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1053),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_1052),
.B(n_896),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1055),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1051),
.B(n_898),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_1048),
.Y(n_1071)
);

NAND4xp75_ASAP7_75t_L g1072 ( 
.A(n_1056),
.B(n_236),
.C(n_238),
.D(n_239),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_1045),
.B(n_904),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1050),
.Y(n_1074)
);

NAND4xp75_ASAP7_75t_L g1075 ( 
.A(n_1057),
.B(n_241),
.C(n_242),
.D(n_243),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1057),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_1065),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1061),
.Y(n_1078)
);

NAND3x1_ASAP7_75t_L g1079 ( 
.A(n_1062),
.B(n_246),
.C(n_247),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1075),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1064),
.B(n_880),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1076),
.A2(n_904),
.B(n_901),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1060),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_1060),
.B(n_249),
.Y(n_1084)
);

NOR2x1p5_ASAP7_75t_L g1085 ( 
.A(n_1069),
.B(n_250),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1068),
.B(n_901),
.Y(n_1086)
);

NOR2x1p5_ASAP7_75t_L g1087 ( 
.A(n_1078),
.B(n_1067),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1083),
.B(n_1071),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1077),
.A2(n_1068),
.B1(n_1074),
.B2(n_1066),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_1084),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1085),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1081),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_1088),
.B(n_1080),
.C(n_1072),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1091),
.A2(n_1090),
.B1(n_1089),
.B2(n_1092),
.C(n_1063),
.Y(n_1094)
);

OAI221xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1087),
.A2(n_1070),
.B1(n_1086),
.B2(n_1082),
.C(n_1079),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_SL g1096 ( 
.A(n_1090),
.B(n_1073),
.C(n_252),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1093),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1097),
.A2(n_1094),
.B(n_1095),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1097),
.B(n_1096),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1098),
.A2(n_1073),
.B1(n_894),
.B2(n_885),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_SL g1101 ( 
.A1(n_1099),
.A2(n_251),
.B(n_253),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1101),
.A2(n_255),
.B(n_256),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1100),
.A2(n_894),
.B1(n_885),
.B2(n_880),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_SL g1104 ( 
.A1(n_1102),
.A2(n_863),
.B1(n_816),
.B2(n_815),
.Y(n_1104)
);

OAI221xp5_ASAP7_75t_R g1105 ( 
.A1(n_1104),
.A2(n_1103),
.B1(n_258),
.B2(n_259),
.C(n_260),
.Y(n_1105)
);

AOI211xp5_ASAP7_75t_L g1106 ( 
.A1(n_1105),
.A2(n_257),
.B(n_262),
.C(n_264),
.Y(n_1106)
);


endmodule