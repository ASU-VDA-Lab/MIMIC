module fake_jpeg_17248_n_158 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_1),
.C(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_38),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_34),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_3),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_16),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_44),
.B1(n_21),
.B2(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_4),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_22),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_16),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_48),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_50),
.Y(n_77)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_76),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_73),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_22),
.B1(n_26),
.B2(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_40),
.B1(n_47),
.B2(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_46),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_92),
.B1(n_59),
.B2(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_97),
.C(n_96),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_63),
.B1(n_51),
.B2(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_96),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_63),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_98),
.C(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_80),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_65),
.C(n_71),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_61),
.B(n_55),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_116),
.B(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_111),
.B1(n_85),
.B2(n_84),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_55),
.C(n_54),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_114),
.C(n_115),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_59),
.B1(n_69),
.B2(n_68),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_79),
.B1(n_91),
.B2(n_83),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_54),
.C(n_68),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_54),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_100),
.Y(n_132)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_90),
.B1(n_98),
.B2(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_86),
.B1(n_90),
.B2(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_138),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_105),
.A3(n_86),
.B1(n_106),
.B2(n_109),
.C(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_88),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_85),
.B1(n_122),
.B2(n_130),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_127),
.B1(n_119),
.B2(n_124),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_120),
.C(n_128),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.C(n_132),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_120),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_149),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_151),
.B(n_144),
.Y(n_154)
);

OAI211xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_142),
.B(n_145),
.C(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

OAI221xp5_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_153),
.B1(n_142),
.B2(n_149),
.C(n_143),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_156),
.Y(n_158)
);


endmodule