module real_jpeg_12845_n_17 (n_5, n_4, n_8, n_0, n_12, n_299, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_299;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_288;
wire n_176;
wire n_292;
wire n_221;
wire n_215;
wire n_249;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_184;
wire n_48;
wire n_164;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx10_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_42),
.B1(n_61),
.B2(n_62),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_104),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_104),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_104),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_34),
.B1(n_61),
.B2(n_62),
.Y(n_76)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_11),
.B(n_142),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_44),
.B(n_82),
.C(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_11),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_11),
.B(n_38),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_156),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_29),
.C(n_65),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_83),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_11),
.A2(n_95),
.B(n_204),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_156),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_12),
.B(n_45),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_13),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_136),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_136),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_136),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_184)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_16),
.A2(n_44),
.B1(n_45),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_16),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_85),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_125),
.B1(n_295),
.B2(n_296),
.Y(n_18)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_19),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_107),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_21),
.B(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_89),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_22),
.A2(n_23),
.B1(n_73),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_56),
.B2(n_72),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B1(n_36),
.B2(n_55),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_26),
.A2(n_36),
.B(n_72),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_26),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_27),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_27),
.A2(n_31),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_27),
.A2(n_31),
.B1(n_94),
.B2(n_184),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_28),
.A2(n_29),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_28),
.B(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_31),
.B(n_159),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_33),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_43),
.B(n_48),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_37),
.A2(n_43),
.B1(n_50),
.B2(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_39),
.A2(n_50),
.B(n_156),
.C(n_165),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_39),
.A2(n_44),
.A3(n_47),
.B1(n_166),
.B2(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_43),
.B(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_43),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_43),
.A2(n_48),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_43),
.A2(n_50),
.B1(n_103),
.B2(n_253),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_50),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_68),
.B2(n_71),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_63),
.B1(n_71),
.B2(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_62),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_61),
.B(n_194),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_62),
.A2(n_81),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_71),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_63),
.B(n_151),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_63),
.A2(n_71),
.B1(n_149),
.B2(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_63),
.A2(n_71),
.B1(n_99),
.B2(n_172),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_67),
.A2(n_171),
.B(n_173),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_67),
.A2(n_173),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_67),
.B(n_156),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_71),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_73),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_88),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_75),
.A2(n_150),
.B(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_78),
.A2(n_86),
.B1(n_135),
.B2(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_78),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_78),
.A2(n_169),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_83),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_83),
.B(n_138),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_86),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_86),
.A2(n_101),
.B(n_137),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

FAx1_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_108),
.CI(n_109),
.CON(n_107),
.SN(n_107)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_89),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.C(n_102),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_90),
.A2(n_91),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_92),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_96),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_95),
.A2(n_96),
.B1(n_146),
.B2(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_95),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_145),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_96),
.A2(n_158),
.B(n_209),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_96),
.B(n_156),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_100),
.B(n_102),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_106),
.B(n_164),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_107),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_125),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_289),
.B(n_294),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_277),
.B(n_288),
.Y(n_127)
);

OAI321xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_245),
.A3(n_270),
.B1(n_275),
.B2(n_276),
.C(n_299),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_185),
.B(n_244),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_160),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_131),
.B(n_160),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_147),
.C(n_152),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_132),
.A2(n_133),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_140),
.C(n_144),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_147),
.A2(n_152),
.B1(n_153),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_154),
.B(n_157),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_175),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_161),
.B(n_176),
.C(n_177),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_174),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_162),
.B(n_168),
.C(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_178),
.B(n_182),
.Y(n_255)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_237),
.B(n_243),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_224),
.B(n_236),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_205),
.B(n_223),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_189),
.B(n_195),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_203),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_213),
.B(n_222),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_211),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_217),
.B(n_221),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_226),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_232),
.C(n_235),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_260),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_260),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_256),
.C(n_259),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_247),
.A2(n_248),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_254),
.C(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_269),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_264),
.C(n_269),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_287),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);


endmodule