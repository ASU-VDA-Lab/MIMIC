module fake_jpeg_3213_n_195 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_69),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_59),
.B1(n_48),
.B2(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_59),
.B1(n_53),
.B2(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_64),
.B1(n_57),
.B2(n_56),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_52),
.B1(n_55),
.B2(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_100),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_101),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_54),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_63),
.C(n_60),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_48),
.C(n_51),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_69),
.B(n_67),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_47),
.B(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_75),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_49),
.B1(n_52),
.B2(n_75),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_75),
.B1(n_62),
.B2(n_44),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_120),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_101),
.B(n_106),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_11),
.B(n_12),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_64),
.B1(n_56),
.B2(n_63),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_62),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_60),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_6),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_105),
.B1(n_93),
.B2(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_66),
.B1(n_61),
.B2(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_1),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_2),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_5),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_58),
.B1(n_26),
.B2(n_27),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_2),
.CI(n_3),
.CON(n_128),
.SN(n_128)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_58),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_136),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_141),
.Y(n_159)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_115),
.A3(n_128),
.B1(n_119),
.B2(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_145),
.Y(n_166)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_25),
.B1(n_42),
.B2(n_39),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_152),
.B(n_16),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_148),
.B(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_19),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_158),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_18),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_24),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_20),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_151),
.B1(n_144),
.B2(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_150),
.A3(n_151),
.B1(n_132),
.B2(n_139),
.C1(n_130),
.C2(n_34),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_21),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_176),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

FAx1_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_155),
.CI(n_165),
.CON(n_179),
.SN(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_181),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_166),
.B(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_167),
.B1(n_154),
.B2(n_157),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_186),
.C(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_175),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_177),
.Y(n_187)
);

OAI21x1_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_178),
.B(n_182),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_188),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_174),
.C(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_29),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_32),
.Y(n_195)
);


endmodule