module fake_jpeg_20915_n_156 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_76),
.B1(n_74),
.B2(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_82),
.B1(n_56),
.B2(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_67),
.B1(n_65),
.B2(n_68),
.Y(n_85)
);

BUFx6f_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_88),
.B1(n_58),
.B2(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_52),
.B1(n_69),
.B2(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_62),
.B1(n_57),
.B2(n_69),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_94),
.B1(n_66),
.B2(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_62),
.B1(n_57),
.B2(n_71),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_60),
.B1(n_53),
.B2(n_51),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_61),
.B1(n_73),
.B2(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_103),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_5),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_11),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_3),
.B(n_5),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_111),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_25),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_113),
.B1(n_18),
.B2(n_19),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_29),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_121),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_10),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_130),
.B(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_20),
.C(n_28),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_134),
.B1(n_30),
.B2(n_31),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_111),
.B1(n_113),
.B2(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_114),
.B1(n_124),
.B2(n_32),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_141),
.B(n_136),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_140),
.CI(n_142),
.CON(n_148),
.SN(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_145),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_148),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_127),
.C(n_131),
.Y(n_153)
);

AOI321xp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_144),
.A3(n_137),
.B1(n_40),
.B2(n_43),
.C(n_37),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_134),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_38),
.Y(n_156)
);


endmodule