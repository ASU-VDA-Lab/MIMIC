module real_jpeg_13687_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_1),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_1),
.B(n_31),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_56),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_25),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_6),
.B(n_51),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_6),
.B(n_35),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_6),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_7),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_25),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_10),
.B(n_25),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_51),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_56),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_14),
.Y(n_107)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_79),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_19),
.B(n_79),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_57),
.C(n_70),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_20),
.A2(n_21),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_39),
.C(n_48),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_29),
.C(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_27),
.B(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_36),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_36),
.B(n_115),
.Y(n_158)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.C(n_44),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_42),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_43),
.B(n_52),
.Y(n_129)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_52),
.B(n_115),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_57),
.A2(n_58),
.B1(n_70),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_69),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_66),
.C(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_62),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_70),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.C(n_76),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_71),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_76),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_95),
.B2(n_116),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_94),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_86),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_86),
.SN(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_95),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.CI(n_104),
.CON(n_95),
.SN(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_103),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_173),
.B(n_179),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_143),
.B(n_172),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_133),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_122),
.B(n_133),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_169),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.CI(n_126),
.CON(n_123),
.SN(n_123)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_142),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_139),
.C(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_166),
.B(n_171),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_156),
.B(n_165),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_160),
.B(n_164),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);


endmodule