module fake_jpeg_28316_n_120 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_16),
.B1(n_12),
.B2(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_16),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_12),
.B(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_46),
.B1(n_47),
.B2(n_19),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_13),
.B1(n_19),
.B2(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_50),
.B1(n_55),
.B2(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_29),
.B1(n_35),
.B2(n_13),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_44),
.B1(n_38),
.B2(n_20),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_35),
.B1(n_13),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_66),
.B1(n_56),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_35),
.B1(n_19),
.B2(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_70),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_23),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_54),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_16),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_11),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_11),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_20),
.C(n_17),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_86),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_69),
.B(n_67),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_74),
.B(n_76),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_65),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_56),
.B(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_71),
.B(n_74),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_95),
.B(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_68),
.B1(n_25),
.B2(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_77),
.C(n_82),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_88),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_22),
.B1(n_0),
.B2(n_2),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_103),
.C(n_94),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_90),
.B(n_93),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_99),
.C(n_97),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_95),
.C(n_89),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_107),
.A2(n_108),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_109),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_98),
.B1(n_96),
.B2(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

AOI31xp67_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_2),
.A3(n_3),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

AOI31xp67_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_3),
.A3(n_7),
.B(n_8),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_116),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_8),
.B(n_9),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_8),
.Y(n_120)
);


endmodule