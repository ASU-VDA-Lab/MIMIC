module fake_jpeg_5750_n_265 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_44),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_50),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_51),
.Y(n_123)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_59),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_48),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_77),
.B(n_96),
.C(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_76),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_16),
.B(n_25),
.C(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_60),
.B(n_72),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_62),
.Y(n_103)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_67),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_16),
.B1(n_17),
.B2(n_14),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_65),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_16),
.B1(n_44),
.B2(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_74),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_18),
.B1(n_29),
.B2(n_26),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_71),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_33),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_20),
.B1(n_22),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_20),
.B1(n_22),
.B2(n_27),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_37),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_89),
.Y(n_100)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_36),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_32),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_36),
.B(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_36),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_36),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_102),
.Y(n_149)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_121),
.B1(n_66),
.B2(n_82),
.Y(n_127)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_32),
.B(n_1),
.C(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_32),
.B(n_24),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_60),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_57),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_58),
.B(n_96),
.C(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_107),
.B(n_19),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_100),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_92),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_133),
.B(n_120),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_136),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_92),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_108),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_72),
.A3(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_54),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_142),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_63),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_73),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_64),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_94),
.B1(n_53),
.B2(n_62),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_154),
.B1(n_109),
.B2(n_102),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_75),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_150),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_146),
.Y(n_166)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_4),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_74),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

OAI22x1_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_55),
.B1(n_87),
.B2(n_69),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_106),
.B1(n_98),
.B2(n_118),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_55),
.B1(n_79),
.B2(n_21),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_109),
.B1(n_99),
.B2(n_113),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_21),
.B1(n_19),
.B2(n_93),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_5),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_130),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_134),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_175),
.B(n_129),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_169),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_185),
.B1(n_157),
.B2(n_128),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_126),
.B1(n_133),
.B2(n_130),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_173),
.B(n_182),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_107),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_180),
.C(n_183),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_120),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_93),
.B(n_6),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_120),
.C(n_115),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_184),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_5),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_178),
.B1(n_171),
.B2(n_177),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_203),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_201),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_136),
.B1(n_143),
.B2(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_140),
.B1(n_156),
.B2(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_198),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_147),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_175),
.C(n_180),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_99),
.B(n_6),
.C(n_7),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_174),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_206),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_129),
.C(n_6),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_7),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_217),
.B1(n_221),
.B2(n_222),
.Y(n_225)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_168),
.B1(n_171),
.B2(n_169),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_206),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_176),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_185),
.B1(n_163),
.B2(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_187),
.C(n_189),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_187),
.C(n_194),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_201),
.B1(n_195),
.B2(n_172),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_231),
.B1(n_235),
.B2(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_204),
.B1(n_192),
.B2(n_166),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_204),
.B1(n_159),
.B2(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_163),
.C(n_162),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_162),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_167),
.C(n_164),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_210),
.B1(n_226),
.B2(n_215),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_217),
.B(n_224),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_243),
.B(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_214),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_211),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_223),
.B(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_228),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_166),
.A3(n_164),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_225),
.B1(n_234),
.B2(n_227),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_237),
.B1(n_239),
.B2(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_8),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_249),
.C(n_250),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_233),
.C(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_256),
.C(n_247),
.Y(n_259)
);

XOR2x2_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_248),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_258),
.C(n_259),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_251),
.C(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_251),
.C(n_253),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_244),
.Y(n_265)
);


endmodule