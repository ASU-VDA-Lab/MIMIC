module fake_jpeg_22067_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_7),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_17),
.B1(n_35),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_64),
.B1(n_25),
.B2(n_17),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_24),
.B1(n_41),
.B2(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_35),
.B1(n_19),
.B2(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_53),
.A2(n_74),
.B1(n_24),
.B2(n_41),
.Y(n_112)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_33),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_60),
.Y(n_106)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_21),
.C(n_28),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_17),
.B1(n_19),
.B2(n_25),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_31),
.Y(n_78)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_45),
.Y(n_94)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_10),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_10),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_13),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_84),
.Y(n_120)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_51),
.Y(n_125)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_113),
.B1(n_114),
.B2(n_24),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_96),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_54),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_29),
.B(n_22),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_115),
.B(n_78),
.C(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_31),
.B1(n_23),
.B2(n_33),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_42),
.B1(n_32),
.B2(n_26),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_56),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_26),
.B1(n_32),
.B2(n_34),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_34),
.B1(n_30),
.B2(n_20),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_47),
.B(n_39),
.C(n_22),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_61),
.C(n_77),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_137),
.C(n_77),
.Y(n_158)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_121),
.Y(n_156)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_142),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_95),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_73),
.B1(n_52),
.B2(n_72),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_131),
.B(n_22),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_141),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_76),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_65),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_52),
.B1(n_74),
.B2(n_73),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_99),
.B1(n_101),
.B2(n_69),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_106),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_161),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_91),
.B(n_83),
.C(n_84),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_160),
.B1(n_165),
.B2(n_178),
.Y(n_184)
);

OR2x4_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_115),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_131),
.B(n_135),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_127),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_115),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_100),
.B(n_90),
.Y(n_204)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_163),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_167),
.C(n_118),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_114),
.B1(n_80),
.B2(n_89),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_139),
.B1(n_118),
.B2(n_81),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_88),
.B1(n_86),
.B2(n_63),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_166),
.B(n_170),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_47),
.C(n_39),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_86),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_174),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_22),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_179),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_103),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_181),
.B(n_195),
.Y(n_217)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_188),
.Y(n_221)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_152),
.B1(n_153),
.B2(n_143),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_193),
.B1(n_147),
.B2(n_177),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_197),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_204),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_138),
.B1(n_135),
.B2(n_49),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_212),
.B1(n_180),
.B2(n_163),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_47),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_155),
.B(n_174),
.C(n_147),
.D(n_149),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_155),
.C(n_162),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_67),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_30),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_22),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_213),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_151),
.A2(n_139),
.B1(n_67),
.B2(n_34),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_22),
.B(n_1),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_205),
.B1(n_3),
.B2(n_5),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_227),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_231),
.B1(n_235),
.B2(n_212),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_232),
.C(n_203),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_206),
.B(n_192),
.C(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_148),
.A3(n_20),
.B1(n_34),
.B2(n_30),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_214),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_173),
.B1(n_30),
.B2(n_20),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_173),
.B1(n_20),
.B2(n_2),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_234),
.A2(n_236),
.B1(n_186),
.B2(n_184),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_11),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_11),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_191),
.C(n_200),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_232),
.C(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_263),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_230),
.A2(n_208),
.B1(n_200),
.B2(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_190),
.B1(n_194),
.B2(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_198),
.B1(n_188),
.B2(n_207),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_261),
.A2(n_216),
.B1(n_236),
.B2(n_234),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_262),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_0),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_5),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_6),
.B(n_9),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_275),
.B1(n_253),
.B2(n_264),
.Y(n_299)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_226),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_248),
.C(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_215),
.C(n_226),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_255),
.C(n_247),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_241),
.B1(n_239),
.B2(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_245),
.B(n_9),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_288),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_261),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_243),
.Y(n_289)
);

OAI321xp33_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_280),
.A3(n_244),
.B1(n_282),
.B2(n_249),
.C(n_266),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_252),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_277),
.C(n_275),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_251),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_298),
.C(n_301),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_274),
.B1(n_278),
.B2(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_250),
.C(n_257),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_298),
.C(n_294),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_314),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_305),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_268),
.B(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_260),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_270),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_315),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_249),
.B1(n_290),
.B2(n_252),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_312),
.B1(n_308),
.B2(n_313),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_321),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_9),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_11),
.Y(n_323)
);

AOI31xp33_ASAP7_75t_SL g324 ( 
.A1(n_319),
.A2(n_304),
.A3(n_303),
.B(n_312),
.Y(n_324)
);

AOI31xp67_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_322),
.A3(n_316),
.B(n_318),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_329),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_12),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_13),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_319),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_331),
.A2(n_332),
.B(n_334),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_326),
.C(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_327),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_336),
.C(n_14),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_14),
.C(n_15),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_15),
.Y(n_340)
);


endmodule