module real_jpeg_4977_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_0),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_0),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_0),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_0),
.B(n_133),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_0),
.B(n_180),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_0),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_0),
.B(n_308),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_1),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_1),
.Y(n_185)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_1),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_1),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_2),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_2),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_3),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_3),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_3),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_4),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_4),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_4),
.B(n_185),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_4),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_4),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_4),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_4),
.B(n_142),
.Y(n_402)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_7),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_7),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_8),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_8),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_97),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_8),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_8),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_8),
.B(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_10),
.B(n_86),
.Y(n_167)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_10),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_10),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_10),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_10),
.B(n_342),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_10),
.B(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_11),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_12),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_12),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_12),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_12),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_12),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_12),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_14),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_14),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_14),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_14),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_14),
.B(n_211),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_14),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_14),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_15),
.B(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_15),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_74),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_15),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_15),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_15),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_15),
.B(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_16),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_16),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_16),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_16),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_18),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_18),
.B(n_72),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_18),
.B(n_196),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_18),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_18),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_18),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_18),
.B(n_383),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_18),
.B(n_408),
.Y(n_407)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_118),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_116),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_100),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_29),
.B(n_100),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_80),
.C(n_81),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_30),
.A2(n_31),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_53),
.C(n_69),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_32),
.A2(n_33),
.B1(n_507),
.B2(n_509),
.Y(n_506)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_37),
.C(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_39),
.Y(n_191)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_40),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_40),
.Y(n_198)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_40),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.C(n_51),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_42),
.B(n_497),
.Y(n_496)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_497)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_48),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_49),
.Y(n_355)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_50),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_50),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_50),
.Y(n_390)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_50),
.Y(n_408)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_53),
.A2(n_69),
.B1(n_70),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_53),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.C(n_64),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_54),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_56),
.Y(n_261)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_59),
.A2(n_60),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_503)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_60),
.B(n_195),
.C(n_200),
.Y(n_504)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_63),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_63),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_77),
.C(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_68),
.Y(n_212)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_68),
.Y(n_335)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_68),
.Y(n_412)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_78),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_93),
.C(n_96),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_80),
.B(n_81),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_89),
.C(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_93),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_113),
.B2(n_114),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_526),
.B(n_531),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_490),
.B(n_523),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_291),
.B(n_489),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_240),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_122),
.B(n_240),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_192),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_123),
.B(n_193),
.C(n_222),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_165),
.C(n_174),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_124),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_139),
.C(n_154),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_125),
.B(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_132),
.C(n_136),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_130),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_130),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_139),
.A2(n_140),
.B1(n_154),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_150),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_141),
.B(n_150),
.Y(n_465)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_144),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_145),
.B(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_154),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_157),
.C(n_162),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_159),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_160),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_200),
.C(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_161),
.A2(n_162),
.B1(n_200),
.B2(n_203),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_165),
.B(n_174),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_171),
.C(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_168),
.A2(n_172),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_170),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_172),
.B(n_227),
.C(n_233),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_186),
.C(n_188),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_175),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_183),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_176),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_179),
.B(n_183),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_185),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_188),
.Y(n_269)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_191),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_222),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_194),
.B(n_205),
.C(n_221),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_202),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_213),
.B1(n_220),
.B2(n_221),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.C(n_210),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_210),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_214),
.B(n_216),
.C(n_219),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_224),
.B(n_226),
.C(n_234),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_238),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.C(n_247),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_242),
.B(n_245),
.Y(n_485)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_247),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_267),
.C(n_270),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_249),
.B(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_258),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_250),
.A2(n_251),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_253),
.A2(n_254),
.B(n_257),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_253),
.B(n_258),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_433)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_264),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_265),
.B(n_368),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_270),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_282),
.C(n_287),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_272),
.B(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.C(n_279),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_273),
.B(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_275),
.A2(n_279),
.B1(n_280),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_275),
.Y(n_446)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_282),
.B(n_287),
.Y(n_467)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_483),
.B(n_488),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_470),
.B(n_482),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_452),
.B(n_469),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_426),
.B(n_451),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_394),
.B(n_425),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_360),
.B(n_393),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_337),
.B(n_359),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_315),
.B(n_336),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_312),
.B(n_314),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_310),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

INVx3_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_317),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_325),
.B2(n_326),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_328),
.C(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_323),
.Y(n_348)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_358),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_358),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_349),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_348),
.C(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_345),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_379),
.C(n_380),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_356),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_356),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_363),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_377),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_364),
.B(n_378),
.C(n_381),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_367),
.C(n_370),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_373),
.B1(n_374),
.B2(n_376),
.Y(n_370)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_371),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_376),
.Y(n_403)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g423 ( 
.A(n_382),
.B(n_388),
.C(n_391),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_388),
.B1(n_391),
.B2(n_392),
.Y(n_384)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_388),
.Y(n_392)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_424),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_424),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_405),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_404),
.C(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_403),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_399),
.Y(n_440)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_440),
.C(n_441),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_415),
.C(n_422),
.Y(n_429)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_406),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_409),
.CI(n_410),
.CON(n_406),
.SN(n_406)
);

MAJx2_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_409),
.C(n_410),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_422),
.B2(n_423),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_421),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_421),
.Y(n_436)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_449),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_449),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_438),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_430),
.C(n_438),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_461),
.C(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_443),
.C(n_448),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_447),
.B2(n_448),
.Y(n_442)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_468),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_468),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_459),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_458),
.C(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_456),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_464),
.C(n_466),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_480),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_480),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_477),
.C(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_486),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_486),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_518),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_L g523 ( 
.A1(n_491),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_511),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_492),
.B(n_511),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_500),
.B2(n_510),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_493),
.B(n_501),
.C(n_506),
.Y(n_530)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.C(n_498),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_514),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_496),
.A2(n_498),
.B1(n_499),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_500),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_506),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.C(n_505),
.Y(n_501)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_502),
.B(n_504),
.CI(n_505),
.CON(n_516),
.SN(n_516)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_507),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_516),
.C(n_517),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_512),
.A2(n_513),
.B1(n_516),
.B2(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_516),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_516),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_517),
.B(n_520),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_519),
.B(n_522),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_522),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_530),
.Y(n_531)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule