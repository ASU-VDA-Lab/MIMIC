module real_jpeg_26677_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_244;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_28),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_38),
.B1(n_43),
.B2(n_45),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_4),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_28),
.B1(n_32),
.B2(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_4),
.A2(n_52),
.B1(n_64),
.B2(n_65),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_57),
.B1(n_59),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_88),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_43),
.B1(n_45),
.B2(n_88),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_5),
.A2(n_28),
.B1(n_32),
.B2(n_88),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_6),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_61),
.B(n_65),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_57),
.B1(n_59),
.B2(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_6),
.B(n_63),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_6),
.A2(n_45),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_45),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_6),
.B(n_82),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_6),
.A2(n_26),
.B1(n_202),
.B2(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_64),
.B(n_218),
.Y(n_217)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_8),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_57),
.B1(n_59),
.B2(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_43),
.B1(n_45),
.B2(n_80),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_28),
.B1(n_32),
.B2(n_80),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_9),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_9),
.A2(n_33),
.B1(n_43),
.B2(n_45),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_10),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_10),
.A2(n_43),
.B1(n_45),
.B2(n_56),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_56),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_12),
.A2(n_57),
.B1(n_59),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_28),
.B1(n_32),
.B2(n_69),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_12),
.A2(n_43),
.B1(n_45),
.B2(n_69),
.Y(n_222)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_28),
.B1(n_32),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_15),
.Y(n_103)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_17),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_17),
.A2(n_42),
.B1(n_64),
.B2(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_17),
.A2(n_28),
.B1(n_32),
.B2(n_42),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_106),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_22),
.B(n_106),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_100),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_23),
.B(n_100),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_53),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_54),
.C(n_70),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_25),
.B(n_39),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_26),
.A2(n_34),
.B1(n_37),
.B2(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_26),
.A2(n_34),
.B(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_26),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_26),
.A2(n_36),
.B1(n_196),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_26),
.A2(n_190),
.B1(n_191),
.B2(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_27),
.A2(n_31),
.B1(n_35),
.B2(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_35),
.B1(n_96),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_27),
.A2(n_35),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_28),
.B(n_48),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_28),
.B(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_32),
.A2(n_45),
.A3(n_50),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g191 ( 
.A(n_35),
.Y(n_191)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_36),
.B(n_93),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_41),
.A2(n_112),
.B1(n_115),
.B2(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_45),
.B1(n_74),
.B2(n_77),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_43),
.A2(n_64),
.A3(n_77),
.B1(n_219),
.B2(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_45),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_46),
.A2(n_47),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_46),
.A2(n_47),
.B1(n_176),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_46),
.A2(n_47),
.B1(n_143),
.B2(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_47),
.B(n_93),
.Y(n_203)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_55),
.Y(n_90)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_67),
.B(n_93),
.C(n_94),
.Y(n_92)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_60),
.A2(n_63),
.B1(n_87),
.B2(n_140),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_73),
.Y(n_75)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_65),
.B(n_93),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_81),
.B1(n_82),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_71),
.A2(n_82),
.B1(n_138),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_76),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_72),
.A2(n_76),
.B1(n_98),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_72),
.A2(n_76),
.B1(n_158),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_77),
.Y(n_228)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.C(n_97),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_95),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_104),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_124),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_116),
.B2(n_117),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_112),
.A2(n_115),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_118),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.CI(n_123),
.CON(n_118),
.SN(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_163),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_146),
.B(n_162),
.Y(n_128)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_134),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_134),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.C(n_141),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_150),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_156),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_159),
.B(n_161),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_160),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.C(n_166),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_248),
.B(n_253),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_234),
.B(n_247),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_212),
.B(n_233),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_192),
.B(n_211),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_171),
.B(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_199),
.B(n_210),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_194),
.B(n_198),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_204),
.B(n_209),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_225),
.B1(n_231),
.B2(n_232),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_224),
.C(n_232),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_243),
.C(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);


endmodule