module fake_jpeg_25226_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx9p33_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_16),
.B1(n_25),
.B2(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_50),
.B1(n_39),
.B2(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_32),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_16),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_31),
.C(n_17),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_38),
.C(n_34),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_18),
.B(n_28),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_24),
.C(n_38),
.Y(n_81)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_29),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_63),
.Y(n_96)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_71),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_32),
.B(n_22),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_82),
.B(n_23),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_41),
.B1(n_24),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_32),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_27),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_30),
.A3(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_77),
.C(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_38),
.B(n_15),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_86),
.B1(n_101),
.B2(n_89),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_47),
.B1(n_48),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_71),
.B1(n_57),
.B2(n_80),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_65),
.B(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_60),
.C(n_62),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_108),
.C(n_118),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_78),
.B1(n_84),
.B2(n_56),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_95),
.C(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_115),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_116),
.B(n_56),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_58),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_100),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_77),
.C(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_63),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_119),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_101),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_67),
.C(n_63),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_88),
.C(n_84),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_102),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_134),
.C(n_67),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_132),
.B1(n_113),
.B2(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_91),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_103),
.C(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_135),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_92),
.B1(n_85),
.B2(n_88),
.C(n_87),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_111),
.B1(n_78),
.B2(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_131),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_78),
.B1(n_107),
.B2(n_105),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_118),
.B(n_109),
.C(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_146),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.C(n_130),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_67),
.C(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_156),
.C(n_143),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_153),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_127),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_124),
.C(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_158),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_148),
.C(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_133),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.C(n_4),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_143),
.C(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_124),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_123),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_162),
.A2(n_154),
.B(n_157),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_170),
.B(n_8),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_169),
.C(n_159),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.C(n_174),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_14),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_10),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_9),
.C(n_11),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_9),
.B(n_11),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_13),
.Y(n_177)
);


endmodule