module fake_jpeg_30740_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_63),
.Y(n_107)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_18),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_70),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_65),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_73),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_77),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_16),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_84),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_94),
.Y(n_115)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_29),
.B(n_15),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_101),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_25),
.C(n_37),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_111),
.B(n_44),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_117),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_31),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_131),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_90),
.B(n_38),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_126),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_49),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_38),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_33),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_32),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_132),
.B(n_135),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_32),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_48),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_136),
.B(n_138),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_49),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_48),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_141),
.B(n_142),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_55),
.B(n_47),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_54),
.B(n_47),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_158),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_77),
.B(n_40),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_40),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_77),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_30),
.Y(n_202)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_164),
.Y(n_228)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_166),
.Y(n_236)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_169),
.B(n_173),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_102),
.A2(n_46),
.B(n_89),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_171),
.B(n_181),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_97),
.B1(n_46),
.B2(n_57),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_194),
.B1(n_195),
.B2(n_199),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_105),
.B(n_87),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_134),
.A2(n_64),
.B1(n_68),
.B2(n_56),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_183),
.A2(n_212),
.B1(n_217),
.B2(n_113),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_112),
.A2(n_45),
.B(n_84),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_215),
.C(n_155),
.Y(n_244)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_191),
.Y(n_272)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_111),
.A2(n_34),
.B(n_45),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_37),
.B(n_113),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_134),
.A2(n_46),
.B1(n_27),
.B2(n_61),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_140),
.A2(n_89),
.B1(n_84),
.B2(n_58),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx5_ASAP7_75t_SL g197 ( 
.A(n_162),
.Y(n_197)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_151),
.A2(n_118),
.B1(n_106),
.B2(n_127),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_28),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_200),
.B(n_209),
.Y(n_242)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_201),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_202),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_30),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_206),
.B(n_208),
.Y(n_238)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

CKINVDCx12_ASAP7_75t_R g208 ( 
.A(n_162),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_125),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_28),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_220),
.B1(n_222),
.B2(n_160),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_59),
.B1(n_72),
.B2(n_76),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_34),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_213),
.B(n_219),
.Y(n_261)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_143),
.A2(n_101),
.B1(n_98),
.B2(n_95),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_154),
.B(n_15),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_146),
.A2(n_129),
.B1(n_106),
.B2(n_118),
.Y(n_220)
);

BUFx4f_ASAP7_75t_SL g221 ( 
.A(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_129),
.A2(n_37),
.B1(n_25),
.B2(n_43),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_190),
.A2(n_127),
.B1(n_152),
.B2(n_151),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_229),
.A2(n_237),
.B1(n_243),
.B2(n_255),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_233),
.A2(n_203),
.B(n_175),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_181),
.A2(n_149),
.B1(n_152),
.B2(n_161),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_234),
.A2(n_262),
.B(n_195),
.C(n_199),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_241),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_205),
.A2(n_159),
.B1(n_121),
.B2(n_149),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_168),
.A2(n_109),
.B1(n_108),
.B2(n_79),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_250),
.A2(n_260),
.B1(n_270),
.B2(n_198),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_159),
.B1(n_121),
.B2(n_108),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_193),
.A2(n_217),
.B1(n_182),
.B2(n_204),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_257),
.A2(n_166),
.B1(n_201),
.B2(n_178),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_170),
.A2(n_79),
.B1(n_67),
.B2(n_58),
.Y(n_260)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_67),
.B1(n_45),
.B2(n_43),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_45),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_185),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_167),
.B(n_188),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_274),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_197),
.A2(n_45),
.B1(n_43),
.B2(n_15),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_172),
.B(n_14),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_211),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_276),
.B(n_282),
.Y(n_345)
);

OA22x2_ASAP7_75t_L g321 ( 
.A1(n_277),
.A2(n_234),
.B1(n_249),
.B2(n_262),
.Y(n_321)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_231),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_281),
.B(n_297),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_189),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_183),
.B1(n_184),
.B2(n_180),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_291),
.A2(n_292),
.B1(n_319),
.B2(n_228),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_164),
.B1(n_186),
.B2(n_165),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_200),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_294),
.B(n_295),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_186),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_308),
.B(n_292),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_244),
.A2(n_185),
.B(n_221),
.C(n_166),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_300),
.Y(n_325)
);

INVx6_ASAP7_75t_SL g300 ( 
.A(n_232),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_316),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_238),
.B(n_218),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_303),
.Y(n_323)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_310),
.Y(n_331)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_233),
.B(n_187),
.C(n_196),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_309),
.C(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_317),
.Y(n_341)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_314),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_313),
.A2(n_230),
.B(n_266),
.Y(n_335)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_228),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_273),
.A2(n_221),
.B1(n_13),
.B2(n_2),
.Y(n_316)
);

AND2x6_ASAP7_75t_L g317 ( 
.A(n_234),
.B(n_13),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_235),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_226),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_234),
.A2(n_237),
.B1(n_262),
.B2(n_242),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_SL g378 ( 
.A1(n_321),
.A2(n_334),
.B(n_304),
.C(n_307),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_262),
.B1(n_249),
.B2(n_253),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_322),
.A2(n_277),
.B1(n_315),
.B2(n_300),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_326),
.B(n_318),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_239),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_330),
.B(n_354),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_332),
.A2(n_350),
.B1(n_319),
.B2(n_348),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_333),
.A2(n_335),
.B1(n_339),
.B2(n_344),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_285),
.A2(n_266),
.B1(n_230),
.B2(n_225),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_224),
.C(n_246),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_348),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_285),
.A2(n_225),
.B1(n_246),
.B2(n_224),
.Y(n_344)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_248),
.C(n_247),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_320),
.A2(n_248),
.B1(n_235),
.B2(n_254),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_311),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_353),
.B(n_358),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_236),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_0),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_361),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_277),
.A2(n_0),
.B(n_4),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_356),
.A2(n_347),
.B(n_361),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_293),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_290),
.Y(n_362)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_373),
.Y(n_397)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_370),
.A2(n_381),
.B1(n_367),
.B2(n_388),
.Y(n_427)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_388),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_332),
.A2(n_334),
.B1(n_350),
.B2(n_326),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_377),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_341),
.A2(n_277),
.B1(n_317),
.B2(n_280),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_384),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_323),
.B(n_283),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_376),
.B(n_383),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_325),
.Y(n_377)
);

OAI21xp33_ASAP7_75t_SL g421 ( 
.A1(n_378),
.A2(n_391),
.B(n_336),
.Y(n_421)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_379),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_333),
.A2(n_310),
.B1(n_306),
.B2(n_312),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_345),
.B(n_288),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_341),
.A2(n_299),
.B1(n_289),
.B2(n_275),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_321),
.C(n_327),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_324),
.B(n_329),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_386),
.B(n_349),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_286),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_390),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_356),
.A2(n_335),
.B(n_325),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_329),
.B(n_351),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_389),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_284),
.Y(n_390)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_321),
.B(n_314),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_4),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_393),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_343),
.B(n_4),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_395),
.Y(n_419)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_337),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_5),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_340),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_330),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_403),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_417),
.C(n_384),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_321),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_382),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_407),
.B(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_365),
.B(n_339),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_413),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_378),
.A2(n_359),
.B(n_346),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_411),
.A2(n_421),
.B(n_378),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_344),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_373),
.B(n_337),
.C(n_360),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_336),
.Y(n_420)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_368),
.B(n_328),
.Y(n_422)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_328),
.Y(n_423)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_425),
.B(n_424),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_340),
.Y(n_426)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_366),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_428),
.A2(n_415),
.B1(n_422),
.B2(n_423),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_397),
.A2(n_367),
.B1(n_372),
.B2(n_378),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_435),
.B1(n_447),
.B2(n_427),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_434),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_420),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_431),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_448),
.C(n_450),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_363),
.C(n_378),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_376),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_436),
.A2(n_441),
.B1(n_414),
.B2(n_444),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_375),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_440),
.B(n_451),
.Y(n_459)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_443),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_398),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_397),
.A2(n_381),
.B1(n_363),
.B2(n_391),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_402),
.C(n_403),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_407),
.B(n_391),
.C(n_387),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_364),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_394),
.C(n_371),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_418),
.C(n_6),
.Y(n_473)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_457),
.A2(n_446),
.B(n_452),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_429),
.A2(n_398),
.B1(n_404),
.B2(n_406),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_447),
.A2(n_404),
.B1(n_406),
.B2(n_412),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_462),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_435),
.A2(n_412),
.B1(n_399),
.B2(n_410),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_466),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_426),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_468),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_430),
.B(n_415),
.CI(n_410),
.CON(n_469),
.SN(n_469)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_469),
.B(n_472),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_470),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_438),
.B(n_395),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_434),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_428),
.A2(n_418),
.B1(n_374),
.B2(n_7),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_474),
.C(n_453),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_5),
.C(n_7),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_483),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_486),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_432),
.C(n_439),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_482),
.C(n_437),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_439),
.C(n_440),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_437),
.Y(n_483)
);

BUFx4f_ASAP7_75t_SL g484 ( 
.A(n_465),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_463),
.B(n_445),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_451),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_490),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_460),
.B(n_450),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_457),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_454),
.B(n_458),
.Y(n_492)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_492),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_476),
.B(n_474),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_496),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_480),
.A2(n_482),
.B(n_484),
.Y(n_495)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_484),
.A2(n_467),
.B(n_461),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_503),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_500),
.C(n_483),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_464),
.C(n_473),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_456),
.C(n_469),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_504),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_475),
.A2(n_471),
.B(n_466),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_456),
.C(n_469),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_496),
.A2(n_488),
.B1(n_487),
.B2(n_472),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_506),
.B(n_513),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_512),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_487),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_479),
.B(n_485),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_514),
.A2(n_505),
.B(n_477),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_500),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_518),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_498),
.C(n_491),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_521),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_505),
.B(n_498),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_515),
.C(n_509),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_525),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_511),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_524),
.A2(n_510),
.B(n_449),
.Y(n_527)
);

O2A1O1Ixp33_ASAP7_75t_SL g528 ( 
.A1(n_527),
.A2(n_523),
.B(n_526),
.C(n_468),
.Y(n_528)
);

O2A1O1Ixp33_ASAP7_75t_SL g529 ( 
.A1(n_528),
.A2(n_462),
.B(n_438),
.C(n_9),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_5),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_5),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_10),
.Y(n_532)
);

OAI332xp33_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_484),
.B3(n_465),
.C1(n_436),
.C2(n_530),
.Y(n_533)
);


endmodule