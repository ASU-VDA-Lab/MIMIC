module fake_jpeg_30751_n_359 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_359);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_23),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_79),
.B1(n_88),
.B2(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_78),
.B(n_84),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_40),
.B1(n_33),
.B2(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_85),
.B1(n_25),
.B2(n_44),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_53),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

HAxp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_30),
.CON(n_84),
.SN(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_35),
.B1(n_25),
.B2(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_34),
.B1(n_30),
.B2(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_43),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_38),
.C(n_31),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_70),
.C(n_69),
.Y(n_150)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_123),
.B1(n_93),
.B2(n_74),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_29),
.B1(n_31),
.B2(n_42),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_29),
.B1(n_32),
.B2(n_42),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_38),
.B1(n_32),
.B2(n_45),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_91),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_27),
.B1(n_36),
.B2(n_3),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_87),
.A2(n_27),
.B1(n_36),
.B2(n_3),
.Y(n_122)
);

NOR2x1_ASAP7_75t_R g146 ( 
.A(n_122),
.B(n_125),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_76),
.B1(n_95),
.B2(n_74),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_36),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_130),
.Y(n_144)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_129),
.Y(n_136)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_36),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_4),
.Y(n_148)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_150),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_148),
.B1(n_105),
.B2(n_131),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_130),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_153),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_93),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_79),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_157),
.C(n_141),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_73),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_111),
.B1(n_88),
.B2(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_173),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_119),
.B1(n_129),
.B2(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_140),
.B1(n_170),
.B2(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_167),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_168),
.A2(n_174),
.B(n_146),
.C(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_156),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_150),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_104),
.B1(n_103),
.B2(n_102),
.Y(n_173)
);

FAx1_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_105),
.CI(n_104),
.CON(n_174),
.SN(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_102),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_178),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_70),
.B(n_106),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_141),
.B(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_188),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_138),
.C(n_145),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_187),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_148),
.B(n_173),
.C(n_137),
.D(n_166),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_156),
.B1(n_159),
.B2(n_152),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_175),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_108),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_194),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_136),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_170),
.C(n_174),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_174),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_172),
.B1(n_163),
.B2(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_208),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_186),
.A2(n_147),
.B1(n_179),
.B2(n_169),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_199),
.B(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_212),
.C(n_217),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_174),
.A3(n_168),
.B1(n_162),
.B2(n_163),
.C1(n_176),
.C2(n_173),
.Y(n_210)
);

OAI221xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_215),
.B1(n_103),
.B2(n_107),
.C(n_121),
.Y(n_242)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_162),
.C(n_164),
.Y(n_212)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_147),
.B1(n_148),
.B2(n_167),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_160),
.C(n_152),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_191),
.B1(n_198),
.B2(n_196),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_160),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_197),
.C(n_143),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_181),
.B1(n_190),
.B2(n_199),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_227),
.B1(n_214),
.B2(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_209),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_184),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_184),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_184),
.B1(n_198),
.B2(n_181),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_4),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_219),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_143),
.C(n_135),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_237),
.C(n_232),
.Y(n_245)
);

AO21x2_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_205),
.B(n_201),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_234),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_135),
.C(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_242),
.B(n_134),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_256),
.C(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_250),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_247),
.B(n_264),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_200),
.B1(n_218),
.B2(n_209),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_255),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_216),
.C(n_220),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_234),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_239),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_112),
.B1(n_128),
.B2(n_126),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_134),
.C(n_124),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_223),
.B1(n_221),
.B2(n_225),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_5),
.C(n_6),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_235),
.C(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_270),
.B(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_236),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_278),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_251),
.A2(n_234),
.B(n_227),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_234),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_234),
.B1(n_7),
.B2(n_8),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_5),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_246),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_20),
.B1(n_10),
.B2(n_11),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_245),
.C(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_296),
.C(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_262),
.C(n_257),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_250),
.C(n_244),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_272),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_277),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_244),
.C(n_247),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_252),
.C(n_261),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_286),
.C(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_302),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_266),
.A2(n_7),
.B(n_10),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_297),
.B(n_292),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_267),
.B1(n_285),
.B2(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_309),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_313),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_290),
.A2(n_280),
.B1(n_270),
.B2(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_301),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_13),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_284),
.C(n_10),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_317),
.C(n_289),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_294),
.B(n_7),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_13),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_318),
.B(n_326),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_324),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_296),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_322),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_298),
.Y(n_323)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_15),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_13),
.C(n_14),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_15),
.B(n_16),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_315),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_338),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_328),
.A2(n_327),
.B1(n_313),
.B2(n_318),
.Y(n_332)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_321),
.A2(n_310),
.B(n_311),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_334),
.A2(n_17),
.B(n_18),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_16),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_340),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_16),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_342),
.A2(n_346),
.B(n_337),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_334),
.A2(n_17),
.B(n_18),
.Y(n_343)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_343),
.Y(n_351)
);

AOI21x1_ASAP7_75t_SL g344 ( 
.A1(n_333),
.A2(n_17),
.B(n_18),
.Y(n_344)
);

AO21x2_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_19),
.B(n_20),
.Y(n_353)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_347),
.A2(n_336),
.B(n_335),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_350),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_348),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_353),
.B(n_341),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_354),
.B(n_351),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_356),
.A2(n_355),
.B(n_345),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_353),
.B(n_19),
.Y(n_358)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_358),
.Y(n_359)
);


endmodule