module real_jpeg_31474_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g424 ( 
.A(n_0),
.Y(n_424)
);

NAND2xp67_ASAP7_75t_SL g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_1),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_1),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_1),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_1),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_1),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_2),
.B(n_559),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_2),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_3),
.Y(n_226)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_5),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_6),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_6),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_6),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_6),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_6),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_7),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_7),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_7),
.B(n_116),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_7),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_8),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_8),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_8),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_8),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_8),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_8),
.B(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_9),
.B(n_286),
.Y(n_285)
);

NAND2x1_ASAP7_75t_L g300 ( 
.A(n_9),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_9),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_9),
.B(n_432),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_9),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_10),
.B(n_72),
.Y(n_71)
);

NAND2x2_ASAP7_75t_L g104 ( 
.A(n_10),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_10),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_10),
.B(n_127),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_56),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_13),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_13),
.B(n_292),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_13),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_13),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_13),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_14),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_15),
.Y(n_559)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_16),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_16),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_16),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_17),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_17),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_17),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_17),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_17),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_17),
.B(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_17),
.B(n_455),
.Y(n_454)
);

OAI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_520),
.B1(n_560),
.B2(n_564),
.C(n_565),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_19),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_243),
.B(n_516),
.Y(n_19)
);

NAND2x1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_194),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_22),
.A2(n_518),
.B(n_519),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_157),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_23),
.B(n_157),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_93),
.C(n_129),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_24),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_62),
.C(n_76),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_26),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_40),
.C(n_49),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_27),
.B(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_27)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_29),
.A2(n_30),
.B1(n_234),
.B2(n_363),
.Y(n_553)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_37),
.C(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_33),
.A2(n_128),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_33),
.A2(n_75),
.B1(n_227),
.B2(n_348),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AO22x1_ASAP7_75t_SL g467 ( 
.A1(n_36),
.A2(n_37),
.B1(n_468),
.B2(n_471),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_46),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_37),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_37),
.B(n_471),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_40),
.B(n_49),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_48),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_44),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_46),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_46),
.A2(n_217),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_46),
.B(n_260),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_47),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_47),
.Y(n_447)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_47),
.Y(n_470)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_48),
.B(n_280),
.C(n_285),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_48),
.B(n_502),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_51),
.A2(n_299),
.B1(n_300),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_51),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_51),
.B(n_104),
.C(n_299),
.Y(n_335)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_53),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_55),
.B(n_58),
.C(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_63),
.A2(n_64),
.B1(n_77),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_66),
.B(n_71),
.C(n_74),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_66),
.A2(n_73),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_66),
.A2(n_73),
.B1(n_90),
.B2(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_66),
.B(n_166),
.C(n_167),
.Y(n_528)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_72),
.Y(n_539)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_78),
.C(n_89),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_78),
.B(n_236),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_86),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_79),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_79),
.B(n_152),
.C(n_153),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_79),
.A2(n_86),
.B1(n_151),
.B2(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_83),
.B(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_85),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_85),
.Y(n_433)
);

CKINVDCx12_ASAP7_75t_R g208 ( 
.A(n_86),
.Y(n_208)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_90),
.Y(n_237)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_92),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_94),
.A2(n_131),
.B1(n_193),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_94),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_111),
.C(n_122),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

AOI21x1_ASAP7_75t_SL g186 ( 
.A1(n_97),
.A2(n_187),
.B(n_190),
.Y(n_186)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_101),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_101),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_103),
.B(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_104),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_104),
.B(n_106),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_104),
.B(n_174),
.C(n_182),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_123),
.C(n_128),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_123),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_106),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_106),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_106),
.B(n_251),
.C(n_253),
.Y(n_324)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_108),
.Y(n_233)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_108),
.Y(n_334)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_108),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_122),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_119),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_112),
.A2(n_136),
.B1(n_234),
.B2(n_363),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_112),
.B(n_179),
.C(n_234),
.Y(n_550)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_119),
.B1(n_120),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_115),
.B(n_174),
.C(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_SL g337 ( 
.A(n_115),
.Y(n_337)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_117),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_142),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.C(n_139),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_142),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_144),
.C(n_192),
.Y(n_191)
);

XOR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_153),
.A2(n_154),
.B1(n_552),
.B2(n_553),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_191),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_159),
.B(n_160),
.C(n_191),
.Y(n_524)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_170),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_161),
.B(n_185),
.C(n_543),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_180),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_171),
.A2(n_181),
.B1(n_182),
.B2(n_544),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_171),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_178),
.B2(n_179),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_174),
.A2(n_179),
.B1(n_210),
.B2(n_339),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_174),
.A2(n_179),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_176),
.Y(n_309)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_176),
.Y(n_458)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_SL g260 ( 
.A(n_189),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_239),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_195),
.B(n_239),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_204),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_196),
.B(n_200),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_204),
.B(n_395),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_218),
.B(n_238),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_205),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_214),
.Y(n_205)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_209),
.A2(n_214),
.B1(n_215),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_209),
.Y(n_370)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_210),
.Y(n_339)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_235),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_235),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_219),
.B(n_235),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_231),
.C(n_234),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_220),
.A2(n_221),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.C(n_227),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_222),
.B(n_224),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_227),
.Y(n_348)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_233),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_234),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_397),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_375),
.B(n_389),
.C(n_396),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_350),
.B(n_374),
.Y(n_245)
);

NAND2x1p5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_325),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g399 ( 
.A(n_247),
.B(n_325),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_277),
.C(n_303),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_249),
.B(n_507),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.C(n_263),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_250),
.B(n_496),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_257),
.A2(n_258),
.B1(n_263),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_262),
.Y(n_414)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_263),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.C(n_272),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_273),
.Y(n_486)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_268),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_278),
.B(n_304),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_289),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_279),
.B(n_290),
.C(n_297),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_280),
.B(n_285),
.Y(n_502)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_297),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_294),
.B(n_296),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_294),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_366),
.C(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_320),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_321),
.C(n_323),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_313),
.C(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_313),
.B1(n_318),
.B2(n_319),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_341),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_342),
.C(n_343),
.Y(n_373)
);

XOR2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_340),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_336),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_340),
.C(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_335),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_331),
.C(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_373),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_373),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_377),
.C(n_378),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_368),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_355),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_360),
.B2(n_364),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_360),
.Y(n_364)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_374),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_379),
.B1(n_390),
.B2(n_394),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_376),
.B(n_379),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.C(n_383),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_387),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_394),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_390),
.B(n_394),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.C(n_393),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_511),
.C(n_512),
.Y(n_397)
);

NOR2x1p5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

AOI21x1_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_505),
.B(n_510),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_493),
.B(n_504),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_473),
.B(n_491),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_449),
.B(n_472),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_426),
.B(n_448),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_406),
.A2(n_421),
.B(n_425),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_412),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_412),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_415),
.B1(n_416),
.B2(n_420),
.Y(n_412)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_413),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_415),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_420),
.Y(n_427)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_443),
.Y(n_442)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_428),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_440),
.B2(n_441),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_434),
.C(n_440),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_444),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_451),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_463),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_464),
.C(n_467),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_459),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_457),
.C(n_459),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_468),
.Y(n_471)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

NAND3xp33_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_487),
.C(n_490),
.Y(n_473)
);

O2A1O1Ixp5_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_475),
.B(n_490),
.C(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_481),
.Y(n_474)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_475),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_480),
.C(n_500),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_478),
.Y(n_500)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_484),
.C(n_488),
.Y(n_503)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_489),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_503),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_503),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_498),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_499),
.C(n_509),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_508),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_515),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVxp67_ASAP7_75t_R g516 ( 
.A(n_517),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_545),
.C(n_557),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

AOI221xp5_ASAP7_75t_SL g565 ( 
.A1(n_522),
.A2(n_557),
.B1(n_561),
.B2(n_566),
.C(n_567),
.Y(n_565)
);

NOR4xp25_ASAP7_75t_L g567 ( 
.A(n_522),
.B(n_546),
.C(n_558),
.D(n_562),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_524),
.B(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_525),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_542),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_528),
.B(n_529),
.C(n_542),
.Y(n_555)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_534),
.B1(n_535),
.B2(n_541),
.Y(n_530)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_531),
.Y(n_541)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_537),
.B1(n_538),
.B2(n_540),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_540),
.C(n_541),
.Y(n_554)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_538),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_558),
.Y(n_561)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_556),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_555),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_555),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_554),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_551),
.Y(n_549)
);

CKINVDCx11_ASAP7_75t_R g552 ( 
.A(n_553),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_558),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_562),
.Y(n_560)
);


endmodule