module fake_jpeg_17908_n_113 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_55),
.B1(n_42),
.B2(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_50),
.B1(n_53),
.B2(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_52),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_87),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_26),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_68),
.C(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_89),
.B(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_99),
.B1(n_10),
.B2(n_12),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_101),
.B1(n_13),
.B2(n_15),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_8),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_20),
.C(n_22),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_30),
.B(n_31),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_33),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_34),
.B(n_37),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_38),
.Y(n_113)
);


endmodule