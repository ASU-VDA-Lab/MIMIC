module fake_jpeg_29751_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_0),
.B(n_2),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_25),
.C(n_24),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_24),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_27),
.B1(n_25),
.B2(n_14),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_53),
.B1(n_60),
.B2(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_14),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_17),
.B1(n_19),
.B2(n_28),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_38),
.B1(n_26),
.B2(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_84),
.B1(n_90),
.B2(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_73),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_30),
.B1(n_23),
.B2(n_21),
.Y(n_74)
);

AO22x2_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_87),
.B1(n_88),
.B2(n_91),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_21),
.Y(n_75)
);

XNOR2x1_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_78),
.Y(n_97)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_10),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_55),
.B(n_9),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_45),
.B(n_5),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_90),
.B1(n_45),
.B2(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_4),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

AOI22x1_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_55),
.B1(n_45),
.B2(n_63),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_94),
.Y(n_120)
);

NOR2xp67_ASAP7_75t_R g112 ( 
.A(n_96),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_88),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_6),
.B1(n_8),
.B2(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_8),
.B1(n_83),
.B2(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_75),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_113),
.B1(n_121),
.B2(n_110),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_68),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_122),
.C(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_85),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_76),
.B(n_77),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_95),
.B(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_87),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_108),
.C(n_98),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_107),
.C(n_99),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_93),
.C(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_111),
.B(n_96),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_120),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_134),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_120),
.B1(n_123),
.B2(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_99),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.C(n_124),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_114),
.C(n_120),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_135),
.C(n_127),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_150),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_92),
.A3(n_95),
.B1(n_105),
.B2(n_139),
.C1(n_134),
.C2(n_132),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_129),
.B(n_130),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_158),
.B(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_148),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_133),
.B1(n_105),
.B2(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_142),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_158),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_151),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_161),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_167),
.C(n_166),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_171),
.B(n_166),
.C(n_172),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_162),
.Y(n_175)
);


endmodule