module fake_jpeg_10997_n_201 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g72 ( 
.A(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.Y(n_103)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_58),
.B1(n_70),
.B2(n_86),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_102),
.B1(n_106),
.B2(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_107),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_62),
.B1(n_79),
.B2(n_61),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_95),
.B1(n_89),
.B2(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_73),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_92),
.B1(n_91),
.B2(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_130),
.B1(n_118),
.B2(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_132),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_92),
.B1(n_64),
.B2(n_80),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_7),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_68),
.B1(n_71),
.B2(n_76),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_126),
.B1(n_4),
.B2(n_6),
.Y(n_145)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_66),
.B(n_72),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_124),
.C(n_0),
.Y(n_140)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_66),
.B(n_83),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_69),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_129),
.C(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_78),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_69),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_73),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_59),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_6),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_71),
.B1(n_68),
.B2(n_76),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_139),
.B1(n_145),
.B2(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_152),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_R g168 ( 
.A(n_140),
.B(n_16),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_17),
.B(n_18),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_156),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_12),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_29),
.B1(n_55),
.B2(n_51),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_14),
.B2(n_15),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_9),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_161),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_10),
.B(n_11),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_141),
.B(n_153),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_171),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_173),
.C(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_139),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_143),
.B(n_153),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_147),
.B(n_155),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_163),
.A3(n_168),
.B1(n_164),
.B2(n_159),
.C1(n_17),
.C2(n_32),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_159),
.B1(n_166),
.B2(n_162),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_174),
.C(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_161),
.B1(n_21),
.B2(n_22),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_179),
.Y(n_192)
);

AOI321xp33_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_192),
.A3(n_184),
.B1(n_183),
.B2(n_188),
.C(n_186),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_184),
.B(n_188),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_191),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_20),
.B(n_31),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_39),
.C(n_40),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_41),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_44),
.B(n_46),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_50),
.Y(n_201)
);


endmodule