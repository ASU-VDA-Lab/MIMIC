module fake_jpeg_12188_n_594 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_594);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_594;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_16),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_61),
.B(n_77),
.Y(n_117)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_68),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_17),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_100),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_37),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_90),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_15),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_48),
.B(n_14),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_108),
.Y(n_156)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_52),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_36),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_52),
.B1(n_50),
.B2(n_43),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_44),
.B1(n_46),
.B2(n_42),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_43),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_145),
.B(n_150),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_41),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_41),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_45),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_80),
.B(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_82),
.B(n_51),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_82),
.B(n_51),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_175),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_62),
.B(n_32),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_44),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx12_ASAP7_75t_R g173 ( 
.A(n_103),
.Y(n_173)
);

CKINVDCx12_ASAP7_75t_R g216 ( 
.A(n_173),
.Y(n_216)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_42),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_55),
.Y(n_176)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_177),
.B(n_185),
.Y(n_245)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_179),
.Y(n_282)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_180),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_182),
.A2(n_192),
.B1(n_206),
.B2(n_218),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_36),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_186),
.Y(n_258)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_117),
.B(n_40),
.C(n_26),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_225),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_126),
.A2(n_105),
.B1(n_96),
.B2(n_93),
.Y(n_192)
);

OR2x4_ASAP7_75t_L g193 ( 
.A(n_114),
.B(n_37),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_193),
.B(n_209),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_136),
.A2(n_92),
.B1(n_87),
.B2(n_60),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_199),
.A2(n_204),
.B1(n_237),
.B2(n_239),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_46),
.B(n_1),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_136),
.A2(n_44),
.B1(n_32),
.B2(n_47),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_111),
.A2(n_89),
.B1(n_109),
.B2(n_84),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_125),
.B(n_36),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_40),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_215),
.B(n_217),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_46),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_112),
.A2(n_71),
.B1(n_70),
.B2(n_69),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_120),
.B(n_13),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_219),
.B(n_229),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_118),
.A2(n_67),
.B1(n_59),
.B2(n_56),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_224),
.A2(n_139),
.B1(n_50),
.B2(n_54),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_122),
.Y(n_225)
);

CKINVDCx6p67_ASAP7_75t_R g226 ( 
.A(n_146),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_227),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_128),
.B(n_13),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_233),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_169),
.A2(n_37),
.B(n_44),
.C(n_47),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_231),
.Y(n_274)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_120),
.B(n_54),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_127),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_141),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_236),
.Y(n_241)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_155),
.Y(n_237)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_32),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_240),
.A2(n_54),
.B(n_47),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_144),
.B1(n_113),
.B2(n_116),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_243),
.A2(n_248),
.B1(n_249),
.B2(n_267),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_259),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_170),
.B1(n_123),
.B2(n_113),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_204),
.A2(n_170),
.B1(n_123),
.B2(n_116),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g252 ( 
.A1(n_191),
.A2(n_146),
.A3(n_169),
.B1(n_168),
.B2(n_155),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_252),
.B(n_0),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_148),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_186),
.B(n_162),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_265),
.B(n_285),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_199),
.A2(n_144),
.B1(n_160),
.B2(n_166),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_231),
.B(n_137),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_284),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_190),
.A2(n_160),
.B1(n_171),
.B2(n_134),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_273),
.A2(n_296),
.B1(n_194),
.B2(n_223),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_178),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_200),
.B(n_171),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_205),
.B(n_139),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_297),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_202),
.B1(n_183),
.B2(n_203),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_239),
.A2(n_39),
.B1(n_38),
.B2(n_2),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_189),
.B(n_39),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_299),
.A2(n_346),
.B1(n_248),
.B2(n_281),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_264),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_302),
.B(n_310),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_235),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_303),
.B(n_313),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_213),
.B1(n_227),
.B2(n_198),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_309),
.A2(n_335),
.B1(n_326),
.B2(n_293),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx13_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_246),
.B(n_256),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_253),
.B(n_230),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_314),
.B(n_316),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_241),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_322),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_259),
.B(n_214),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_318),
.Y(n_366)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_201),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_324),
.B(n_329),
.Y(n_370)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_327),
.B(n_328),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_261),
.B(n_269),
.Y(n_328)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_226),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_226),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_331),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_265),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_184),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_334),
.Y(n_390)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_336),
.Y(n_393)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_262),
.B(n_187),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_338),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_266),
.B(n_220),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_340),
.Y(n_358)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

INVx13_ASAP7_75t_L g341 ( 
.A(n_260),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_274),
.B(n_195),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_0),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_344),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_234),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_271),
.B(n_234),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_345),
.B(n_286),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_254),
.A2(n_39),
.B1(n_38),
.B2(n_3),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_347),
.A2(n_291),
.B(n_242),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_271),
.B(n_1),
.C(n_3),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_297),
.C(n_288),
.Y(n_354)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_276),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_349),
.A2(n_336),
.B1(n_282),
.B2(n_289),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_350),
.A2(n_359),
.B1(n_384),
.B2(n_391),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_354),
.B(n_337),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_332),
.A2(n_266),
.B(n_251),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_356),
.A2(n_368),
.B(n_371),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_347),
.A2(n_254),
.B1(n_297),
.B2(n_289),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_292),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_362),
.B(n_363),
.C(n_375),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_286),
.C(n_295),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_367),
.B1(n_336),
.B2(n_340),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_326),
.A2(n_260),
.B1(n_290),
.B2(n_282),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_339),
.A2(n_270),
.B(n_280),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_275),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_295),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_385),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_335),
.A2(n_306),
.B1(n_343),
.B2(n_311),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_332),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_348),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_301),
.B(n_275),
.C(n_291),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_287),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_320),
.C(n_341),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_332),
.A2(n_242),
.B1(n_257),
.B2(n_287),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_301),
.A2(n_280),
.B(n_270),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_392),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_353),
.B(n_315),
.Y(n_395)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_395),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_356),
.A2(n_308),
.B(n_324),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_421),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_399),
.B(n_391),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_365),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_400),
.B(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_401),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_402),
.B(n_354),
.C(n_361),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_327),
.Y(n_403)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_351),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_407),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_412),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_381),
.B(n_298),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_410),
.B(n_411),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_322),
.Y(n_411)
);

OAI32xp33_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_329),
.A3(n_349),
.B1(n_325),
.B2(n_336),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_317),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_413),
.B(n_416),
.Y(n_463)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_318),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_419),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_319),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_373),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_372),
.B(n_305),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_431),
.C(n_433),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_312),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_334),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_422),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_392),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_363),
.B(n_321),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_424),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_369),
.B(n_307),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_304),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_427),
.Y(n_455)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_4),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_257),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_385),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_393),
.B(n_4),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_429),
.A2(n_368),
.B(n_358),
.Y(n_436)
);

AO22x1_ASAP7_75t_L g479 ( 
.A1(n_436),
.A2(n_418),
.B1(n_405),
.B2(n_421),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_395),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_438),
.B(n_439),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_403),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_430),
.A2(n_383),
.B1(n_372),
.B2(n_374),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_443),
.A2(n_454),
.B1(n_456),
.B2(n_466),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_396),
.A2(n_399),
.B1(n_404),
.B2(n_401),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_419),
.B1(n_415),
.B2(n_427),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_460),
.C(n_450),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_457),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_358),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_453),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_409),
.A2(n_374),
.B1(n_350),
.B2(n_361),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_425),
.A2(n_378),
.B1(n_366),
.B2(n_360),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_406),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_398),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_371),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_420),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_465),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_412),
.A2(n_360),
.B1(n_382),
.B2(n_379),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_468),
.A2(n_453),
.B1(n_405),
.B2(n_422),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_414),
.Y(n_469)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_470),
.A2(n_490),
.B1(n_479),
.B2(n_437),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_435),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_472),
.B(n_492),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_447),
.B(n_397),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_475),
.Y(n_503)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_442),
.Y(n_476)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_476),
.Y(n_518)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_477),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_408),
.C(n_432),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_480),
.C(n_484),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_R g519 ( 
.A(n_479),
.B(n_7),
.C(n_8),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_397),
.C(n_426),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_481),
.A2(n_493),
.B1(n_496),
.B2(n_466),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_428),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_489),
.Y(n_509)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_483),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_379),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_485),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_382),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_394),
.C(n_352),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_456),
.C(n_436),
.Y(n_505)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_455),
.A2(n_352),
.B1(n_394),
.B2(n_355),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_459),
.A2(n_355),
.B(n_6),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_495),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_5),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_462),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_497),
.B(n_440),
.Y(n_511)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_486),
.B(n_446),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_500),
.B(n_517),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_487),
.A2(n_444),
.B1(n_468),
.B2(n_437),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_504),
.A2(n_496),
.B1(n_477),
.B2(n_476),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_515),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_463),
.Y(n_506)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_445),
.C(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_508),
.B(n_511),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_510),
.A2(n_487),
.B1(n_473),
.B2(n_479),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_445),
.C(n_453),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_521),
.C(n_471),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_488),
.A2(n_455),
.B1(n_452),
.B2(n_441),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_497),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_480),
.B(n_468),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_467),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_8),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_491),
.B(n_462),
.Y(n_517)
);

AO21x1_ASAP7_75t_L g541 ( 
.A1(n_519),
.A2(n_11),
.B(n_12),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_474),
.B(n_482),
.C(n_470),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_523),
.B(n_529),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_524),
.A2(n_520),
.B1(n_501),
.B2(n_518),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_513),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_534),
.Y(n_543)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_507),
.Y(n_528)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_469),
.B(n_485),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_530),
.A2(n_523),
.B(n_527),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_521),
.B(n_489),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_531),
.B(n_536),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_495),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_505),
.A2(n_7),
.B(n_8),
.Y(n_535)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_535),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_9),
.C(n_10),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_539),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_9),
.C(n_10),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_9),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_537),
.Y(n_546)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_541),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_538),
.Y(n_544)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_544),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_499),
.C(n_503),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_546),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_522),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_548),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_549),
.B(n_551),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_530),
.A2(n_519),
.B(n_520),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_509),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_555),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_509),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_547),
.A2(n_529),
.B1(n_541),
.B2(n_533),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_567),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_550),
.Y(n_561)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_561),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_545),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_565),
.A2(n_558),
.B(n_559),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_543),
.A2(n_539),
.B(n_531),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_549),
.A2(n_532),
.B(n_503),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_569),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_554),
.B(n_512),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_536),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_571),
.B(n_546),
.C(n_540),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_572),
.B(n_573),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_566),
.B(n_559),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_574),
.A2(n_570),
.B(n_563),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_564),
.B(n_551),
.C(n_557),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_577),
.B(n_579),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_556),
.C(n_552),
.Y(n_579)
);

OA21x2_ASAP7_75t_SL g581 ( 
.A1(n_576),
.A2(n_575),
.B(n_578),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_581),
.B(n_512),
.C(n_11),
.Y(n_587)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_582),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_574),
.A2(n_570),
.B1(n_563),
.B2(n_561),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_583),
.B(n_571),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_585),
.A2(n_587),
.B(n_584),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_588),
.B(n_589),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_586),
.B(n_583),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_580),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_591),
.B(n_11),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_12),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_593),
.B(n_12),
.Y(n_594)
);


endmodule