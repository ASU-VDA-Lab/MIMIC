module fake_jpeg_27231_n_159 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_159);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_23),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_28),
.Y(n_70)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_48),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_34),
.B1(n_21),
.B2(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_59),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_32),
.B(n_17),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_19),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_29),
.B(n_23),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_65),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_23),
.B(n_35),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_61),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_16),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_69),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_42),
.B1(n_39),
.B2(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_80),
.Y(n_103)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_42),
.B1(n_17),
.B2(n_27),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_58),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_96),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_52),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_101),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_51),
.C(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_100),
.C(n_105),
.Y(n_121)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_66),
.C(n_49),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_53),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_20),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_26),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_25),
.C(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_87),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_87),
.B1(n_71),
.B2(n_76),
.C(n_90),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_111),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_84),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_79),
.B(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_25),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_18),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_102),
.B1(n_100),
.B2(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_94),
.C(n_105),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_134),
.C(n_122),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_18),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_131),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_24),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_26),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

OA21x2_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_115),
.B(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_120),
.B(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_127),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_146),
.A2(n_140),
.B1(n_125),
.B2(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_141),
.C(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_26),
.C(n_7),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_5),
.B1(n_11),
.B2(n_9),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_152),
.A3(n_144),
.B1(n_143),
.B2(n_13),
.C1(n_8),
.C2(n_4),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_149),
.B1(n_3),
.B2(n_4),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_157),
.C(n_153),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);


endmodule