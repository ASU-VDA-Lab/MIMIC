module fake_jpeg_8189_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_12),
.B1(n_18),
.B2(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_33),
.B1(n_12),
.B2(n_29),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_40),
.B1(n_25),
.B2(n_14),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_23),
.B1(n_22),
.B2(n_14),
.Y(n_53)
);

OA22x2_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_16),
.Y(n_45)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_39),
.B1(n_34),
.B2(n_43),
.Y(n_75)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_12),
.A3(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_20),
.B1(n_17),
.B2(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_25),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_45),
.B(n_52),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

XOR2x1_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_16),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_46),
.B(n_39),
.C(n_38),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_67),
.B1(n_72),
.B2(n_75),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_53),
.B(n_54),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_44),
.B1(n_36),
.B2(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_17),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_83),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_94),
.B1(n_75),
.B2(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_49),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_75),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_65),
.C(n_72),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_104),
.C(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_62),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_106),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_113),
.C(n_117),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_86),
.C(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_93),
.A3(n_89),
.B1(n_80),
.B2(n_90),
.C(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_109),
.B1(n_104),
.B2(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_101),
.B1(n_93),
.B2(n_100),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_125),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_101),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_124),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_92),
.B1(n_76),
.B2(n_38),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_3),
.B(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_8),
.C(n_11),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_10),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_7),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_131),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.C(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_120),
.B1(n_125),
.B2(n_118),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_118),
.C(n_128),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_138),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_131),
.B(n_130),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_39),
.CI(n_4),
.CON(n_139),
.SN(n_139)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_3),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_140),
.B1(n_138),
.B2(n_141),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_5),
.CI(n_39),
.CON(n_145),
.SN(n_145)
);


endmodule