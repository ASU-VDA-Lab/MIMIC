module fake_aes_11364_n_615 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_615);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_615;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_51), .Y(n_72) );
BUFx3_ASAP7_75t_L g73 ( .A(n_43), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_19), .Y(n_74) );
NOR2xp67_ASAP7_75t_L g75 ( .A(n_57), .B(n_29), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_8), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_41), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_39), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_48), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_56), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_15), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_2), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_11), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_16), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_64), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_7), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_32), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_54), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_65), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_37), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_68), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_4), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_28), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_25), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_23), .B(n_38), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_7), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_27), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_40), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_35), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_33), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_66), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_17), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_11), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_62), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_1), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_73), .B(n_0), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_73), .B(n_0), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_99), .B(n_2), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
XNOR2x2_ASAP7_75t_L g125 ( .A(n_84), .B(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
INVx5_ASAP7_75t_L g128 ( .A(n_99), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_115), .B(n_3), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_86), .B(n_4), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_89), .B(n_5), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_99), .B(n_5), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_94), .B(n_6), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_96), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_102), .B(n_8), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_95), .A2(n_44), .B(n_63), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_105), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_99), .B(n_9), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_98), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_111), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_104), .B(n_10), .Y(n_152) );
OAI21x1_ASAP7_75t_L g153 ( .A1(n_112), .A2(n_45), .B(n_60), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_121), .B(n_92), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_116), .B(n_92), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_120), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_116), .B(n_72), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_117), .B(n_72), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_118), .B(n_113), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_128), .Y(n_163) );
OR2x2_ASAP7_75t_L g164 ( .A(n_141), .B(n_110), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_118), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
INVx6_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
OR2x6_ASAP7_75t_L g169 ( .A(n_150), .B(n_101), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_119), .A2(n_74), .B1(n_91), .B2(n_110), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_117), .B(n_109), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_123), .B(n_109), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_123), .B(n_100), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_124), .B(n_88), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_119), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_124), .B(n_107), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_126), .B(n_91), .Y(n_179) );
OR2x2_ASAP7_75t_L g180 ( .A(n_132), .B(n_12), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_119), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_129), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_126), .B(n_107), .Y(n_185) );
BUFx10_ASAP7_75t_L g186 ( .A(n_119), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_127), .B(n_107), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_130), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_128), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_127), .B(n_74), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_131), .B(n_107), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_132), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_131), .B(n_107), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_128), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_134), .B(n_101), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_134), .B(n_154), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_138), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_125), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_167), .A2(n_154), .B1(n_151), .B2(n_149), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_201), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_194), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_171), .A2(n_145), .B1(n_146), .B2(n_151), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_201), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_202), .Y(n_209) );
BUFx12f_ASAP7_75t_L g210 ( .A(n_164), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_179), .A2(n_146), .B1(n_145), .B2(n_149), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_186), .B(n_153), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_167), .A2(n_135), .B1(n_138), .B2(n_148), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_194), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_155), .B(n_135), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_155), .A2(n_140), .B1(n_152), .B2(n_133), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_186), .B(n_153), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_164), .B(n_142), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_186), .B(n_148), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_161), .B(n_144), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_202), .Y(n_221) );
OR2x4_ASAP7_75t_L g222 ( .A(n_180), .B(n_125), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_202), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_200), .A2(n_144), .B1(n_147), .B2(n_136), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g225 ( .A(n_190), .B(n_13), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_192), .B(n_122), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_172), .B(n_143), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_180), .B(n_13), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_176), .B(n_143), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_176), .B(n_143), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_192), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_157), .B(n_143), .Y(n_233) );
INVxp67_ASAP7_75t_L g234 ( .A(n_156), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_160), .B(n_75), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_158), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_174), .B(n_139), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_173), .B(n_14), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_162), .B(n_18), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_200), .B(n_20), .Y(n_241) );
NOR2x2_ASAP7_75t_L g242 ( .A(n_169), .B(n_21), .Y(n_242) );
OR2x6_ASAP7_75t_L g243 ( .A(n_169), .B(n_22), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_158), .Y(n_244) );
AND2x4_ASAP7_75t_SL g245 ( .A(n_162), .B(n_24), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_167), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_167), .A2(n_26), .B1(n_31), .B2(n_42), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_162), .B(n_46), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_165), .A2(n_47), .B1(n_49), .B2(n_50), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
AND2x6_ASAP7_75t_SL g251 ( .A(n_169), .B(n_53), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_159), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_159), .B(n_55), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_190), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_170), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_203), .Y(n_256) );
NOR2xp67_ASAP7_75t_L g257 ( .A(n_203), .B(n_69), .Y(n_257) );
OAI21xp33_ASAP7_75t_SL g258 ( .A1(n_204), .A2(n_182), .B(n_177), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_255), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_255), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_205), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_230), .A2(n_185), .B(n_178), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_252), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_218), .A2(n_169), .B1(n_197), .B2(n_188), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_231), .A2(n_188), .B(n_197), .C(n_191), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_227), .Y(n_266) );
INVxp67_ASAP7_75t_SL g267 ( .A(n_234), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_215), .Y(n_268) );
AOI221x1_ASAP7_75t_L g269 ( .A1(n_228), .A2(n_187), .B1(n_193), .B2(n_195), .C(n_191), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_253), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_208), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_232), .B(n_184), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_207), .A2(n_184), .B(n_168), .C(n_163), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_237), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_233), .A2(n_163), .B(n_166), .C(n_168), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_212), .A2(n_217), .B(n_219), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_226), .B(n_196), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_233), .A2(n_166), .B(n_175), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_244), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_240), .B(n_175), .Y(n_281) );
BUFx4f_ASAP7_75t_SL g282 ( .A(n_210), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_213), .A2(n_189), .B1(n_196), .B2(n_199), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
NAND2x2_ASAP7_75t_L g286 ( .A(n_222), .B(n_58), .Y(n_286) );
BUFx8_ASAP7_75t_L g287 ( .A(n_229), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
NAND4xp25_ASAP7_75t_SL g289 ( .A(n_204), .B(n_189), .C(n_59), .D(n_199), .Y(n_289) );
BUFx10_ASAP7_75t_L g290 ( .A(n_245), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_211), .B(n_181), .Y(n_292) );
BUFx8_ASAP7_75t_L g293 ( .A(n_240), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_220), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
BUFx12f_ASAP7_75t_L g297 ( .A(n_251), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_214), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_243), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_221), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_272), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_276), .A2(n_217), .B(n_212), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_295), .B(n_216), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_299), .A2(n_256), .B1(n_243), .B2(n_246), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_270), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_275), .A2(n_241), .B(n_248), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_278), .A2(n_247), .B(n_249), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_267), .B(n_213), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_267), .B(n_224), .Y(n_310) );
OAI21x1_ASAP7_75t_SL g311 ( .A1(n_266), .A2(n_247), .B(n_243), .Y(n_311) );
NOR2xp33_ASAP7_75t_SL g312 ( .A(n_293), .B(n_257), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_293), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_264), .B(n_222), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_259), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_268), .B(n_235), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_261), .B(n_236), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_262), .A2(n_238), .B(n_225), .Y(n_318) );
CKINVDCx6p67_ASAP7_75t_R g319 ( .A(n_290), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_269), .A2(n_219), .B(n_239), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_270), .Y(n_323) );
INVx5_ASAP7_75t_L g324 ( .A(n_260), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_260), .B(n_254), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_270), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_287), .A2(n_236), .B1(n_239), .B2(n_242), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_274), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_328), .A2(n_286), .B1(n_298), .B2(n_288), .C(n_271), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_327), .A2(n_297), .B1(n_286), .B2(n_287), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_302), .A2(n_297), .B1(n_283), .B2(n_277), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_302), .A2(n_277), .B1(n_270), .B2(n_296), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_296), .B1(n_281), .B2(n_285), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_324), .Y(n_335) );
BUFx12f_ASAP7_75t_L g336 ( .A(n_327), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_321), .B(n_280), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_322), .Y(n_338) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_312), .B(n_275), .C(n_265), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_322), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_314), .A2(n_277), .B1(n_296), .B2(n_281), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g344 ( .A1(n_304), .A2(n_258), .B(n_265), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_314), .A2(n_296), .B1(n_289), .B2(n_280), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_309), .A2(n_285), .B1(n_259), .B2(n_273), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_324), .B(n_301), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_305), .A2(n_282), .B1(n_263), .B2(n_279), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_313), .A2(n_282), .B1(n_263), .B2(n_279), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_317), .A2(n_300), .B1(n_292), .B2(n_284), .C(n_291), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_310), .A2(n_291), .B1(n_294), .B2(n_290), .C(n_198), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_313), .A2(n_294), .B1(n_183), .B2(n_198), .Y(n_354) );
AND2x4_ASAP7_75t_SL g355 ( .A(n_335), .B(n_343), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_349), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_335), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_349), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_335), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_338), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_337), .B(n_321), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_335), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_337), .B(n_329), .Y(n_365) );
INVx5_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_340), .B(n_329), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_344), .Y(n_368) );
CKINVDCx16_ASAP7_75t_R g369 ( .A(n_336), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_353), .B(n_329), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_347), .B(n_310), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_347), .B(n_315), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_343), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
AO31x2_ASAP7_75t_L g376 ( .A1(n_334), .A2(n_311), .A3(n_308), .B(n_318), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_343), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_303), .Y(n_378) );
INVx3_ASAP7_75t_SL g379 ( .A(n_343), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_330), .B(n_315), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_345), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_378), .B(n_318), .Y(n_386) );
NAND3xp33_ASAP7_75t_SL g387 ( .A(n_383), .B(n_331), .C(n_312), .Y(n_387) );
OAI221xp5_ASAP7_75t_SL g388 ( .A1(n_383), .A2(n_332), .B1(n_348), .B2(n_368), .C(n_384), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_363), .B(n_341), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_365), .B(n_363), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_365), .B(n_303), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_362), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_366), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_379), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_367), .B(n_320), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_382), .B(n_333), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_382), .B(n_350), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_366), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_366), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_367), .B(n_320), .Y(n_405) );
OAI33xp33_ASAP7_75t_L g406 ( .A1(n_381), .A2(n_311), .A3(n_319), .B1(n_352), .B2(n_307), .B3(n_308), .Y(n_406) );
OAI31xp33_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_325), .A3(n_315), .B(n_306), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_382), .B(n_326), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_381), .A2(n_307), .B(n_354), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_356), .Y(n_411) );
OR2x6_ASAP7_75t_L g412 ( .A(n_378), .B(n_325), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_371), .B(n_326), .Y(n_413) );
AOI21xp5_ASAP7_75t_SL g414 ( .A1(n_358), .A2(n_370), .B(n_377), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_371), .B(n_323), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_358), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_366), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_368), .A2(n_323), .B(n_306), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_359), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_376), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_366), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_373), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_384), .A2(n_181), .B1(n_183), .B2(n_198), .C(n_325), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_373), .Y(n_428) );
NAND4xp25_ASAP7_75t_SL g429 ( .A(n_369), .B(n_319), .C(n_324), .D(n_198), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_379), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_394), .B(n_374), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_422), .B(n_390), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_422), .B(n_376), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_397), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_424), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_424), .Y(n_436) );
NAND2xp33_ASAP7_75t_R g437 ( .A(n_403), .B(n_369), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_403), .B(n_372), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_391), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_422), .B(n_376), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_390), .B(n_376), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_392), .B(n_376), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_398), .B(n_417), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_392), .B(n_399), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_417), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_389), .B(n_384), .Y(n_450) );
AND2x4_ASAP7_75t_SL g451 ( .A(n_403), .B(n_372), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_399), .B(n_376), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_405), .B(n_376), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_396), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_416), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_416), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_393), .B(n_385), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_405), .B(n_375), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_403), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_396), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_388), .B(n_418), .C(n_407), .Y(n_465) );
OAI21xp33_ASAP7_75t_SL g466 ( .A1(n_407), .A2(n_377), .B(n_385), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_401), .B(n_385), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_426), .B(n_375), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_386), .B(n_366), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_387), .B(n_380), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_426), .B(n_377), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_430), .Y(n_475) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_402), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_379), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_414), .B(n_364), .C(n_357), .D(n_360), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_425), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_414), .B(n_355), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_432), .B(n_386), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_475), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_470), .B(n_406), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_432), .B(n_412), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_454), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_465), .B(n_425), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_434), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_437), .A2(n_429), .B1(n_386), .B2(n_400), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_440), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_438), .Y(n_494) );
NAND2xp33_ASAP7_75t_L g495 ( .A(n_479), .B(n_404), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_450), .A2(n_386), .B1(n_415), .B2(n_413), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_448), .B(n_423), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g498 ( .A(n_466), .B(n_467), .C(n_447), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_448), .B(n_412), .Y(n_499) );
AND2x2_ASAP7_75t_SL g500 ( .A(n_481), .B(n_425), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_431), .B(n_412), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_438), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_459), .B(n_412), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_444), .B(n_415), .Y(n_505) );
AND3x2_ASAP7_75t_L g506 ( .A(n_460), .B(n_423), .C(n_410), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_481), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_459), .B(n_412), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_444), .B(n_423), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_443), .B(n_413), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_445), .Y(n_511) );
NOR2x1p5_ASAP7_75t_L g512 ( .A(n_478), .B(n_425), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_445), .B(n_410), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_460), .B(n_366), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_431), .B(n_435), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g516 ( .A1(n_449), .A2(n_408), .B1(n_420), .B2(n_410), .C(n_419), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_461), .B(n_395), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_449), .B(n_395), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_436), .B(n_404), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_469), .B(n_419), .Y(n_521) );
NOR2xp33_ASAP7_75t_SL g522 ( .A(n_473), .B(n_357), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_441), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_441), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_446), .B(n_409), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_446), .B(n_409), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_452), .B(n_409), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_468), .B(n_420), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_468), .B(n_355), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_521), .B(n_469), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_485), .A2(n_458), .B1(n_477), .B2(n_463), .C(n_474), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_485), .A2(n_453), .B1(n_452), .B2(n_469), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_500), .A2(n_451), .B(n_439), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_515), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_486), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_500), .A2(n_451), .B(n_439), .C(n_477), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_517), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_494), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_507), .A2(n_476), .B1(n_453), .B2(n_474), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_493), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_498), .B(n_442), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_488), .A2(n_463), .B(n_472), .C(n_464), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_507), .A2(n_472), .B1(n_464), .B2(n_456), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_503), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_511), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_484), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_494), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_507), .A2(n_457), .B1(n_364), .B2(n_357), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_520), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_505), .B(n_471), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_524), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_509), .B(n_433), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_509), .B(n_433), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_526), .B(n_442), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_497), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_517), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_483), .B(n_471), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_512), .A2(n_355), .B(n_364), .C(n_360), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_492), .A2(n_482), .B1(n_462), .B2(n_455), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_549), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_532), .Y(n_566) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_544), .A2(n_528), .B1(n_527), .B2(n_526), .C1(n_529), .C2(n_510), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_531), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_545), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_550), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_536), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_533), .A2(n_495), .B1(n_489), .B2(n_496), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_539), .A2(n_527), .B1(n_528), .B2(n_504), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_557), .B(n_483), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_535), .B(n_487), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_563), .A2(n_495), .B1(n_516), .B2(n_501), .C(n_514), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_531), .B(n_521), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_563), .B(n_506), .C(n_519), .Y(n_578) );
AOI211x1_ASAP7_75t_L g579 ( .A1(n_534), .A2(n_499), .B(n_518), .C(n_508), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_560), .B(n_521), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_559), .A2(n_530), .B1(n_522), .B2(n_506), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_558), .Y(n_582) );
AO22x2_ASAP7_75t_L g583 ( .A1(n_541), .A2(n_546), .B1(n_542), .B2(n_538), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_566), .A2(n_541), .B(n_546), .C(n_537), .Y(n_584) );
AOI221x1_ASAP7_75t_L g585 ( .A1(n_569), .A2(n_561), .B1(n_554), .B2(n_547), .C(n_543), .Y(n_585) );
OAI322xp33_ASAP7_75t_SL g586 ( .A1(n_576), .A2(n_562), .A3(n_556), .B1(n_555), .B2(n_552), .C1(n_548), .C2(n_513), .Y(n_586) );
OAI211xp5_ASAP7_75t_SL g587 ( .A1(n_564), .A2(n_551), .B(n_553), .C(n_427), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_568), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_579), .A2(n_514), .B1(n_523), .B2(n_525), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_583), .A2(n_525), .B1(n_523), .B2(n_502), .C(n_455), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_571), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_582), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_572), .A2(n_502), .B1(n_482), .B2(n_462), .Y(n_593) );
OA21x2_ASAP7_75t_SL g594 ( .A1(n_577), .A2(n_360), .B(n_324), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_577), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g596 ( .A1(n_584), .A2(n_572), .B1(n_581), .B2(n_573), .C(n_567), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_586), .A2(n_583), .B1(n_579), .B2(n_578), .C(n_575), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_595), .B(n_580), .Y(n_598) );
AOI221xp5_ASAP7_75t_SL g599 ( .A1(n_590), .A2(n_574), .B1(n_570), .B2(n_565), .C(n_360), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_592), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_587), .B(n_324), .C(n_183), .Y(n_601) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_587), .A2(n_181), .B(n_183), .C(n_198), .Y(n_602) );
NAND3x1_ASAP7_75t_L g603 ( .A(n_597), .B(n_593), .C(n_594), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_600), .B(n_591), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_598), .B(n_588), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_599), .B(n_589), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_605), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_604), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_608), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_607), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_610), .B(n_607), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_611), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_612), .A2(n_610), .B1(n_609), .B2(n_596), .C(n_606), .Y(n_613) );
AOI322xp5_ASAP7_75t_L g614 ( .A1(n_613), .A2(n_601), .A3(n_603), .B1(n_585), .B2(n_602), .C1(n_181), .C2(n_183), .Y(n_614) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_614), .B(n_181), .Y(n_615) );
endmodule