module fake_jpeg_19119_n_155 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_74),
.Y(n_83)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_75),
.Y(n_82)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_61),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_47),
.B1(n_62),
.B2(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_92),
.B1(n_58),
.B2(n_53),
.Y(n_97)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_65),
.B1(n_71),
.B2(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_56),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_65),
.B1(n_49),
.B2(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_79),
.B(n_52),
.C(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_98),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_83),
.B1(n_63),
.B2(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_73),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_70),
.B(n_67),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_1),
.Y(n_118)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_64),
.B1(n_60),
.B2(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_104),
.B1(n_83),
.B2(n_48),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_52),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_115),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_4),
.B(n_5),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_66),
.B1(n_91),
.B2(n_29),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_66),
.C(n_24),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_10),
.C(n_12),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_2),
.Y(n_122)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_126),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_127),
.B1(n_129),
.B2(n_106),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_113),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_117),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_110),
.C(n_32),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_120),
.B(n_130),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_141),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_142),
.B1(n_143),
.B2(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_137),
.C(n_33),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_23),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_34),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_35),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_39),
.C(n_40),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_44),
.C(n_42),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_43),
.C(n_41),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);


endmodule