module fake_jpeg_4268_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_46),
.B1(n_50),
.B2(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_19),
.B1(n_29),
.B2(n_21),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_57),
.B1(n_31),
.B2(n_23),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_18),
.CON(n_46),
.SN(n_46)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_16),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_52),
.B(n_13),
.Y(n_84)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_36),
.B1(n_41),
.B2(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_67),
.B1(n_43),
.B2(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_28),
.B1(n_20),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_56),
.B1(n_23),
.B2(n_14),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_18),
.B1(n_30),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_15),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_55),
.B1(n_50),
.B2(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_74),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_92),
.Y(n_95)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_77),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_52),
.B1(n_57),
.B2(n_47),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_93),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_92),
.B(n_77),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_115),
.B(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_118),
.B1(n_68),
.B2(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_51),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_110),
.B1(n_88),
.B2(n_69),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_63),
.B(n_59),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_60),
.B1(n_53),
.B2(n_48),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_65),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_124),
.B1(n_126),
.B2(n_110),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_133),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_72),
.B1(n_80),
.B2(n_73),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_75),
.C(n_84),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_135),
.C(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_85),
.B1(n_49),
.B2(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_83),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_87),
.B(n_48),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_136),
.B(n_97),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_140),
.B1(n_146),
.B2(n_113),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_49),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_139),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_115),
.C(n_101),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_59),
.B(n_65),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_81),
.B(n_65),
.C(n_53),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_144),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_94),
.A2(n_65),
.B(n_82),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_96),
.B(n_97),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_83),
.B1(n_58),
.B2(n_60),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_58),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_83),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_108),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_93),
.B1(n_86),
.B2(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_112),
.B(n_99),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_137),
.B1(n_130),
.B2(n_122),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_166),
.B1(n_170),
.B2(n_126),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_103),
.B1(n_119),
.B2(n_110),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_141),
.B1(n_146),
.B2(n_86),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_113),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_120),
.B(n_121),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_114),
.B(n_103),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_168),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_103),
.B1(n_114),
.B2(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_152),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_114),
.B(n_98),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_86),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_142),
.C(n_129),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_93),
.B1(n_98),
.B2(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_102),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_131),
.C(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_125),
.C(n_124),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_196),
.B1(n_186),
.B2(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_184),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_136),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_195),
.B(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_190),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_155),
.B1(n_150),
.B2(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_197),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_137),
.B1(n_145),
.B2(n_132),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_178),
.B1(n_171),
.B2(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_141),
.B1(n_102),
.B2(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_169),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_206),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_163),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_168),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_211),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_220),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_164),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_153),
.C(n_157),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_153),
.C(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_195),
.B(n_193),
.C(n_180),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_181),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_190),
.B(n_184),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_231),
.B(n_237),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_194),
.B(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_238),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_236),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_147),
.B(n_151),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_240),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_172),
.B(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_0),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_199),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_205),
.C(n_201),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_205),
.C(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_252),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_214),
.C(n_206),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_256),
.C(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_216),
.C(n_210),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_172),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_261),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_219),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_240),
.B(n_208),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_208),
.C(n_204),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_207),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_230),
.B1(n_232),
.B2(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_224),
.B(n_227),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_227),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_245),
.B(n_232),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_275),
.C(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_233),
.B1(n_226),
.B2(n_228),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_272),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_244),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_276),
.B(n_12),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_221),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_263),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_232),
.B(n_1),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_256),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_288),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_0),
.B(n_4),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_283),
.Y(n_296)
);

AOI31xp33_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_248),
.A3(n_250),
.B(n_246),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_12),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_10),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_10),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_271),
.C(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_298),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_271),
.C(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_266),
.B1(n_275),
.B2(n_270),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_289),
.B(n_8),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_5),
.C(n_6),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_5),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_311),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_288),
.B(n_281),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_295),
.C(n_294),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_312),
.B(n_301),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_315),
.Y(n_319)
);

AOI321xp33_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_317),
.A3(n_318),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_305),
.A2(n_298),
.B(n_304),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_300),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_7),
.B(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_7),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.C(n_316),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_9),
.Y(n_324)
);


endmodule