module fake_jpeg_14215_n_481 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_481);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_481;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_80),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g83 ( 
.A(n_24),
.B(n_0),
.CON(n_83),
.SN(n_83)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_1),
.B(n_2),
.Y(n_102)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_86),
.Y(n_105)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_85),
.A2(n_87),
.B(n_95),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_18),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_1),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_91),
.Y(n_132)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_93),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_43),
.Y(n_97)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_43),
.B1(n_39),
.B2(n_35),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_97),
.B(n_102),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_120),
.B1(n_138),
.B2(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_50),
.A2(n_46),
.B1(n_45),
.B2(n_48),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_106),
.A2(n_86),
.B1(n_82),
.B2(n_68),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_110),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_52),
.A2(n_42),
.B1(n_36),
.B2(n_34),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_47),
.B1(n_20),
.B2(n_44),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_54),
.A2(n_26),
.B1(n_44),
.B2(n_30),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_26),
.B1(n_30),
.B2(n_40),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_151),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_38),
.B1(n_36),
.B2(n_41),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_38),
.B1(n_48),
.B2(n_34),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_56),
.B(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_93),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_53),
.A2(n_33),
.B1(n_23),
.B2(n_21),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_23),
.B(n_42),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_140),
.A2(n_149),
.B(n_123),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_55),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_154),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_64),
.B1(n_60),
.B2(n_59),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_150),
.B1(n_141),
.B2(n_109),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_72),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_156),
.B(n_165),
.Y(n_239)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_103),
.A2(n_73),
.B1(n_66),
.B2(n_67),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_159),
.A2(n_179),
.B1(n_181),
.B2(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_163),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_87),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_164),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_101),
.B(n_72),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_200),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_92),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_98),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_80),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_97),
.B(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_173),
.B(n_14),
.Y(n_246)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_176),
.A2(n_197),
.B1(n_198),
.B2(n_133),
.Y(n_241)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_177),
.Y(n_221)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_182),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_184),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_105),
.A2(n_71),
.B1(n_63),
.B2(n_5),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_185),
.Y(n_236)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_189),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_61),
.C(n_77),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_14),
.Y(n_243)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_191),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_121),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_121),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_199),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_102),
.A2(n_61),
.B(n_6),
.C(n_8),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_9),
.C(n_13),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_108),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_196),
.A2(n_142),
.B(n_146),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_122),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_122),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_111),
.B(n_8),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_202),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_135),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_204),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_104),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_109),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_17),
.B1(n_200),
.B2(n_154),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_182),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_163),
.B1(n_204),
.B2(n_152),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_208),
.A2(n_213),
.B1(n_235),
.B2(n_238),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_160),
.B1(n_186),
.B2(n_190),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_214),
.B(n_243),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_162),
.A2(n_146),
.B(n_135),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_194),
.B(n_164),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_SL g286 ( 
.A1(n_220),
.A2(n_237),
.B(n_174),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_167),
.B(n_123),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_222),
.B(n_251),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_173),
.B(n_124),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_223),
.B(n_229),
.Y(n_275)
);

OAI22x1_ASAP7_75t_SL g225 ( 
.A1(n_160),
.A2(n_133),
.B1(n_108),
.B2(n_118),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_225),
.A2(n_241),
.B(n_177),
.C(n_195),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_226),
.A2(n_248),
.B1(n_166),
.B2(n_205),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_162),
.B(n_124),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_231),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_150),
.B1(n_141),
.B2(n_139),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_158),
.A2(n_114),
.B1(n_139),
.B2(n_118),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_158),
.A2(n_114),
.B1(n_137),
.B2(n_133),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_158),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_176),
.B1(n_175),
.B2(n_169),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_246),
.B(n_254),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_162),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_248)
);

NOR2x1_ASAP7_75t_R g250 ( 
.A(n_188),
.B(n_15),
.Y(n_250)
);

AND2x4_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_184),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_170),
.B(n_153),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_255),
.B(n_265),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_257),
.A2(n_286),
.B1(n_291),
.B2(n_238),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_157),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_261),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_158),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_208),
.B(n_171),
.C(n_164),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_272),
.C(n_216),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_263),
.B(n_231),
.C(n_236),
.Y(n_337)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_189),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_193),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_266),
.B(n_268),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_206),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_269),
.A2(n_292),
.B1(n_294),
.B2(n_252),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_215),
.B(n_201),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_271),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_232),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_185),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_218),
.Y(n_273)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_215),
.B(n_183),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_199),
.Y(n_277)
);

INVx6_ASAP7_75t_SL g278 ( 
.A(n_221),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_209),
.Y(n_279)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_210),
.B1(n_234),
.B2(n_224),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_203),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_191),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_247),
.A2(n_177),
.B(n_178),
.C(n_187),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_252),
.B(n_240),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_227),
.B(n_169),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_288),
.B(n_293),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_175),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_290),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_232),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_227),
.A2(n_214),
.B1(n_229),
.B2(n_247),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_211),
.B(n_230),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_221),
.Y(n_312)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_297),
.B(n_253),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_267),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_309),
.B1(n_310),
.B2(n_319),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_261),
.A2(n_245),
.B1(n_226),
.B2(n_219),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_314),
.B1(n_331),
.B2(n_332),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_228),
.B1(n_222),
.B2(n_235),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_228),
.B1(n_222),
.B2(n_251),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_312),
.B(n_335),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_281),
.A2(n_219),
.B1(n_222),
.B2(n_248),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_250),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_316),
.C(n_266),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_272),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_267),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_225),
.B1(n_252),
.B2(n_231),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_288),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_327),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_259),
.B(n_242),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_260),
.B(n_242),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_330),
.Y(n_353)
);

NAND2x1p5_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_236),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_260),
.A2(n_225),
.B1(n_231),
.B2(n_240),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_287),
.B(n_224),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_274),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_276),
.B(n_249),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g362 ( 
.A1(n_337),
.A2(n_284),
.B(n_220),
.Y(n_362)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_310),
.A2(n_281),
.B1(n_262),
.B2(n_268),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_349),
.B1(n_317),
.B2(n_332),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_308),
.A2(n_258),
.B(n_291),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_342),
.C(n_344),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_323),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_343),
.B(n_348),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_271),
.C(n_290),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_345),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_SL g348 ( 
.A(n_302),
.B(n_324),
.C(n_304),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_305),
.A2(n_270),
.B1(n_257),
.B2(n_269),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_297),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_354),
.C(n_355),
.Y(n_378)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_293),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_263),
.C(n_279),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_357),
.B(n_365),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_263),
.C(n_236),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_362),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_292),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_366),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_324),
.C(n_337),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_364),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_232),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_264),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_269),
.C(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_307),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_368),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_301),
.B(n_244),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_326),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_349),
.A2(n_314),
.B1(n_322),
.B2(n_306),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_370),
.A2(n_391),
.B1(n_353),
.B2(n_356),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_346),
.A2(n_309),
.B1(n_319),
.B2(n_301),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_379),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_372),
.A2(n_380),
.B1(n_381),
.B2(n_345),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_307),
.Y(n_375)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_358),
.A2(n_318),
.B1(n_304),
.B2(n_303),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_339),
.A2(n_336),
.B1(n_311),
.B2(n_325),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_336),
.B1(n_269),
.B2(n_318),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_361),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_384),
.B(n_385),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_357),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_303),
.Y(n_388)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

NOR4xp25_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_269),
.C(n_326),
.D(n_220),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_394),
.C(n_359),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_356),
.A2(n_328),
.B1(n_299),
.B2(n_313),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_396),
.A2(n_407),
.B1(n_416),
.B2(n_395),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_342),
.C(n_344),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_412),
.C(n_415),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_347),
.B1(n_353),
.B2(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_388),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_399),
.A2(n_413),
.B1(n_338),
.B2(n_393),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_341),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_401),
.Y(n_430)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_405),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_348),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_406),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_350),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_380),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_355),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_377),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_383),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_409),
.B(n_383),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_364),
.C(n_369),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_345),
.C(n_340),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_410),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_418),
.B(n_420),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_415),
.A2(n_386),
.B(n_381),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_419),
.A2(n_422),
.B(n_394),
.Y(n_437)
);

BUFx24_ASAP7_75t_SL g420 ( 
.A(n_403),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_417),
.A2(n_372),
.B(n_370),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_395),
.B(n_379),
.Y(n_423)
);

AO221x1_ASAP7_75t_L g445 ( 
.A1(n_423),
.A2(n_389),
.B1(n_401),
.B2(n_382),
.C(n_413),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_371),
.B1(n_414),
.B2(n_385),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_424),
.A2(n_425),
.B1(n_376),
.B2(n_405),
.Y(n_439)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_402),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_434),
.C(n_435),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_400),
.C(n_404),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_377),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_419),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_423),
.A2(n_376),
.B(n_411),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_438),
.A2(n_445),
.B(n_446),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_439),
.A2(n_448),
.B1(n_430),
.B2(n_422),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_382),
.B1(n_391),
.B2(n_412),
.Y(n_440)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_443),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_408),
.C(n_407),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_425),
.A2(n_354),
.B(n_299),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_392),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_447),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_424),
.A2(n_392),
.B1(n_328),
.B2(n_313),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_421),
.A2(n_300),
.B1(n_256),
.B2(n_294),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_300),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_444),
.B(n_433),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_451),
.A2(n_456),
.B(n_457),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_439),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_447),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_453),
.A2(n_459),
.B1(n_448),
.B2(n_441),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_433),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_431),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_438),
.Y(n_466)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_428),
.C(n_442),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_463),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_436),
.C(n_442),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_464),
.B(n_466),
.Y(n_471)
);

AOI322xp5_ASAP7_75t_L g467 ( 
.A1(n_455),
.A2(n_437),
.A3(n_445),
.B1(n_446),
.B2(n_443),
.C1(n_431),
.C2(n_449),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_467),
.A2(n_454),
.B(n_452),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_460),
.A2(n_432),
.B(n_428),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_468),
.A2(n_435),
.B(n_454),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_285),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_472),
.A2(n_465),
.B(n_462),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g478 ( 
.A(n_474),
.B(n_476),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_473),
.A2(n_467),
.B1(n_273),
.B2(n_256),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_475),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_471),
.C(n_469),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_478),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_480),
.B(n_244),
.Y(n_481)
);


endmodule