module fake_jpeg_12366_n_571 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_571);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_571;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_12),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_17),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_61),
.B(n_95),
.Y(n_152)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_71),
.B(n_79),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_73),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_49),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_0),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_83),
.B(n_20),
.Y(n_153)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_1),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_40),
.B1(n_50),
.B2(n_52),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_113),
.A2(n_125),
.B1(n_129),
.B2(n_28),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_30),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_115),
.B(n_126),
.Y(n_223)
);

INVx6_ASAP7_75t_SL g120 ( 
.A(n_78),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_26),
.B1(n_30),
.B2(n_43),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_27),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_149),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_52),
.B1(n_50),
.B2(n_40),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_158),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_76),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_91),
.A2(n_52),
.B1(n_50),
.B2(n_46),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_101),
.B1(n_28),
.B2(n_51),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_76),
.B(n_47),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_37),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_57),
.B(n_47),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_51),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_59),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_106),
.Y(n_191)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_176),
.B(n_190),
.Y(n_236)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_177),
.Y(n_251)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_96),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_179),
.B(n_181),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_114),
.Y(n_181)
);

OR2x4_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_46),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_182),
.B(n_122),
.Y(n_258)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_183),
.Y(n_262)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_111),
.B(n_75),
.C(n_67),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_135),
.C(n_162),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_43),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_192),
.B(n_205),
.Y(n_252)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_194),
.A2(n_204),
.B1(n_155),
.B2(n_107),
.Y(n_271)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_74),
.B1(n_98),
.B2(n_94),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_196),
.A2(n_199),
.B1(n_167),
.B2(n_127),
.Y(n_253)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_198),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_113),
.A2(n_86),
.B1(n_87),
.B2(n_77),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_122),
.A2(n_46),
.B1(n_81),
.B2(n_102),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_217),
.B1(n_218),
.B2(n_221),
.Y(n_243)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_41),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_41),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_207),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_37),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_136),
.B(n_103),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_213),
.Y(n_246)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_142),
.Y(n_212)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_141),
.B(n_68),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_214),
.Y(n_272)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_34),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_216),
.B(n_219),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_109),
.B(n_32),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_222),
.B(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_109),
.B(n_32),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_225),
.Y(n_279)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_230),
.B1(n_231),
.B2(n_122),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_151),
.A2(n_54),
.B1(n_50),
.B2(n_51),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_228),
.A2(n_45),
.B(n_42),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_161),
.B(n_2),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_229),
.B(n_35),
.Y(n_264)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_156),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_34),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_143),
.A2(n_39),
.B1(n_35),
.B2(n_28),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_23),
.B1(n_35),
.B2(n_39),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_143),
.B1(n_168),
.B2(n_112),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_244),
.B1(n_256),
.B2(n_268),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_167),
.B1(n_127),
.B2(n_157),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_245),
.A2(n_280),
.B1(n_284),
.B2(n_228),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_258),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_194),
.A2(n_157),
.B1(n_155),
.B2(n_146),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_166),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_266),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_177),
.A2(n_118),
.B1(n_116),
.B2(n_162),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_261),
.A2(n_265),
.B1(n_285),
.B2(n_198),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_274),
.C(n_210),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_197),
.A2(n_116),
.B1(n_162),
.B2(n_123),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_166),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_204),
.B(n_156),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_268),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_208),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_39),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_287),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_182),
.A2(n_147),
.B1(n_142),
.B2(n_138),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_213),
.A2(n_147),
.B1(n_23),
.B2(n_107),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_212),
.A2(n_138),
.B1(n_23),
.B2(n_42),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_175),
.B(n_188),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_220),
.B(n_174),
.Y(n_300)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_289),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_297),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_248),
.B(n_223),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_291),
.B(n_301),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_292),
.A2(n_337),
.B1(n_338),
.B2(n_270),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_295),
.A2(n_305),
.B1(n_321),
.B2(n_328),
.Y(n_346)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_241),
.Y(n_298)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_326),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_237),
.B(n_183),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_173),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_302),
.B(n_304),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_222),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_231),
.B1(n_226),
.B2(n_202),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_178),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_316),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_246),
.Y(n_339)
);

BUFx8_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_248),
.B(n_280),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_314),
.A2(n_320),
.B(n_329),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_277),
.A2(n_191),
.B(n_200),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_278),
.B(n_243),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_184),
.Y(n_317)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_317),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_230),
.Y(n_318)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_253),
.A2(n_201),
.B1(n_193),
.B2(n_211),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_319),
.A2(n_322),
.B1(n_327),
.B2(n_251),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_172),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_279),
.B(n_203),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_271),
.A2(n_266),
.B1(n_259),
.B2(n_288),
.Y(n_322)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_323),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_264),
.B(n_172),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_221),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_271),
.A2(n_218),
.B1(n_217),
.B2(n_209),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_268),
.A2(n_180),
.B1(n_200),
.B2(n_187),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_238),
.B(n_186),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_334),
.Y(n_351)
);

BUFx16f_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_331),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_271),
.A2(n_45),
.B1(n_42),
.B2(n_4),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_251),
.B1(n_275),
.B2(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_335),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_262),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_255),
.B(n_186),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_274),
.B(n_45),
.C(n_42),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_278),
.C(n_282),
.Y(n_345)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_235),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_247),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_345),
.Y(n_407)
);

AND2x6_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_246),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_339),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_342),
.A2(n_365),
.B(n_311),
.Y(n_397)
);

AO21x2_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_329),
.B(n_327),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_343),
.A2(n_356),
.B1(n_332),
.B2(n_305),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_276),
.C(n_262),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_348),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_276),
.C(n_254),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_350),
.A2(n_372),
.B1(n_293),
.B2(n_313),
.Y(n_394)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_309),
.A2(n_283),
.A3(n_269),
.B1(n_270),
.B2(n_254),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_328),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_239),
.C(n_263),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_364),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_324),
.B(n_239),
.C(n_263),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_300),
.A2(n_250),
.B(n_247),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_294),
.B(n_250),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_293),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_368),
.A2(n_313),
.B1(n_319),
.B2(n_292),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_306),
.A2(n_45),
.B(n_3),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_370),
.A2(n_311),
.B(n_312),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_295),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_322),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_374),
.A2(n_379),
.B1(n_296),
.B2(n_298),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_294),
.B(n_2),
.C(n_5),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_376),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_7),
.C(n_8),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_329),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_382),
.A2(n_397),
.B(n_362),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_394),
.Y(n_420)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_409),
.B1(n_411),
.B2(n_350),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_293),
.B(n_306),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_386),
.A2(n_405),
.B(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_387),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_359),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_399),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_314),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_314),
.Y(n_391)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_393),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_320),
.B(n_321),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_395),
.A2(n_360),
.B(n_344),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_333),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_410),
.Y(n_431)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_402),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_346),
.A2(n_291),
.B1(n_338),
.B2(n_297),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_401),
.A2(n_356),
.B1(n_343),
.B2(n_342),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_331),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_373),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_408),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_352),
.B(n_326),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_404),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_331),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_343),
.A2(n_289),
.B1(n_337),
.B2(n_307),
.Y(n_409)
);

INVx8_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_343),
.A2(n_307),
.B1(n_316),
.B2(n_299),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_323),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_414),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_7),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_416),
.Y(n_444)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_373),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_311),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_361),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_366),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_364),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_347),
.C(n_363),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_435),
.C(n_413),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_395),
.B1(n_362),
.B2(n_379),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_425),
.A2(n_427),
.B1(n_429),
.B2(n_372),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_383),
.A2(n_343),
.B1(n_365),
.B2(n_374),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_389),
.A2(n_391),
.B1(n_401),
.B2(n_394),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_409),
.B1(n_411),
.B2(n_403),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_430),
.A2(n_434),
.B1(n_10),
.B2(n_11),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_439),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_345),
.C(n_344),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_417),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_375),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_388),
.B(n_377),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_441),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_360),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_447),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_397),
.A2(n_340),
.B(n_370),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_449),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_358),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_404),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_404),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_454),
.C(n_471),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_413),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_457),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_390),
.C(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_456),
.A2(n_458),
.B1(n_461),
.B2(n_474),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_387),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_422),
.A2(n_384),
.B1(n_392),
.B2(n_400),
.Y(n_458)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_393),
.B1(n_376),
.B2(n_396),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_428),
.B(n_410),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_473),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_387),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_469),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_465),
.A2(n_468),
.B1(n_420),
.B2(n_433),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_399),
.B1(n_405),
.B2(n_406),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_444),
.B(n_446),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_355),
.C(n_380),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_410),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_472),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_9),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_423),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_475),
.A2(n_438),
.B1(n_450),
.B2(n_419),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_11),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_477),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_13),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_445),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_431),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_467),
.A2(n_426),
.B(n_449),
.Y(n_480)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g481 ( 
.A(n_459),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_481),
.B(n_500),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_437),
.C(n_439),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_487),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_469),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_437),
.C(n_426),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_474),
.B1(n_436),
.B2(n_451),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_447),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_477),
.Y(n_517)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_470),
.Y(n_494)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_494),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_457),
.B(n_420),
.C(n_433),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_499),
.Y(n_508)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_496),
.Y(n_509)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_425),
.C(n_446),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_428),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_503),
.Y(n_516)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_472),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_488),
.A2(n_464),
.B(n_436),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_512),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_476),
.Y(n_510)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_510),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_471),
.C(n_464),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_482),
.B(n_468),
.C(n_479),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_513),
.B(n_515),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_519),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_460),
.C(n_465),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_517),
.B(n_484),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_427),
.Y(n_519)
);

CKINVDCx14_ASAP7_75t_R g520 ( 
.A(n_486),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_520),
.A2(n_506),
.B1(n_504),
.B2(n_509),
.Y(n_536)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_521),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_499),
.A2(n_475),
.B1(n_431),
.B2(n_441),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_522),
.A2(n_423),
.B1(n_489),
.B2(n_501),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_512),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_527),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_495),
.Y(n_526)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_526),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_497),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_508),
.B(n_490),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_SL g546 ( 
.A(n_529),
.B(n_531),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_530),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_490),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_535),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_505),
.B(n_493),
.C(n_485),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_510),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_493),
.Y(n_535)
);

OAI21x1_ASAP7_75t_SL g547 ( 
.A1(n_536),
.A2(n_424),
.B(n_450),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_434),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_484),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_523),
.A2(n_507),
.B(n_511),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_539),
.A2(n_540),
.B(n_547),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_533),
.A2(n_501),
.B(n_516),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_525),
.A2(n_521),
.B1(n_522),
.B2(n_424),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_542),
.B(n_545),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_548),
.B(n_531),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_438),
.C(n_419),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_528),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_537),
.Y(n_551)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_551),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_541),
.A2(n_529),
.B1(n_526),
.B2(n_532),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_556),
.Y(n_558)
);

NOR2x1_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_535),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_555),
.A2(n_546),
.B(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_549),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_552),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_561),
.A2(n_555),
.B(n_540),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_562),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_553),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_564),
.Y(n_566)
);

BUFx24_ASAP7_75t_SL g567 ( 
.A(n_566),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_565),
.C(n_558),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_557),
.B(n_551),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_550),
.B(n_14),
.Y(n_570)
);

AO21x1_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_14),
.B(n_507),
.Y(n_571)
);


endmodule