module fake_jpeg_28863_n_326 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_326);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_47),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_60),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_22),
.B(n_0),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_74),
.B1(n_100),
.B2(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_86),
.B1(n_20),
.B2(n_4),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_43),
.B1(n_21),
.B2(n_30),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_79),
.B1(n_85),
.B2(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_43),
.B1(n_21),
.B2(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_91),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_43),
.B1(n_30),
.B2(n_38),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_39),
.B1(n_22),
.B2(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_34),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_32),
.B1(n_26),
.B2(n_33),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_98),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_32),
.CON(n_98),
.SN(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_26),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_108),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_25),
.B1(n_20),
.B2(n_31),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_53),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_25),
.B1(n_20),
.B2(n_3),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_20),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_25),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_67),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_18),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_66),
.B1(n_64),
.B2(n_47),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_143),
.B1(n_101),
.B2(n_110),
.Y(n_153)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_128),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_68),
.B1(n_65),
.B2(n_64),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_104),
.B1(n_111),
.B2(n_106),
.Y(n_177)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_80),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_134),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_83),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_17),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_145),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_93),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_177),
.B1(n_179),
.B2(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_105),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_154),
.B(n_180),
.Y(n_211)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_71),
.B(n_82),
.C(n_78),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_128),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_109),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_83),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_109),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_113),
.B(n_148),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_112),
.B(n_82),
.C(n_78),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_135),
.B(n_133),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_97),
.B(n_112),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_126),
.B(n_141),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_125),
.B1(n_147),
.B2(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_8),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_109),
.B1(n_111),
.B2(n_94),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_104),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_94),
.B1(n_97),
.B2(n_87),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_117),
.B1(n_146),
.B2(n_137),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_119),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_193),
.B(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_139),
.C(n_134),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_198),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_151),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_130),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_201),
.B1(n_199),
.B2(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_138),
.B1(n_127),
.B2(n_124),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_115),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_121),
.B1(n_120),
.B2(n_10),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_160),
.B(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_121),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_87),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_120),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_214),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_8),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_94),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_184),
.B(n_160),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_234),
.B(n_240),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_172),
.B1(n_177),
.B2(n_181),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_228),
.B1(n_187),
.B2(n_167),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_238),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_173),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_153),
.B1(n_175),
.B2(n_163),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_168),
.B(n_158),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_235),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_212),
.B1(n_210),
.B2(n_187),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_164),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_164),
.B(n_156),
.Y(n_240)
);

OAI322xp33_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_211),
.A3(n_180),
.B1(n_205),
.B2(n_209),
.C1(n_185),
.C2(n_206),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_242),
.Y(n_272)
);

AOI221xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_211),
.B1(n_186),
.B2(n_214),
.C(n_188),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_192),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_248),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_190),
.B(n_202),
.Y(n_244)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_261),
.B(n_252),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_255),
.B1(n_259),
.B2(n_217),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_236),
.B1(n_224),
.B2(n_219),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_167),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_215),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_215),
.B1(n_161),
.B2(n_156),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_218),
.B1(n_249),
.B2(n_261),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_220),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_165),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_165),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_216),
.C(n_227),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_161),
.B(n_162),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_266),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_227),
.C(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.C(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_226),
.C(n_225),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_240),
.B(n_221),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_270),
.B(n_271),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_229),
.B(n_222),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_254),
.B1(n_245),
.B2(n_248),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_238),
.B1(n_229),
.B2(n_230),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_229),
.B1(n_230),
.B2(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_257),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_280),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_264),
.C(n_273),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_284),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_289),
.B(n_239),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_272),
.B1(n_269),
.B2(n_250),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_247),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_251),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_275),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_268),
.B1(n_271),
.B2(n_262),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_288),
.A2(n_274),
.B1(n_270),
.B2(n_245),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_297),
.B1(n_162),
.B2(n_11),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_295),
.B(n_300),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_277),
.B1(n_286),
.B2(n_287),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_282),
.B1(n_231),
.B2(n_176),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_299),
.C(n_281),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_265),
.C(n_239),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_285),
.A2(n_231),
.B(n_155),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_285),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_307),
.C(n_9),
.Y(n_315)
);

NAND4xp25_ASAP7_75t_SL g303 ( 
.A(n_294),
.B(n_278),
.C(n_11),
.D(n_12),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_305),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_308),
.B1(n_297),
.B2(n_298),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_176),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_9),
.B(n_13),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_9),
.B(n_13),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_301),
.B1(n_293),
.B2(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_292),
.B1(n_299),
.B2(n_14),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_15),
.B(n_16),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_14),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_311),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_322),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_317),
.C(n_318),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_15),
.B(n_16),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_324),
.Y(n_326)
);


endmodule