module fake_jpeg_14387_n_487 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_50),
.Y(n_141)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_60),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_70),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_1),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

CKINVDCx6p67_ASAP7_75t_R g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_2),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_30),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_89),
.Y(n_123)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_92),
.Y(n_137)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_47),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_97),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_33),
.B1(n_42),
.B2(n_26),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_102),
.A2(n_110),
.B1(n_112),
.B2(n_116),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_33),
.B1(n_42),
.B2(n_26),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_33),
.B1(n_42),
.B2(n_26),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_46),
.B1(n_44),
.B2(n_35),
.Y(n_116)
);

AND2x4_ASAP7_75t_SL g118 ( 
.A(n_51),
.B(n_46),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_81),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_54),
.A2(n_46),
.B1(n_44),
.B2(n_49),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_25),
.B1(n_43),
.B2(n_39),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_122),
.A2(n_151),
.B1(n_79),
.B2(n_76),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_25),
.B1(n_40),
.B2(n_37),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_25),
.B1(n_49),
.B2(n_40),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_125),
.A2(n_130),
.B1(n_152),
.B2(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_48),
.B1(n_32),
.B2(n_45),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_36),
.B1(n_30),
.B2(n_45),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_48),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_19),
.Y(n_158)
);

OR2x4_ASAP7_75t_SL g149 ( 
.A(n_59),
.B(n_47),
.Y(n_149)
);

OR2x4_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_81),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_66),
.A2(n_36),
.B1(n_41),
.B2(n_34),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_61),
.A2(n_41),
.B1(n_34),
.B2(n_32),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_65),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_153),
.B(n_157),
.Y(n_228)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_97),
.B1(n_94),
.B2(n_83),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_155),
.A2(n_177),
.B1(n_197),
.B2(n_144),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_62),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_168),
.Y(n_218)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_69),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_171),
.Y(n_215)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_90),
.B(n_67),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_101),
.B(n_72),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_106),
.B(n_70),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_70),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_176),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx6_ASAP7_75t_SL g175 ( 
.A(n_115),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_58),
.Y(n_176)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_184),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_57),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_3),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_191),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_115),
.B(n_117),
.C(n_144),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_135),
.B1(n_143),
.B2(n_139),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_192),
.Y(n_216)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_88),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_107),
.B(n_81),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_3),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_195),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_118),
.B(n_56),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_103),
.A2(n_52),
.B1(n_50),
.B2(n_6),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_138),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_199),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_123),
.B(n_128),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_128),
.B(n_4),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_4),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_133),
.B1(n_109),
.B2(n_111),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_201),
.A2(n_206),
.B1(n_227),
.B2(n_232),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_210),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_109),
.B1(n_133),
.B2(n_111),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_214),
.B1(n_225),
.B2(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_160),
.A2(n_103),
.B1(n_146),
.B2(n_139),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_146),
.B1(n_132),
.B2(n_100),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_188),
.A2(n_143),
.B1(n_135),
.B2(n_113),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_100),
.B1(n_132),
.B2(n_113),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_170),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_185),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_272),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_165),
.C(n_172),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_259),
.C(n_266),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_269),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_198),
.B1(n_189),
.B2(n_193),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_243),
.A2(n_219),
.B1(n_223),
.B2(n_237),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_249),
.A2(n_250),
.B(n_251),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_186),
.B(n_184),
.C(n_178),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_191),
.B(n_168),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_204),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_252),
.B(n_253),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_228),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_177),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_222),
.B(n_158),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_258),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_176),
.C(n_171),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_191),
.B(n_194),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_267),
.B(n_217),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_163),
.B1(n_182),
.B2(n_199),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_254),
.B1(n_225),
.B2(n_241),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_219),
.A2(n_173),
.B1(n_200),
.B2(n_175),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_238),
.B1(n_207),
.B2(n_230),
.Y(n_284)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_196),
.C(n_190),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_161),
.B(n_156),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_216),
.B(n_181),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_213),
.A2(n_166),
.B1(n_174),
.B2(n_142),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_273),
.B1(n_226),
.B2(n_232),
.Y(n_281)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_271),
.B(n_274),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_215),
.A2(n_142),
.B1(n_154),
.B2(n_150),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_291),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_224),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_277),
.B(n_164),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_280),
.B(n_273),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_281),
.A2(n_290),
.B1(n_299),
.B2(n_263),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_263),
.B(n_267),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_229),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_305),
.C(n_260),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_251),
.A2(n_206),
.B1(n_226),
.B2(n_229),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_261),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_255),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_297),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_264),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_304),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_244),
.A2(n_237),
.B1(n_236),
.B2(n_212),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_236),
.B1(n_220),
.B2(n_209),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_303),
.A2(n_248),
.B1(n_247),
.B2(n_270),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_249),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_220),
.C(n_217),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_249),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_233),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_307),
.B(n_304),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_309),
.A2(n_319),
.B(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_310),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_313),
.C(n_324),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_323),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_250),
.C(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_316),
.A2(n_337),
.B1(n_303),
.B2(n_280),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_317),
.A2(n_320),
.B1(n_314),
.B2(n_321),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_294),
.A2(n_250),
.B(n_271),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_250),
.B(n_245),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_250),
.C(n_274),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_245),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_331),
.C(n_334),
.Y(n_365)
);

XOR2x2_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_278),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_328),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_279),
.Y(n_328)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_330),
.B(n_281),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_268),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_278),
.A2(n_159),
.B(n_164),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_299),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_279),
.B(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_126),
.C(n_173),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_117),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_287),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_203),
.B1(n_167),
.B2(n_238),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_239),
.Y(n_339)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_286),
.B(n_239),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_340),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_340),
.Y(n_342)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_290),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_362),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_347),
.Y(n_380)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_321),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_350),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_323),
.B(n_286),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_361),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g350 ( 
.A(n_312),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_351),
.A2(n_368),
.B1(n_369),
.B2(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_360),
.B(n_336),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_318),
.B(n_328),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_317),
.A2(n_287),
.B1(n_297),
.B2(n_276),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_318),
.B(n_302),
.Y(n_370)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_329),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_371),
.A2(n_339),
.B1(n_335),
.B2(n_334),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_357),
.A2(n_326),
.B(n_319),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_373),
.A2(n_354),
.B(n_352),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_324),
.C(n_313),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_378),
.Y(n_414)
);

AO22x1_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_355),
.B1(n_346),
.B2(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_325),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_381),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_331),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_368),
.A2(n_309),
.B1(n_315),
.B2(n_322),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_379),
.A2(n_384),
.B1(n_295),
.B2(n_293),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_330),
.Y(n_381)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_353),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_345),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_363),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_332),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_393),
.C(n_394),
.Y(n_399)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_353),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_335),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_302),
.C(n_275),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_337),
.B1(n_296),
.B2(n_292),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_395),
.A2(n_293),
.B1(n_275),
.B2(n_203),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_364),
.C(n_343),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_366),
.C(n_356),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_400),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_379),
.A2(n_357),
.B(n_363),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_401),
.A2(n_404),
.B(n_373),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_389),
.B(n_350),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_405),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_366),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_376),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_408),
.A2(n_411),
.B1(n_167),
.B2(n_126),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_390),
.B(n_296),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_230),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_367),
.C(n_369),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_396),
.C(n_377),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_383),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_413),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_418),
.B1(n_388),
.B2(n_387),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_295),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_416),
.A2(n_381),
.B(n_375),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_396),
.B1(n_385),
.B2(n_393),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_419),
.A2(n_425),
.B1(n_401),
.B2(n_402),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_420),
.A2(n_412),
.B(n_98),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_423),
.B(n_399),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_434),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_427),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_374),
.C(n_376),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_429),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_399),
.C(n_410),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_432),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_179),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_404),
.A2(n_164),
.B(n_117),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_433),
.A2(n_405),
.B(n_400),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_438),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_417),
.C(n_407),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_407),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_415),
.C(n_408),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_444),
.A2(n_445),
.B(n_449),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_422),
.A2(n_402),
.B1(n_435),
.B2(n_428),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_446),
.A2(n_15),
.B(n_11),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_423),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_421),
.A2(n_420),
.B(n_433),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_430),
.A2(n_150),
.B1(n_141),
.B2(n_98),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_10),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_5),
.B(n_8),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_451),
.A2(n_446),
.B(n_437),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_444),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_440),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_463),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_15),
.C(n_9),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_457),
.B(n_464),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_447),
.A2(n_8),
.B(n_9),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_461),
.A2(n_460),
.B(n_464),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_462),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_13),
.C(n_14),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_458),
.A2(n_445),
.B(n_451),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_470),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_472),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_455),
.B(n_441),
.Y(n_472)
);

AOI211xp5_ASAP7_75t_L g473 ( 
.A1(n_459),
.A2(n_441),
.B(n_439),
.C(n_450),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_457),
.C(n_456),
.Y(n_474)
);

AO21x1_ASAP7_75t_L g480 ( 
.A1(n_474),
.A2(n_479),
.B(n_467),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_462),
.C(n_14),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_477),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_480),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_476),
.A2(n_478),
.B(n_474),
.C(n_475),
.Y(n_481)
);

AOI31xp67_ASAP7_75t_SL g484 ( 
.A1(n_481),
.A2(n_467),
.A3(n_465),
.B(n_15),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_482),
.B(n_14),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_486),
.B(n_483),
.Y(n_487)
);


endmodule