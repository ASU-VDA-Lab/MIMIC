module fake_jpeg_32007_n_377 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_377);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_377;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_64),
.B(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_68),
.Y(n_84)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_71),
.Y(n_122)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_28),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_77),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_20),
.A2(n_11),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_9),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_6),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_0),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_42),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_0),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_81),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_42),
.B1(n_30),
.B2(n_29),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_94),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_38),
.B1(n_25),
.B2(n_23),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_39),
.B1(n_41),
.B2(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_92),
.B(n_98),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_38),
.B1(n_19),
.B2(n_18),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_23),
.B(n_25),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_110),
.B1(n_98),
.B2(n_127),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_38),
.B1(n_25),
.B2(n_41),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_105),
.B1(n_113),
.B2(n_115),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_41),
.B1(n_21),
.B2(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_116),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_43),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_24),
.B1(n_22),
.B2(n_16),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_56),
.A2(n_22),
.B1(n_16),
.B2(n_34),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_127),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_6),
.B(n_7),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_96),
.B1(n_94),
.B2(n_45),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_48),
.B(n_4),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_154),
.Y(n_184)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_141),
.Y(n_190)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_69),
.B(n_70),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_139),
.B(n_149),
.Y(n_212)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_63),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_143),
.B(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_144),
.A2(n_8),
.B1(n_176),
.B2(n_135),
.Y(n_199)
);

AO22x2_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_51),
.B1(n_59),
.B2(n_80),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_145),
.A2(n_162),
.B1(n_179),
.B2(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_84),
.B(n_71),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_150),
.A2(n_151),
.B(n_155),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_84),
.B(n_44),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_86),
.Y(n_154)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_86),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_172),
.Y(n_193)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

AO22x2_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_88),
.B1(n_90),
.B2(n_129),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_53),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_61),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_177),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_84),
.B(n_50),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_8),
.A3(n_141),
.B1(n_149),
.B2(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_53),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_176),
.A3(n_95),
.B1(n_8),
.B2(n_9),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_171),
.Y(n_207)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_6),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_104),
.B(n_66),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_68),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_134),
.Y(n_202)
);

OA22x2_ASAP7_75t_SL g179 ( 
.A1(n_95),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_88),
.B1(n_90),
.B2(n_108),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_180),
.A2(n_185),
.B1(n_187),
.B2(n_199),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_93),
.B1(n_112),
.B2(n_102),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_130),
.B1(n_132),
.B2(n_102),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_130),
.B1(n_132),
.B2(n_112),
.Y(n_187)
);

NAND2x1_ASAP7_75t_SL g228 ( 
.A(n_192),
.B(n_204),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_8),
.B1(n_149),
.B2(n_139),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_201),
.B1(n_214),
.B2(n_156),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_145),
.B1(n_179),
.B2(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_207),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_161),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_162),
.B(n_145),
.C(n_164),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_200),
.B(n_185),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_143),
.B1(n_137),
.B2(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_137),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_147),
.B1(n_163),
.B2(n_174),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_138),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_235),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_238),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_190),
.B(n_140),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_237),
.B(n_219),
.Y(n_274)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_244),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_193),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_153),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_160),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_245),
.A2(n_250),
.B1(n_204),
.B2(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_249),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_188),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_199),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_215),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_210),
.A2(n_204),
.B1(n_201),
.B2(n_180),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_211),
.B(n_237),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_187),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_218),
.C(n_189),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_242),
.B1(n_250),
.B2(n_227),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_204),
.B1(n_203),
.B2(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_256),
.A2(n_277),
.B1(n_251),
.B2(n_249),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_257),
.B(n_272),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_218),
.C(n_219),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_245),
.C(n_243),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_262),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_189),
.B(n_216),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_267),
.A2(n_232),
.B(n_230),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_226),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_274),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_215),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_233),
.B(n_198),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_278),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_228),
.A2(n_198),
.B1(n_181),
.B2(n_211),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_233),
.B(n_181),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_279),
.A2(n_228),
.B(n_243),
.Y(n_302)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_284),
.B1(n_298),
.B2(n_303),
.Y(n_314)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

AOI221xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_227),
.B1(n_247),
.B2(n_228),
.C(n_240),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_289),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_280),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_280),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_290),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_241),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_297),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_253),
.C(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_275),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_274),
.B(n_263),
.Y(n_299)
);

OA21x2_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_259),
.B(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_266),
.B(n_220),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

AOI211xp5_ASAP7_75t_SL g317 ( 
.A1(n_302),
.A2(n_256),
.B(n_277),
.C(n_264),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_311),
.C(n_315),
.Y(n_323)
);

AOI321xp33_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_260),
.A3(n_271),
.B1(n_259),
.B2(n_272),
.C(n_267),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_308),
.B(n_282),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_309),
.B(n_289),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g332 ( 
.A1(n_310),
.A2(n_317),
.B(n_301),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_272),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_257),
.C(n_261),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_261),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_319),
.C(n_287),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_281),
.B(n_236),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_276),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_254),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_331),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g326 ( 
.A(n_305),
.B(n_283),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_334),
.B1(n_337),
.B2(n_320),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_290),
.C(n_288),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_328),
.C(n_335),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_311),
.C(n_316),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_298),
.B1(n_284),
.B2(n_302),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_329),
.A2(n_270),
.B1(n_269),
.B2(n_265),
.Y(n_348)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_332),
.B(n_329),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_295),
.B1(n_297),
.B2(n_292),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_338),
.B1(n_313),
.B2(n_321),
.Y(n_340)
);

NOR3xp33_ASAP7_75t_SL g334 ( 
.A(n_304),
.B(n_300),
.C(n_303),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_295),
.C(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_336),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_312),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_313),
.A2(n_276),
.B1(n_270),
.B2(n_269),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_350),
.Y(n_359)
);

OAI31xp33_ASAP7_75t_L g341 ( 
.A1(n_332),
.A2(n_305),
.A3(n_306),
.B(n_309),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_341),
.B(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_344),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_319),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_SL g345 ( 
.A(n_334),
.B(n_308),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_345),
.A2(n_341),
.B(n_346),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_349),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_333),
.A2(n_265),
.B(n_262),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_347),
.B(n_327),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_357),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_323),
.C(n_344),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_353),
.B(n_358),
.C(n_339),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_355),
.A2(n_349),
.B(n_340),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_239),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_323),
.C(n_325),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_338),
.C(n_238),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_360),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_362),
.B(n_363),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_359),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_354),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.C(n_366),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_348),
.C(n_350),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_361),
.A2(n_355),
.B(n_358),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_360),
.B(n_365),
.C(n_366),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_362),
.C(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_371),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_SL g374 ( 
.A(n_372),
.B(n_373),
.C(n_368),
.Y(n_374)
);

NAND4xp25_ASAP7_75t_SL g373 ( 
.A(n_370),
.B(n_354),
.C(n_235),
.D(n_224),
.Y(n_373)
);

OAI311xp33_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_221),
.A3(n_222),
.B1(n_244),
.C1(n_246),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_375),
.Y(n_377)
);


endmodule