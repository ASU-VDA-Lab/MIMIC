module real_jpeg_33334_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_0),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_1),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_1),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_1),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_1),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g473 ( 
.A(n_1),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_1),
.B(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_2),
.B(n_20),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_4),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_47),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_4),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_4),
.B(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_6),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_6),
.B(n_87),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_6),
.B(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_6),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_6),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_6),
.B(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_7),
.Y(n_248)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_7),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_7),
.Y(n_516)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_8),
.B(n_79),
.Y(n_78)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_8),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_8),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_10),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_10),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_11),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_11),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_11),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_11),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_11),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_11),
.B(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_13),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_13),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_13),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g356 ( 
.A(n_13),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_13),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_13),
.B(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_13),
.B(n_476),
.Y(n_475)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_14),
.Y(n_260)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_14),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_15),
.Y(n_292)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_15),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_16),
.B(n_250),
.Y(n_249)
);

BUFx24_ASAP7_75t_L g301 ( 
.A(n_16),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_16),
.B(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_16),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_16),
.B(n_101),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_17),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_17),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_17),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_17),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_17),
.B(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_17),
.B(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_17),
.B(n_522),
.Y(n_521)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_109),
.B(n_560),
.C(n_563),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_20),
.B(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_22),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_108),
.Y(n_22)
);

NAND2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_70),
.Y(n_23)
);

OR2x6_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_70),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_48),
.Y(n_24)
);

BUFx24_ASAP7_75t_SL g566 ( 
.A(n_25),
.Y(n_566)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_41),
.CI(n_44),
.CON(n_25),
.SN(n_25)
);

MAJx2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.C(n_38),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_28),
.B(n_244),
.C(n_256),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_29),
.A2(n_30),
.B1(n_256),
.B2(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_31),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_32),
.Y(n_319)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_34),
.B(n_129),
.C(n_132),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_34),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_37),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_54),
.C(n_58),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_38),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_40),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_40),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_40),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_86),
.C(n_90),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_41),
.B(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_43),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_43),
.Y(n_188)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_43),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_45),
.A2(n_46),
.B1(n_124),
.B2(n_125),
.Y(n_194)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_46),
.B(n_125),
.C(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_47),
.B(n_301),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_63),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_52),
.B(n_145),
.C(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_52),
.B(n_234),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_63),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_96),
.C(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_54),
.A2(n_55),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_54),
.B(n_153),
.C(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_54),
.B(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2x2_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_61),
.Y(n_213)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_62),
.Y(n_311)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.C(n_105),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_71),
.A2(n_72),
.B1(n_105),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_74),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_95),
.C(n_103),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_81),
.B(n_84),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_81),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_77),
.B(n_162),
.C(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_77),
.A2(n_78),
.B1(n_166),
.B2(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_77),
.B(n_202),
.C(n_211),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_77),
.A2(n_78),
.B1(n_212),
.B2(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_85),
.B(n_106),
.C(n_107),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_86),
.B(n_90),
.Y(n_160)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_91),
.B(n_203),
.C(n_207),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_91),
.B(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2x1_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_103),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_98),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_123),
.C(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_121),
.B1(n_123),
.B2(n_141),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_99),
.B(n_354),
.C(n_356),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_99),
.A2(n_121),
.B1(n_354),
.B2(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_102),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_109),
.B(n_561),
.Y(n_560)
);

AOI21x1_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_172),
.B(n_557),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_169),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_114),
.B(n_169),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_135),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_116),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_128),
.Y(n_118)
);

XNOR2x2_ASAP7_75t_SL g214 ( 
.A(n_119),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_122),
.B(n_128),
.Y(n_215)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_125),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_125),
.B(n_252),
.Y(n_436)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_127),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_129),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_158),
.C(n_161),
.Y(n_136)
);

XNOR2x2_ASAP7_75t_L g216 ( 
.A(n_137),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B1(n_156),
.B2(n_157),
.Y(n_137)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_138),
.Y(n_228)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_143),
.B(n_146),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_145),
.B(n_363),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_153),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_154),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_153),
.A2(n_154),
.B1(n_310),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_159),
.B(n_161),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_163),
.B(n_441),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_163),
.A2(n_164),
.B1(n_441),
.B2(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_190),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_164),
.B(n_241),
.Y(n_240)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_165),
.Y(n_351)
);

INVx8_ASAP7_75t_L g519 ( 
.A(n_165),
.Y(n_519)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_268),
.B(n_552),
.Y(n_172)
);

NAND2x1_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_221),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_175),
.A2(n_554),
.B(n_555),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_218),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_177),
.B(n_556),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_214),
.C(n_216),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_179),
.B(n_214),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_195),
.C(n_200),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_193),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_182),
.B(n_185),
.Y(n_326)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_190),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_190),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_190),
.A2(n_242),
.B1(n_348),
.B2(n_349),
.Y(n_391)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_192),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_192),
.A2(n_415),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_193),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_193),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_202),
.B(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_206),
.Y(n_499)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_218),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_266),
.Y(n_221)
);

NAND2xp67_ASAP7_75t_SL g554 ( 
.A(n_222),
.B(n_266),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_230),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_224),
.B(n_227),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_230),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.C(n_261),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_232),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.C(n_240),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_233),
.B(n_240),
.Y(n_369)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_238),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_262),
.B1(n_263),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_244),
.A2(n_245),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.C(n_252),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_249),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_254),
.Y(n_476)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_259),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_373),
.B(n_543),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_333),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_330),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_271),
.A2(n_330),
.B1(n_334),
.B2(n_371),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_329),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_272),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_279),
.B(n_324),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_279),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_274),
.A2(n_275),
.B1(n_324),
.B2(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_281),
.B(n_372),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_306),
.C(n_320),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_282),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.C(n_293),
.Y(n_282)
);

XOR2x2_ASAP7_75t_L g422 ( 
.A(n_283),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_286),
.A2(n_287),
.B(n_289),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_286),
.B(n_294),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.C(n_302),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_296),
.B(n_344),
.Y(n_343)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_298),
.B(n_355),
.Y(n_354)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_300),
.A2(n_302),
.B1(n_303),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_301),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_301),
.B(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_305),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_307),
.B(n_321),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.C(n_316),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_310),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_316),
.Y(n_340)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_315),
.Y(n_439)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_329),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_330),
.B(n_550),
.C(n_551),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_371),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g544 ( 
.A(n_334),
.B(n_371),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_364),
.C(n_367),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_336),
.B(n_427),
.Y(n_426)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.C(n_361),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_338),
.B(n_362),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_418),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_346),
.B(n_360),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_342),
.A2(n_343),
.B1(n_397),
.B2(n_399),
.Y(n_396)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_352),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_347),
.A2(n_352),
.B1(n_353),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_355),
.B(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_356),
.B(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_365),
.B(n_368),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_424),
.C(n_429),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_416),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_375),
.B(n_416),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_395),
.C(n_400),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_449),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_391),
.C(n_392),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_377),
.B(n_391),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_385),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g484 ( 
.A(n_379),
.B(n_386),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_381),
.B(n_484),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_R g537 ( 
.A(n_381),
.B(n_484),
.Y(n_537)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_L g449 ( 
.A(n_396),
.B(n_400),
.Y(n_449)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_397),
.Y(n_399)
);

XOR2x2_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_406),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_406),
.C(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_411),
.C(n_415),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_407),
.A2(n_408),
.B1(n_411),
.B2(n_412),
.Y(n_446)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_420),
.C(n_422),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g545 ( 
.A1(n_425),
.A2(n_546),
.B(n_547),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_426),
.B(n_428),
.Y(n_546)
);

OAI21x1_ASAP7_75t_SL g429 ( 
.A1(n_430),
.A2(n_450),
.B(n_541),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_448),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_432),
.B(n_542),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_445),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_539),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_435),
.B(n_445),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.C(n_440),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_436),
.A2(n_437),
.B1(n_438),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_436),
.Y(n_489)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_440),
.B(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_441),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_448),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_534),
.B(n_540),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_490),
.B(n_533),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_480),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_453),
.B(n_480),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_472),
.C(n_477),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_454),
.A2(n_455),
.B1(n_501),
.B2(n_503),
.Y(n_500)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_466),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_461),
.B2(n_465),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_465),
.C(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_461),
.Y(n_465)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_472),
.A2(n_477),
.B1(n_478),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_475),
.Y(n_493)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_487),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_485),
.B2(n_486),
.Y(n_481)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_482),
.Y(n_486)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_483),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_536),
.C(n_537),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_487),
.Y(n_536)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_504),
.B(n_532),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_500),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_500),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.C(n_495),
.Y(n_492)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_529),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_494),
.Y(n_529)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_501),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_525),
.B(n_531),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_520),
.B(n_524),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_511),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_511),
.Y(n_524)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_517),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_512),
.B(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_517),
.Y(n_526)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_519),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_527),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_530),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_538),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_535),
.B(n_538),
.Y(n_540)
);

O2A1O1Ixp33_ASAP7_75t_SL g543 ( 
.A1(n_544),
.A2(n_545),
.B(n_548),
.C(n_549),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_564),
.Y(n_563)
);


endmodule