module fake_jpeg_29069_n_448 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_9),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_47),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_63),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_51),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_57),
.Y(n_140)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_15),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_73),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_77),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_13),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_89),
.Y(n_122)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_94),
.Y(n_123)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_17),
.B1(n_20),
.B2(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_99),
.A2(n_143),
.B1(n_52),
.B2(n_66),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_101),
.B(n_128),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_48),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_72),
.B1(n_67),
.B2(n_30),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_50),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_25),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_7),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_29),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_29),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_92),
.B(n_40),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_0),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_58),
.A2(n_17),
.B1(n_20),
.B2(n_44),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_148),
.B1(n_151),
.B2(n_69),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_93),
.A2(n_39),
.B1(n_19),
.B2(n_44),
.Y(n_143)
);

AND2x4_ASAP7_75t_SL g146 ( 
.A(n_68),
.B(n_44),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_8),
.B(n_9),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_46),
.A2(n_19),
.B1(n_30),
.B2(n_4),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_49),
.A2(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_12),
.B(n_11),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_153),
.Y(n_228)
);

NAND2x1_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_30),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_154),
.B(n_165),
.Y(n_236)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g242 ( 
.A1(n_156),
.A2(n_181),
.B(n_174),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_106),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_162),
.Y(n_208)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_0),
.B(n_6),
.C(n_7),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_161),
.A2(n_191),
.B(n_174),
.C(n_165),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_62),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_199),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_30),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_183),
.B1(n_198),
.B2(n_125),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_169),
.A2(n_174),
.B1(n_184),
.B2(n_147),
.Y(n_205)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_176),
.Y(n_212)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_102),
.B1(n_140),
.B2(n_98),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_96),
.B(n_6),
.C(n_7),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_139),
.C(n_133),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_100),
.B(n_6),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_180),
.Y(n_217)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_144),
.B(n_8),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_118),
.B(n_8),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_123),
.A2(n_9),
.B1(n_122),
.B2(n_99),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_9),
.B1(n_119),
.B2(n_142),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx9p33_ASAP7_75t_R g186 ( 
.A(n_97),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_113),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_101),
.B(n_131),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_190),
.Y(n_235)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_149),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_148),
.B(n_130),
.C(n_140),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_107),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_200),
.Y(n_240)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_145),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_119),
.A2(n_147),
.B1(n_145),
.B2(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_126),
.B(n_141),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_150),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_201),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_150),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_126),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_225),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_205),
.A2(n_211),
.B1(n_242),
.B2(n_198),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_164),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_215),
.B1(n_241),
.B2(n_202),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_167),
.A2(n_111),
.B1(n_127),
.B2(n_183),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_166),
.B(n_180),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_216),
.B(n_225),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_168),
.B(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_165),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_162),
.B(n_179),
.C(n_199),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_154),
.B(n_186),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_191),
.A2(n_184),
.B1(n_200),
.B2(n_172),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_165),
.B(n_184),
.Y(n_243)
);

OR2x4_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_165),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_245),
.A2(n_258),
.B(n_264),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_247),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_205),
.A2(n_184),
.B1(n_174),
.B2(n_161),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_248),
.A2(n_251),
.B1(n_268),
.B2(n_211),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_157),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_250),
.B(n_260),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_275),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_SL g258 ( 
.A(n_228),
.B(n_154),
.C(n_201),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_217),
.B(n_195),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_262),
.B1(n_220),
.B2(n_204),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_213),
.A2(n_178),
.B1(n_158),
.B2(n_170),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_163),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_263),
.B(n_276),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_197),
.B(n_192),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

AO21x2_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_197),
.B(n_189),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_206),
.A2(n_194),
.B(n_185),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_207),
.B(n_234),
.Y(n_293)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_160),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_216),
.B(n_185),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_218),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_278),
.Y(n_301)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_280),
.A2(n_305),
.B1(n_254),
.B2(n_255),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_268),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_291),
.B1(n_292),
.B2(n_268),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_298),
.C(n_306),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_220),
.B1(n_227),
.B2(n_226),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_273),
.B1(n_218),
.B2(n_258),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_236),
.C(n_224),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_275),
.A2(n_236),
.B(n_207),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_299),
.B(n_284),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_236),
.B(n_212),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_308),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_262),
.A2(n_222),
.B1(n_229),
.B2(n_234),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_229),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_209),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_259),
.C(n_266),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_247),
.A2(n_185),
.B(n_214),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_316),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_313),
.A2(n_335),
.B1(n_311),
.B2(n_312),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_294),
.A2(n_268),
.B1(n_277),
.B2(n_264),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_260),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_320),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_318),
.A2(n_331),
.B(n_332),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g319 ( 
.A1(n_295),
.A2(n_253),
.B(n_245),
.C(n_272),
.D(n_270),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_291),
.Y(n_342)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_322),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_323),
.B(n_325),
.Y(n_347)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_329),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_294),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_328),
.Y(n_343)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_330),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_265),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_333),
.B(n_284),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_271),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_337),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_285),
.A2(n_268),
.B1(n_274),
.B2(n_278),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_336),
.A2(n_281),
.B(n_293),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_269),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_288),
.C(n_298),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_348),
.C(n_351),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_339),
.A2(n_355),
.B1(n_362),
.B2(n_296),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_350),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_299),
.C(n_289),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_289),
.C(n_307),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_354),
.C(n_359),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_309),
.C(n_302),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_315),
.A2(n_296),
.B1(n_290),
.B2(n_297),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_309),
.C(n_302),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_327),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_233),
.C(n_244),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_313),
.A2(n_332),
.B1(n_336),
.B2(n_334),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_328),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_352),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_340),
.A2(n_331),
.B1(n_335),
.B2(n_326),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_368),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_346),
.A2(n_329),
.B(n_321),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_366),
.B(n_369),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_345),
.A2(n_320),
.B1(n_330),
.B2(n_324),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_349),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_371),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_297),
.B(n_210),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_378),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_256),
.B1(n_214),
.B2(n_232),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_373),
.A2(n_380),
.B1(n_382),
.B2(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_232),
.Y(n_374)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_356),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_362),
.A2(n_233),
.B(n_244),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_379),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_355),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_344),
.A2(n_155),
.B1(n_359),
.B2(n_342),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_341),
.B(n_348),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_383),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_338),
.C(n_347),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_384),
.B(n_396),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_394),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_363),
.Y(n_404)
);

AND3x1_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_350),
.C(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_393),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_367),
.B(n_352),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_351),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_353),
.C(n_358),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_381),
.C(n_382),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_398),
.B(n_364),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_375),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_406),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_394),
.C(n_387),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_372),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_408),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_363),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_410),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_385),
.B(n_366),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_413),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_397),
.A2(n_379),
.B(n_374),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_412),
.A2(n_387),
.B(n_368),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_399),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_396),
.B(n_398),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_414),
.A2(n_416),
.B(n_424),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_416),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_409),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_415),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_422),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_406),
.C(n_402),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_405),
.C(n_400),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_391),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_426),
.B(n_427),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_410),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_431),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_391),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_432),
.A2(n_418),
.B(n_404),
.Y(n_436)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_429),
.A2(n_418),
.B(n_423),
.C(n_389),
.Y(n_433)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_433),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_436),
.B(n_437),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_365),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_438),
.Y(n_441)
);

NOR3xp33_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_442),
.C(n_435),
.Y(n_443)
);

A2O1A1Ixp33_ASAP7_75t_SL g442 ( 
.A1(n_438),
.A2(n_432),
.B(n_434),
.C(n_425),
.Y(n_442)
);

NOR3xp33_ASAP7_75t_SL g445 ( 
.A(n_443),
.B(n_444),
.C(n_439),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_431),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_371),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_447),
.B(n_373),
.Y(n_448)
);


endmodule