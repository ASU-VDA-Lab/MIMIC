module fake_netlist_1_12408_n_743 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_743);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_743;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_21), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_17), .Y(n_110) );
INVx4_ASAP7_75t_R g111 ( .A(n_75), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_28), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_96), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_93), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_12), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_59), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_101), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_44), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_65), .Y(n_122) );
INVx2_ASAP7_75t_SL g123 ( .A(n_51), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_43), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_99), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_108), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_54), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_62), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_2), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_63), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_9), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_90), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_3), .Y(n_133) );
BUFx2_ASAP7_75t_SL g134 ( .A(n_104), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_55), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_70), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_58), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_83), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_89), .Y(n_140) );
INVxp33_ASAP7_75t_L g141 ( .A(n_100), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_102), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
NOR2xp67_ASAP7_75t_L g144 ( .A(n_60), .B(n_31), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_46), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_23), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_91), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_25), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
NOR2xp67_ASAP7_75t_L g151 ( .A(n_95), .B(n_35), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_107), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_50), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_112), .B(n_24), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_112), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_150), .B(n_0), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_150), .B(n_0), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_113), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_109), .B(n_1), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_130), .B(n_1), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_109), .B(n_2), .Y(n_166) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_113), .A2(n_3), .B(n_4), .Y(n_167) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_116), .A2(n_42), .B(n_105), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_123), .B(n_4), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_114), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
NOR2xp33_ASAP7_75t_R g174 ( .A(n_147), .B(n_45), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_170), .B(n_147), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_164), .B(n_141), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_161), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_173), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_160), .B(n_123), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_170), .B(n_128), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_156), .A2(n_146), .B1(n_118), .B2(n_129), .Y(n_181) );
NAND2xp33_ASAP7_75t_SL g182 ( .A(n_174), .B(n_110), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_157), .B(n_120), .Y(n_184) );
INVx6_ASAP7_75t_L g185 ( .A(n_161), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_156), .B(n_114), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_173), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_165), .B(n_115), .C(n_138), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_164), .A2(n_154), .B1(n_152), .B2(n_119), .Y(n_189) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_156), .B(n_119), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_160), .B(n_117), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_170), .B(n_125), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_164), .B(n_131), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_173), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_157), .B(n_120), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_190), .B(n_174), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_176), .B(n_164), .Y(n_204) );
INVxp67_ASAP7_75t_L g205 ( .A(n_176), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_177), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
NOR2x2_ASAP7_75t_L g209 ( .A(n_181), .B(n_166), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_197), .B(n_157), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_195), .B(n_156), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_197), .B(n_163), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_200), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_185), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_188), .B(n_165), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_175), .B(n_163), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g217 ( .A1(n_190), .A2(n_156), .B1(n_167), .B2(n_138), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_189), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_193), .B(n_170), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_195), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_163), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_183), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_190), .B(n_162), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_195), .B(n_172), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_200), .B(n_172), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_185), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_182), .B(n_162), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_192), .A2(n_172), .B(n_162), .C(n_168), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_200), .B(n_166), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_202), .B(n_166), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_194), .Y(n_234) );
BUFx6f_ASAP7_75t_SL g235 ( .A(n_196), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_196), .B(n_166), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_185), .B(n_162), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_186), .B(n_126), .Y(n_238) );
NOR2x2_ASAP7_75t_L g239 ( .A(n_181), .B(n_116), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_219), .A2(n_202), .B(n_199), .C(n_168), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_229), .A2(n_226), .B(n_223), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_225), .A2(n_199), .B(n_191), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_205), .B(n_186), .Y(n_244) );
BUFx12f_ASAP7_75t_L g245 ( .A(n_204), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_217), .B(n_186), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_211), .A2(n_189), .B1(n_179), .B2(n_201), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_228), .A2(n_168), .B(n_184), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_216), .A2(n_168), .B(n_189), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_211), .A2(n_189), .B1(n_160), .B2(n_167), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_220), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_212), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_204), .B(n_131), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_232), .B(n_160), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_213), .A2(n_198), .B(n_187), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_236), .B(n_160), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_215), .B(n_160), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_213), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_230), .A2(n_124), .B(n_142), .C(n_121), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_211), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_218), .Y(n_261) );
NOR3xp33_ASAP7_75t_SL g262 ( .A(n_209), .B(n_135), .C(n_153), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_221), .B(n_167), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_206), .A2(n_187), .B(n_178), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_206), .B(n_167), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_207), .A2(n_198), .B(n_178), .Y(n_267) );
OAI22xp5_ASAP7_75t_SL g268 ( .A1(n_239), .A2(n_167), .B1(n_134), .B2(n_140), .Y(n_268) );
OR2x6_ASAP7_75t_SL g269 ( .A(n_235), .B(n_132), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_207), .B(n_167), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_214), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_265), .A2(n_208), .B(n_234), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_268), .A2(n_217), .B1(n_235), .B2(n_203), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_249), .A2(n_231), .B(n_208), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_259), .A2(n_237), .B(n_231), .C(n_222), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_SL g276 ( .A1(n_240), .A2(n_222), .B(n_234), .C(n_233), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_233), .B1(n_235), .B2(n_238), .C(n_227), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_270), .A2(n_220), .B(n_227), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_243), .A2(n_224), .B(n_214), .C(n_121), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_269), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_241), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_240), .A2(n_144), .B(n_151), .Y(n_283) );
BUFx10_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_244), .A2(n_224), .B1(n_214), .B2(n_133), .C(n_124), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_244), .A2(n_224), .B1(n_167), .B2(n_142), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_245), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_260), .A2(n_133), .B1(n_152), .B2(n_154), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_245), .A2(n_134), .B1(n_139), .B2(n_122), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_SL g291 ( .A1(n_246), .A2(n_148), .B(n_143), .C(n_136), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_246), .A2(n_151), .B(n_144), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_242), .A2(n_145), .B(n_137), .C(n_127), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_248), .A2(n_267), .B(n_264), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_250), .A2(n_145), .B(n_137), .C(n_127), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_274), .A2(n_263), .B(n_257), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_295), .A2(n_247), .B(n_256), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_275), .A2(n_254), .B(n_262), .C(n_258), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_292), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_284), .A2(n_260), .B1(n_271), .B2(n_266), .Y(n_301) );
AOI21xp33_ASAP7_75t_L g302 ( .A1(n_283), .A2(n_136), .B(n_143), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_282), .B(n_251), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_272), .B(n_251), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
AOI222xp33_ASAP7_75t_L g307 ( .A1(n_280), .A2(n_133), .B1(n_251), .B2(n_266), .C1(n_148), .C2(n_158), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_284), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_276), .A2(n_255), .B(n_266), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_286), .A2(n_171), .B(n_158), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_276), .A2(n_158), .B(n_171), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_287), .B(n_5), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
CKINVDCx6p67_ASAP7_75t_R g316 ( .A(n_277), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_273), .A2(n_133), .B1(n_158), .B2(n_171), .Y(n_317) );
OAI21xp33_ASAP7_75t_SL g318 ( .A1(n_285), .A2(n_171), .B(n_173), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_315), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_300), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_302), .A2(n_293), .B(n_296), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_300), .Y(n_324) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_308), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_311), .A2(n_291), .B(n_294), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_312), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_308), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_310), .B(n_293), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_312), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_305), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_310), .B(n_279), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_315), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_315), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_318), .A2(n_278), .B(n_291), .Y(n_338) );
AO21x2_ASAP7_75t_L g339 ( .A1(n_302), .A2(n_290), .B(n_169), .Y(n_339) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_312), .A2(n_298), .B(n_311), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_313), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_297), .B(n_304), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_298), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_298), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_306), .A2(n_133), .B1(n_173), .B2(n_159), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_335), .B(n_297), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_336), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_330), .B(n_297), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_330), .B(n_297), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_329), .B(n_314), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_320), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_322), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_336), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_319), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_336), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_323), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_337), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
INVx5_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
INVx5_ASAP7_75t_SL g367 ( .A(n_331), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_337), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_323), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_328), .B(n_314), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_328), .B(n_303), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_325), .B(n_309), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_324), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_335), .B(n_297), .Y(n_375) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_327), .B(n_309), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_330), .B(n_313), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_333), .B(n_313), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_333), .B(n_316), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_327), .B(n_309), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_333), .B(n_316), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_325), .B(n_316), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_342), .B(n_301), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_329), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_332), .B(n_317), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_332), .B(n_133), .Y(n_388) );
INVx3_ASAP7_75t_SL g389 ( .A(n_324), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_334), .B(n_299), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_324), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_376), .B(n_345), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_376), .B(n_327), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_350), .B(n_342), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_365), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_353), .B(n_334), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_366), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_344), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_368), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_350), .B(n_344), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_352), .B(n_344), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_372), .B(n_334), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_352), .B(n_341), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_368), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_347), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_347), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_372), .B(n_307), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_371), .B(n_307), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_347), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_351), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_360), .B(n_341), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_352), .B(n_343), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_360), .B(n_343), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_377), .B(n_343), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_371), .B(n_321), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_360), .B(n_343), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_385), .B(n_345), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_351), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_390), .B(n_321), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_390), .B(n_321), .Y(n_430) );
OAI222xp33_ASAP7_75t_L g431 ( .A1(n_383), .A2(n_346), .B1(n_327), .B2(n_326), .C1(n_299), .C2(n_339), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_377), .B(n_340), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_377), .B(n_340), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_378), .B(n_340), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_381), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_351), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_381), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_378), .B(n_340), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_378), .B(n_340), .Y(n_440) );
NOR3xp33_ASAP7_75t_SL g441 ( .A(n_348), .B(n_318), .C(n_338), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_357), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_357), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_379), .B(n_340), .Y(n_444) );
AND2x4_ASAP7_75t_SL g445 ( .A(n_388), .B(n_327), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_384), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_384), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_357), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_384), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_367), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_379), .B(n_321), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_379), .B(n_331), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_382), .B(n_331), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_359), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_382), .B(n_321), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_359), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_382), .B(n_331), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_359), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_388), .B(n_331), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_348), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_398), .B(n_375), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_410), .B(n_386), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_445), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_392), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_392), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_398), .B(n_389), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_393), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_400), .B(n_386), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_433), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_393), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_410), .B(n_388), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_399), .B(n_380), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_405), .B(n_385), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_405), .B(n_361), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_432), .B(n_434), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_396), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_408), .B(n_409), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_415), .B(n_383), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_411), .B(n_420), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_408), .B(n_361), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_432), .B(n_375), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_434), .B(n_354), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_399), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_411), .B(n_354), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_445), .Y(n_487) );
AOI211xp5_ASAP7_75t_L g488 ( .A1(n_431), .A2(n_380), .B(n_389), .C(n_373), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_409), .B(n_362), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_396), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_452), .B(n_389), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_460), .B(n_362), .Y(n_492) );
AND2x4_ASAP7_75t_SL g493 ( .A(n_399), .B(n_358), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_420), .B(n_354), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_397), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_436), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_369), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_453), .B(n_369), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_397), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_453), .B(n_369), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_457), .B(n_373), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_422), .B(n_374), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_422), .B(n_374), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_457), .B(n_355), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_401), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_395), .B(n_394), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_401), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_402), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_444), .B(n_435), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_438), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_425), .B(n_355), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_460), .B(n_387), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_402), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_425), .B(n_355), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_423), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_403), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_444), .B(n_364), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_403), .B(n_387), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_404), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_459), .B(n_364), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_459), .B(n_364), .Y(n_521) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_395), .B(n_370), .Y(n_522) );
AOI222xp33_ASAP7_75t_L g523 ( .A1(n_416), .A2(n_387), .B1(n_338), .B2(n_370), .C1(n_365), .C2(n_358), .Y(n_523) );
OAI21xp33_ASAP7_75t_L g524 ( .A1(n_428), .A2(n_430), .B(n_455), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_435), .B(n_370), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_394), .B(n_358), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_439), .B(n_358), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_419), .B(n_367), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_404), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_439), .B(n_365), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_406), .B(n_387), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_450), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_438), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_427), .B(n_339), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_406), .B(n_365), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_407), .B(n_365), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_407), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_419), .B(n_367), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_412), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_440), .B(n_367), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_412), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_450), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_451), .A2(n_339), .B1(n_440), .B2(n_427), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_446), .B(n_367), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_394), .B(n_365), .Y(n_545) );
NOR2x1p5_ASAP7_75t_L g546 ( .A(n_506), .B(n_473), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_450), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_515), .B(n_429), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_480), .B(n_421), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_462), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_508), .Y(n_552) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_545), .B(n_394), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_479), .B(n_478), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_476), .B(n_429), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_510), .Y(n_556) );
AOI21xp33_ASAP7_75t_SL g557 ( .A1(n_484), .A2(n_421), .B(n_424), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_509), .B(n_446), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_464), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_509), .B(n_424), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_466), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_465), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_484), .B(n_447), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_515), .B(n_447), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_482), .B(n_449), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_467), .Y(n_566) );
BUFx3_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
NOR2xp67_ASAP7_75t_L g568 ( .A(n_506), .B(n_449), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_483), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_479), .B(n_5), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_471), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_523), .B(n_346), .C(n_456), .D(n_454), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_474), .B(n_454), .Y(n_573) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_473), .B(n_456), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_483), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_524), .B(n_458), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_513), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_482), .B(n_458), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_477), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_485), .B(n_413), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_461), .B(n_413), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_488), .B(n_441), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_545), .A2(n_326), .B(n_443), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
BUFx3_ASAP7_75t_L g585 ( .A(n_493), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_490), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_494), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_495), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_499), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_505), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_501), .B(n_448), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_461), .B(n_414), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_534), .B(n_414), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_507), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_469), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_489), .B(n_417), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_473), .B(n_417), .Y(n_597) );
NOR2xp67_ASAP7_75t_L g598 ( .A(n_506), .B(n_418), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_468), .B(n_418), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_535), .B(n_173), .C(n_443), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_426), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_540), .B(n_426), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_469), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_475), .B(n_437), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_516), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_492), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_472), .A2(n_448), .B1(n_442), .B2(n_437), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_481), .B(n_442), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_519), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_463), .B(n_6), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_534), .B(n_331), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_502), .B(n_331), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_529), .B(n_331), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_537), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_539), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_491), .B(n_339), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_541), .B(n_339), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_503), .B(n_169), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_470), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_470), .Y(n_620) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_517), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_486), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_530), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_512), .B(n_169), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_582), .A2(n_543), .B1(n_542), .B2(n_532), .C(n_487), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_574), .A2(n_522), .B(n_536), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_548), .Y(n_627) );
AOI21xp33_ASAP7_75t_SL g628 ( .A1(n_621), .A2(n_526), .B(n_528), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_595), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_546), .B(n_527), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_610), .A2(n_543), .B1(n_531), .B2(n_518), .C(n_514), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_557), .B(n_526), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_552), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_548), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_564), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_570), .A2(n_500), .B1(n_497), .B2(n_498), .C1(n_504), .C2(n_520), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_603), .Y(n_638) );
AOI32xp33_ASAP7_75t_L g639 ( .A1(n_584), .A2(n_544), .A3(n_521), .B1(n_526), .B2(n_538), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_568), .A2(n_511), .B1(n_533), .B2(n_486), .C(n_496), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_600), .B(n_544), .C(n_533), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_554), .A2(n_496), .B1(n_169), .B2(n_159), .C(n_155), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_624), .A2(n_6), .B(n_7), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_564), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_547), .A2(n_169), .B(n_159), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_555), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_551), .Y(n_647) );
AOI211xp5_ASAP7_75t_SL g648 ( .A1(n_598), .A2(n_7), .B(n_8), .C(n_9), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_606), .B(n_577), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_578), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_567), .B(n_585), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_593), .B(n_169), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_563), .A2(n_169), .B(n_159), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_607), .B(n_169), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_581), .Y(n_655) );
BUFx2_ASAP7_75t_L g656 ( .A(n_577), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_602), .A2(n_159), .B1(n_155), .B2(n_169), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_581), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_572), .A2(n_169), .B1(n_159), .B2(n_155), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_607), .B(n_159), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_592), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_593), .B(n_159), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_550), .A2(n_159), .B1(n_155), .B2(n_11), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_592), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_553), .B(n_159), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_624), .B(n_155), .C(n_10), .Y(n_666) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_597), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_618), .B(n_8), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_560), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_558), .B(n_155), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_559), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_549), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_569), .A2(n_155), .B1(n_11), .B2(n_12), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_562), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_566), .Y(n_675) );
XNOR2xp5_ASAP7_75t_L g676 ( .A(n_561), .B(n_10), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_628), .A2(n_633), .B1(n_625), .B2(n_656), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_670), .Y(n_678) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_634), .A2(n_575), .B1(n_623), .B2(n_587), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_627), .B(n_576), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_636), .Y(n_681) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_676), .A2(n_556), .A3(n_576), .B(n_565), .Y(n_682) );
OAI31xp33_ASAP7_75t_L g683 ( .A1(n_648), .A2(n_616), .A3(n_611), .B(n_599), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_632), .A2(n_573), .B1(n_571), .B2(n_590), .C(n_594), .Y(n_684) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_654), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_644), .Y(n_686) );
AOI311xp33_ASAP7_75t_L g687 ( .A1(n_649), .A2(n_579), .A3(n_605), .B(n_586), .C(n_615), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_659), .B(n_611), .C(n_588), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_635), .A2(n_614), .B1(n_609), .B2(n_589), .C(n_601), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_655), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g691 ( .A1(n_648), .A2(n_583), .B(n_617), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_629), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_630), .B(n_591), .Y(n_693) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_651), .B(n_622), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_673), .A2(n_617), .B(n_613), .Y(n_695) );
AOI332xp33_ASAP7_75t_L g696 ( .A1(n_650), .A2(n_619), .A3(n_620), .B1(n_613), .B2(n_608), .B3(n_604), .C1(n_596), .C2(n_580), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_647), .B(n_612), .Y(n_697) );
AOI31xp33_ASAP7_75t_L g698 ( .A1(n_668), .A2(n_14), .A3(n_15), .B(n_16), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_639), .A2(n_155), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_658), .Y(n_700) );
AOI21xp33_ASAP7_75t_SL g701 ( .A1(n_631), .A2(n_14), .B(n_18), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_673), .A2(n_18), .B(n_19), .C(n_20), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g703 ( .A1(n_667), .A2(n_155), .B1(n_20), .B2(n_21), .C1(n_22), .C2(n_19), .Y(n_703) );
NAND2x1_ASAP7_75t_L g704 ( .A(n_626), .B(n_155), .Y(n_704) );
OAI221xp5_ASAP7_75t_SL g705 ( .A1(n_637), .A2(n_22), .B1(n_111), .B2(n_27), .C(n_29), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_694), .B(n_661), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_677), .A2(n_640), .B1(n_664), .B2(n_671), .C(n_674), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_701), .A2(n_643), .B(n_668), .C(n_665), .Y(n_708) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_683), .B(n_645), .C(n_642), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_687), .A2(n_641), .B1(n_638), .B2(n_675), .C(n_663), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g711 ( .A1(n_685), .A2(n_646), .B1(n_660), .B2(n_652), .C1(n_672), .C2(n_662), .Y(n_711) );
NAND4xp75_ASAP7_75t_L g712 ( .A(n_699), .B(n_643), .C(n_653), .D(n_652), .Y(n_712) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_679), .A2(n_657), .B(n_666), .C(n_669), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_682), .A2(n_657), .B1(n_111), .B2(n_32), .C(n_33), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_684), .A2(n_26), .B1(n_30), .B2(n_34), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_696), .A2(n_36), .B(n_37), .C(n_38), .Y(n_716) );
AOI221x1_ASAP7_75t_L g717 ( .A1(n_695), .A2(n_39), .B1(n_40), .B2(n_41), .C(n_47), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_692), .B(n_48), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g719 ( .A1(n_703), .A2(n_49), .B(n_52), .C(n_53), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_693), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_707), .B(n_705), .C(n_702), .D(n_691), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_716), .B(n_692), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_720), .B(n_678), .Y(n_723) );
NAND5xp2_ASAP7_75t_L g724 ( .A(n_714), .B(n_685), .C(n_678), .D(n_689), .E(n_698), .Y(n_724) );
NOR4xp25_ASAP7_75t_L g725 ( .A(n_709), .B(n_681), .C(n_686), .D(n_690), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_708), .A2(n_704), .B(n_680), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g727 ( .A(n_713), .B(n_711), .C(n_719), .D(n_717), .Y(n_727) );
OAI222xp33_ASAP7_75t_L g728 ( .A1(n_722), .A2(n_710), .B1(n_706), .B2(n_715), .C1(n_700), .C2(n_718), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_723), .Y(n_729) );
NOR3xp33_ASAP7_75t_L g730 ( .A(n_727), .B(n_712), .C(n_688), .Y(n_730) );
NAND3xp33_ASAP7_75t_SL g731 ( .A(n_725), .B(n_697), .C(n_57), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_729), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_730), .A2(n_721), .B1(n_726), .B2(n_724), .Y(n_733) );
NAND4xp75_ASAP7_75t_L g734 ( .A(n_728), .B(n_56), .C(n_61), .D(n_64), .Y(n_734) );
AOI221xp5_ASAP7_75t_SL g735 ( .A1(n_733), .A2(n_731), .B1(n_67), .B2(n_68), .C(n_69), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_732), .Y(n_736) );
OA22x2_ASAP7_75t_L g737 ( .A1(n_736), .A2(n_734), .B1(n_72), .B2(n_73), .Y(n_737) );
AOI22x1_ASAP7_75t_L g738 ( .A1(n_735), .A2(n_66), .B1(n_74), .B2(n_76), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_737), .A2(n_77), .B1(n_78), .B2(n_80), .Y(n_739) );
OA22x2_ASAP7_75t_L g740 ( .A1(n_738), .A2(n_82), .B1(n_85), .B2(n_86), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_740), .A2(n_87), .B1(n_92), .B2(n_94), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_741), .A2(n_739), .B(n_103), .Y(n_742) );
AOI21xp33_ASAP7_75t_SL g743 ( .A1(n_742), .A2(n_98), .B(n_106), .Y(n_743) );
endmodule