module fake_jpeg_8617_n_282 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_23),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_46),
.A3(n_30),
.B1(n_17),
.B2(n_28),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_54),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_63),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_20),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_62),
.B1(n_18),
.B2(n_19),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_25),
.B(n_19),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_19),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_78),
.C(n_16),
.Y(n_105)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

OR2x4_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_70),
.B(n_75),
.CI(n_78),
.CON(n_100),
.SN(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_81),
.B1(n_42),
.B2(n_41),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_16),
.B1(n_32),
.B2(n_33),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_36),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_42),
.B1(n_41),
.B2(n_36),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_88),
.B1(n_32),
.B2(n_64),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_42),
.B1(n_21),
.B2(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_97),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_92),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_84),
.B(n_83),
.C(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_106),
.B1(n_113),
.B2(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_105),
.B(n_32),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_66),
.B1(n_73),
.B2(n_38),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_55),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_111),
.Y(n_137)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_109),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_73),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_48),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_54),
.B1(n_48),
.B2(n_64),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_68),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_118),
.B(n_31),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_98),
.B(n_111),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_79),
.B(n_77),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_140),
.B(n_126),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_94),
.B1(n_113),
.B2(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_141),
.B1(n_110),
.B2(n_17),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_69),
.B(n_31),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_21),
.B1(n_28),
.B2(n_22),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_138),
.B1(n_97),
.B2(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_17),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_72),
.B1(n_86),
.B2(n_65),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_95),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_66),
.B(n_71),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_144),
.B1(n_165),
.B2(n_141),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_151),
.B(n_160),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_92),
.B1(n_100),
.B2(n_107),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_157),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_119),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_162),
.B1(n_166),
.B2(n_17),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_140),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_100),
.C(n_15),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_119),
.C(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_159),
.C(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_100),
.C(n_38),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_107),
.C(n_51),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_13),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_163),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_109),
.B1(n_110),
.B2(n_53),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_128),
.B1(n_116),
.B2(n_117),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_10),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_51),
.C(n_109),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_51),
.C(n_24),
.Y(n_192)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_143),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_162),
.A2(n_131),
.B1(n_133),
.B2(n_132),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_189),
.B1(n_169),
.B2(n_163),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_184),
.B1(n_186),
.B2(n_26),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_118),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_177),
.C(n_192),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_151),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_134),
.B1(n_135),
.B2(n_129),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_182),
.B1(n_194),
.B2(n_0),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_122),
.B1(n_53),
.B2(n_49),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_122),
.B1(n_29),
.B2(n_27),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_49),
.B1(n_51),
.B2(n_29),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_24),
.B(n_26),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_152),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_165),
.B1(n_150),
.B2(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_199),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_161),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_156),
.C(n_168),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_206),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_211),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_29),
.C(n_27),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_27),
.C(n_26),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_174),
.B1(n_193),
.B2(n_178),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_188),
.B1(n_174),
.B2(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_218),
.A2(n_225),
.B1(n_9),
.B2(n_13),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

OAI322xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_193),
.A3(n_198),
.B1(n_171),
.B2(n_197),
.C1(n_195),
.C2(n_170),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_232),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_190),
.CI(n_192),
.CON(n_222),
.SN(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_181),
.B1(n_178),
.B2(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_206),
.B1(n_210),
.B2(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_8),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_200),
.C(n_202),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_242),
.C(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_213),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_232),
.C(n_219),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_216),
.B1(n_211),
.B2(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_226),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_8),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_15),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_8),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_223),
.C(n_224),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_7),
.B(n_13),
.Y(n_244)
);

OAI321xp33_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_11),
.A3(n_12),
.B1(n_6),
.B2(n_5),
.C(n_4),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_217),
.B1(n_226),
.B2(n_11),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_219),
.B(n_236),
.C(n_245),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_253),
.B(n_241),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_12),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_254),
.C(n_235),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_6),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_234),
.C1(n_249),
.C2(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_234),
.C(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_271),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_254),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_259),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_261),
.B(n_249),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_275),
.B(n_276),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_2),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_267),
.B(n_269),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_274),
.C(n_2),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_277),
.C(n_3),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_3),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);


endmodule