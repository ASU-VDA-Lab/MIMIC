module fake_jpeg_18627_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_31),
.B1(n_18),
.B2(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_46),
.B1(n_44),
.B2(n_35),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_67),
.Y(n_89)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_70),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_31),
.B1(n_18),
.B2(n_29),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_41),
.B1(n_34),
.B2(n_29),
.Y(n_97)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_44),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_21),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_76),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_84),
.Y(n_125)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_43),
.CON(n_79),
.SN(n_79)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_81),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_44),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_33),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_31),
.B1(n_18),
.B2(n_47),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_97),
.B1(n_98),
.B2(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_21),
.B(n_19),
.C(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_96),
.B(n_108),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_101),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_19),
.B(n_16),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_41),
.C(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_105),
.Y(n_140)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_42),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_113),
.B1(n_39),
.B2(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_68),
.B(n_42),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_42),
.C(n_39),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_73),
.B1(n_68),
.B2(n_35),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_126),
.B1(n_133),
.B2(n_136),
.Y(n_152)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_105),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_82),
.B1(n_106),
.B2(n_93),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_20),
.B1(n_26),
.B2(n_34),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_143),
.B1(n_109),
.B2(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_113),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_39),
.B1(n_26),
.B2(n_20),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_82),
.A2(n_39),
.B1(n_60),
.B2(n_24),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_82),
.A2(n_60),
.B1(n_24),
.B2(n_33),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_108),
.B(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_150),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_149),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_140),
.B1(n_120),
.B2(n_138),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_106),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_159),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_81),
.C(n_88),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_164),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_110),
.B1(n_99),
.B2(n_102),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_162),
.B1(n_177),
.B2(n_136),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_100),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_176),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_120),
.B1(n_118),
.B2(n_122),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_89),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_160),
.B(n_161),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_81),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_99),
.B1(n_90),
.B2(n_111),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_178),
.B(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_96),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_80),
.C(n_94),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_166),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_94),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_112),
.C(n_27),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_95),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_27),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_171),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_25),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_25),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_116),
.A2(n_109),
.B1(n_76),
.B2(n_33),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_112),
.B1(n_23),
.B2(n_24),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_203),
.B1(n_208),
.B2(n_152),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_182),
.A2(n_184),
.B(n_186),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_144),
.B(n_138),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_188),
.B1(n_197),
.B2(n_199),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_134),
.B(n_138),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_123),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_133),
.B1(n_115),
.B2(n_130),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_205),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_145),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_194),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_122),
.B(n_107),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_200),
.B(n_178),
.Y(n_229)
);

OAI22x1_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_118),
.B1(n_91),
.B2(n_17),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_117),
.B1(n_118),
.B2(n_128),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_114),
.B(n_17),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_137),
.B1(n_25),
.B2(n_23),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_162),
.B1(n_172),
.B2(n_147),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_164),
.B1(n_170),
.B2(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_147),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_137),
.B1(n_91),
.B2(n_128),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_8),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_194),
.B1(n_3),
.B2(n_4),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_221),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_224),
.B1(n_188),
.B2(n_179),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_165),
.C(n_161),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_210),
.C(n_198),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_163),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_169),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_187),
.Y(n_227)
);

XOR2x2_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_184),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_167),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_233),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_146),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_160),
.B(n_3),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_201),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_182),
.B1(n_200),
.B2(n_195),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_9),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_215),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_243),
.C(n_246),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_250),
.B(n_214),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_202),
.C(n_185),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_254),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_202),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_202),
.C(n_201),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_255),
.C(n_218),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_207),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_179),
.B1(n_194),
.B2(n_4),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_224),
.B1(n_214),
.B2(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_257),
.B(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_264),
.B1(n_267),
.B2(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_274),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_216),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_217),
.B1(n_219),
.B2(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_228),
.C(n_237),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_243),
.C(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_233),
.C(n_228),
.Y(n_269)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_273),
.B1(n_242),
.B2(n_6),
.Y(n_288)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_240),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_214),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_240),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_285),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_244),
.B(n_250),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_289),
.B(n_274),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_242),
.B(n_7),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_11),
.C(n_7),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_277),
.C(n_9),
.Y(n_302)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_267),
.B1(n_264),
.B2(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_300),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_298),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_299),
.B1(n_283),
.B2(n_290),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_281),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_272),
.B1(n_266),
.B2(n_273),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_268),
.B1(n_265),
.B2(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_10),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_15),
.B1(n_10),
.B2(n_12),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_301),
.C(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_310),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_303),
.B1(n_297),
.B2(n_294),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_278),
.C(n_285),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_284),
.C(n_280),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_302),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_316),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_301),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_293),
.Y(n_316)
);

OA21x2_ASAP7_75t_SL g321 ( 
.A1(n_318),
.A2(n_299),
.B(n_308),
.Y(n_321)
);

OAI211xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_315),
.B(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.C(n_320),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_320),
.B1(n_282),
.B2(n_14),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_12),
.B(n_14),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_14),
.C(n_15),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_1),
.Y(n_328)
);


endmodule