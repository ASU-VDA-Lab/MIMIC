module fake_jpeg_2949_n_222 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_11),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_1),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_13),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_27),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_77),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_66),
.Y(n_98)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_72),
.B1(n_58),
.B2(n_63),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_57),
.B(n_77),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_71),
.Y(n_113)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_58),
.B1(n_67),
.B2(n_63),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_79),
.B1(n_73),
.B2(n_64),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_69),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2x1p5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_82),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_107),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_68),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_78),
.B1(n_80),
.B2(n_85),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_113),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_59),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_64),
.A3(n_62),
.B1(n_75),
.B2(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_80),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_61),
.B1(n_59),
.B2(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_0),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_30),
.B1(n_51),
.B2(n_50),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_106),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_126),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g125 ( 
.A(n_101),
.Y(n_125)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_70),
.C(n_53),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_136),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_78),
.B1(n_53),
.B2(n_70),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_85),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_108),
.B1(n_91),
.B2(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_61),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_28),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_99),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_143),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_116),
.B(n_93),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_125),
.B(n_120),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_144),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_105),
.B1(n_61),
.B2(n_59),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_148),
.B1(n_20),
.B2(n_46),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_99),
.B1(n_3),
.B2(n_4),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_154),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_2),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_R g167 ( 
.A(n_157),
.B(n_3),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_2),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_8),
.Y(n_183)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_24),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_4),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_125),
.B(n_134),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_173),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_173),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_52),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_163),
.C(n_156),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_31),
.B(n_47),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_182),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_6),
.B(n_7),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_168),
.B1(n_166),
.B2(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_179),
.Y(n_192)
);

AOI21x1_ASAP7_75t_SL g179 ( 
.A1(n_153),
.A2(n_33),
.B(n_45),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_19),
.B(n_42),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_140),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_162),
.C(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_176),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_193),
.A2(n_177),
.B1(n_166),
.B2(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_170),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_164),
.B(n_170),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_187),
.C(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_194),
.C(n_190),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_197),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_154),
.B1(n_10),
.B2(n_11),
.Y(n_205)
);

AOI31xp67_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_9),
.A3(n_10),
.B(n_13),
.Y(n_207)
);

OAI322xp33_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_211),
.A3(n_204),
.B1(n_36),
.B2(n_18),
.C1(n_39),
.C2(n_40),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_203),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_37),
.B(n_41),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_38),
.B(n_48),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_212),
.B(n_213),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_213),
.B1(n_210),
.B2(n_17),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_216),
.B(n_14),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_16),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_16),
.Y(n_222)
);


endmodule