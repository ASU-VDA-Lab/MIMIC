module fake_ariane_15_n_1021 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1021);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1021;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx2_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_97),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_129),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_48),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_148),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_56),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_161),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_147),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_92),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_20),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_150),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_118),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_146),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_143),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_84),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_198),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_115),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_9),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_90),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_59),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_0),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_55),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_18),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_47),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_30),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_142),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_57),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_60),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_26),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_138),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_13),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_42),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_67),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_53),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_43),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_14),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_164),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_80),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_119),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_26),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_177),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_163),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_79),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_188),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_104),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_3),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_113),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_193),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_189),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_185),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_186),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_50),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_180),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_289),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_289),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_216),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_217),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_226),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_226),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_210),
.B(n_0),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_219),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_243),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_243),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_228),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_242),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_246),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_214),
.B(n_1),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_252),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_255),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_240),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_258),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_266),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_211),
.B(n_1),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_275),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_261),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_280),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_284),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_255),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_222),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_222),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_222),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_213),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_290),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_293),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_224),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_270),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_234),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_291),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_299),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_301),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_300),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_291),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_313),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_313),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_325),
.B(n_285),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_306),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_314),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_310),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_209),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_319),
.A2(n_292),
.B(n_259),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_220),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_336),
.Y(n_371)
);

OAI21x1_ASAP7_75t_L g372 ( 
.A1(n_328),
.A2(n_263),
.B(n_250),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_297),
.B(n_268),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_315),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_318),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_207),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_317),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_207),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_311),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_320),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_323),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_323),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_320),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_294),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_294),
.B(n_281),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_334),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_296),
.B(n_327),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_347),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_296),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

OR2x6_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_354),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

AO21x2_ASAP7_75t_L g410 ( 
.A1(n_372),
.A2(n_283),
.B(n_269),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_396),
.B(n_329),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

AO21x2_ASAP7_75t_L g414 ( 
.A1(n_372),
.A2(n_358),
.B(n_356),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_362),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_329),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_331),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_331),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_383),
.B1(n_368),
.B2(n_379),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_332),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_392),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_368),
.B(n_332),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_L g427 ( 
.A1(n_376),
.A2(n_341),
.B1(n_340),
.B2(n_231),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_380),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_355),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_340),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_379),
.Y(n_435)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_281),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_354),
.B(n_341),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_2),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_354),
.B(n_288),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_238),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_208),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_212),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_349),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_215),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_400),
.B(n_218),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

BUFx8_ASAP7_75t_SL g453 ( 
.A(n_348),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_365),
.B(n_221),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_367),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_400),
.B(n_223),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_366),
.B(n_225),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_400),
.B(n_262),
.Y(n_458)
);

AND3x2_ASAP7_75t_L g459 ( 
.A(n_364),
.B(n_2),
.C(n_3),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_378),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_349),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_370),
.B(n_262),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_370),
.B(n_4),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_371),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_349),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_384),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_405),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_403),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_227),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_371),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_373),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_424),
.B(n_393),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_424),
.A2(n_408),
.B1(n_420),
.B2(n_470),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_452),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_452),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_383),
.B1(n_369),
.B2(n_376),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_418),
.B(n_399),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_401),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_420),
.B(n_363),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_421),
.B(n_401),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_377),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_408),
.B(n_393),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_419),
.B(n_381),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_423),
.B(n_388),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_433),
.B(n_394),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_416),
.A2(n_425),
.B(n_449),
.C(n_444),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_408),
.A2(n_397),
.B1(n_391),
.B2(n_375),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_426),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_428),
.B(n_383),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_350),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_408),
.A2(n_386),
.B1(n_398),
.B2(n_361),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_413),
.B(n_351),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_470),
.A2(n_361),
.B1(n_369),
.B2(n_385),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_435),
.B(n_403),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_429),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_448),
.B(n_385),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_469),
.A2(n_369),
.B1(n_374),
.B2(n_349),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_455),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_458),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_438),
.B(n_412),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_357),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_467),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_406),
.B(n_374),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_5),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_448),
.B(n_422),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_440),
.B(n_6),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_415),
.A2(n_369),
.B1(n_287),
.B2(n_286),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_446),
.B(n_230),
.C(n_229),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_432),
.A2(n_235),
.B(n_232),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_427),
.B(n_236),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_415),
.B(n_237),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

O2A1O1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_460),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_415),
.A2(n_282),
.B1(n_276),
.B2(n_274),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_469),
.A2(n_429),
.B1(n_465),
.B2(n_478),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

CKINVDCx11_ASAP7_75t_R g536 ( 
.A(n_407),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_469),
.A2(n_262),
.B1(n_267),
.B2(n_271),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_407),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_461),
.A2(n_273),
.B1(n_264),
.B2(n_257),
.Y(n_540)
);

O2A1O1Ixp5_ASAP7_75t_L g541 ( 
.A1(n_434),
.A2(n_267),
.B(n_262),
.C(n_12),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_8),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_407),
.B(n_10),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_434),
.A2(n_241),
.B(n_239),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_12),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_464),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_456),
.B(n_244),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_469),
.A2(n_267),
.B1(n_262),
.B2(n_256),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_441),
.B(n_245),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_441),
.B(n_247),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_453),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_466),
.B(n_248),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_411),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_471),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_439),
.B(n_249),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_454),
.B(n_253),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_439),
.B(n_262),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_469),
.A2(n_267),
.B1(n_262),
.B2(n_15),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_469),
.A2(n_267),
.B1(n_14),
.B2(n_16),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_457),
.B(n_267),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_507),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_519),
.B(n_417),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_494),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_499),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_518),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_484),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_494),
.B(n_474),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_536),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_553),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_483),
.A2(n_436),
.B1(n_451),
.B2(n_472),
.Y(n_577)
);

INVx6_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_488),
.B(n_490),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_486),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_556),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

NOR2xp67_ASAP7_75t_L g584 ( 
.A(n_539),
.B(n_474),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_503),
.B(n_475),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_497),
.B(n_458),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_482),
.B(n_521),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_514),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_492),
.B(n_458),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_501),
.B(n_453),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_543),
.Y(n_594)
);

A2O1A1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_563),
.A2(n_479),
.B(n_477),
.C(n_447),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_522),
.B(n_458),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_509),
.B(n_477),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_SL g600 ( 
.A(n_491),
.B(n_459),
.C(n_479),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_517),
.B(n_458),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_506),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_489),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

AO22x1_ASAP7_75t_L g606 ( 
.A1(n_559),
.A2(n_437),
.B1(n_458),
.B2(n_436),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_521),
.Y(n_608)
);

AND3x1_ASAP7_75t_SL g609 ( 
.A(n_516),
.B(n_13),
.C(n_16),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_515),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_523),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_515),
.B(n_447),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_517),
.B(n_437),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_500),
.B(n_480),
.Y(n_614)
);

NOR3xp33_ASAP7_75t_SL g615 ( 
.A(n_496),
.B(n_17),
.C(n_18),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_493),
.B(n_437),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_523),
.B(n_436),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_515),
.B(n_437),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

INVx3_ASAP7_75t_SL g621 ( 
.A(n_561),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_520),
.B(n_437),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_520),
.B(n_437),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_495),
.B(n_480),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_515),
.B(n_436),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_546),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_595),
.A2(n_541),
.B(n_562),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_586),
.Y(n_631)
);

AOI221x1_ASAP7_75t_L g632 ( 
.A1(n_595),
.A2(n_546),
.B1(n_542),
.B2(n_544),
.C(n_530),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_596),
.A2(n_541),
.B(n_513),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_579),
.B(n_487),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_613),
.A2(n_513),
.B(n_564),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_622),
.A2(n_548),
.B(n_560),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_624),
.A2(n_542),
.A3(n_554),
.B(n_552),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_618),
.A2(n_562),
.B(n_534),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_601),
.A2(n_534),
.B(n_563),
.Y(n_639)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_591),
.A2(n_508),
.B(n_538),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_587),
.A2(n_414),
.B(n_526),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_551),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_577),
.A2(n_549),
.B(n_472),
.Y(n_643)
);

NAND2x1_ASAP7_75t_L g644 ( 
.A(n_610),
.B(n_557),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_627),
.A2(n_549),
.B(n_472),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_627),
.A2(n_468),
.B(n_538),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_572),
.B(n_504),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_583),
.B(n_529),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_612),
.A2(n_468),
.B(n_550),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_625),
.A2(n_414),
.B(n_499),
.Y(n_650)
);

NOR2x1_ASAP7_75t_L g651 ( 
.A(n_584),
.B(n_557),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_568),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_583),
.B(n_487),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_623),
.B(n_535),
.Y(n_654)
);

AO31x2_ASAP7_75t_L g655 ( 
.A1(n_629),
.A2(n_528),
.A3(n_410),
.B(n_540),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_612),
.A2(n_468),
.B(n_550),
.Y(n_656)
);

OA21x2_ASAP7_75t_L g657 ( 
.A1(n_604),
.A2(n_525),
.B(n_410),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_603),
.A2(n_532),
.B(n_414),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_598),
.A2(n_533),
.B(n_463),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_603),
.A2(n_410),
.B(n_535),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_604),
.A2(n_555),
.B(n_535),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_607),
.A2(n_555),
.B(n_535),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_574),
.B(n_555),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_588),
.B(n_608),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_565),
.A2(n_555),
.B1(n_442),
.B2(n_431),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_588),
.A2(n_442),
.B1(n_431),
.B2(n_411),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_569),
.A2(n_442),
.B1(n_431),
.B2(n_411),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_607),
.Y(n_668)
);

AO31x2_ASAP7_75t_L g669 ( 
.A1(n_582),
.A2(n_442),
.A3(n_431),
.B(n_463),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_570),
.A2(n_463),
.B(n_442),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_599),
.A2(n_431),
.B(n_463),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_597),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_615),
.A2(n_463),
.B(n_19),
.C(n_20),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_582),
.A2(n_267),
.A3(n_100),
.B(n_101),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_589),
.B(n_46),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_573),
.A2(n_17),
.B(n_19),
.Y(n_676)
);

AO31x2_ASAP7_75t_L g677 ( 
.A1(n_590),
.A2(n_102),
.A3(n_205),
.B(n_203),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_588),
.B(n_21),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_580),
.B(n_21),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_574),
.B(n_22),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_574),
.B(n_611),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_581),
.B(n_22),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_614),
.A2(n_616),
.B(n_626),
.C(n_600),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_567),
.B(n_23),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_590),
.A2(n_99),
.B(n_200),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_567),
.B(n_23),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_620),
.A2(n_103),
.B(n_197),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_589),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_647),
.A2(n_594),
.B1(n_602),
.B2(n_578),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_SL g690 ( 
.A1(n_676),
.A2(n_609),
.B(n_592),
.C(n_593),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_652),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_652),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_681),
.B(n_566),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_650),
.A2(n_660),
.B(n_641),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_642),
.A2(n_617),
.B(n_605),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_642),
.A2(n_617),
.B(n_605),
.Y(n_696)
);

BUFx2_ASAP7_75t_SL g697 ( 
.A(n_678),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_668),
.Y(n_698)
);

OA21x2_ASAP7_75t_L g699 ( 
.A1(n_632),
.A2(n_641),
.B(n_650),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_661),
.A2(n_619),
.B(n_606),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_653),
.A2(n_578),
.B1(n_621),
.B2(n_609),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_663),
.B(n_617),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_659),
.B(n_568),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_631),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_664),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_648),
.A2(n_638),
.B1(n_676),
.B2(n_634),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_672),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_665),
.A2(n_610),
.A3(n_619),
.B(n_571),
.Y(n_708)
);

OA21x2_ASAP7_75t_L g709 ( 
.A1(n_630),
.A2(n_571),
.B(n_568),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_678),
.B(n_578),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_662),
.A2(n_571),
.B(n_568),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_659),
.B(n_571),
.Y(n_712)
);

NAND2x1p5_ASAP7_75t_L g713 ( 
.A(n_664),
.B(n_585),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_680),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_SL g715 ( 
.A1(n_630),
.A2(n_575),
.B(n_25),
.C(n_27),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_679),
.Y(n_716)
);

AOI221xp5_ASAP7_75t_L g717 ( 
.A1(n_638),
.A2(n_585),
.B1(n_576),
.B2(n_621),
.C(n_575),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_652),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_658),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_679),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_634),
.B(n_49),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_635),
.A2(n_98),
.B(n_196),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_639),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_105),
.B(n_194),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_669),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_646),
.A2(n_685),
.B(n_687),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_688),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_727)
);

AOI21x1_ASAP7_75t_L g728 ( 
.A1(n_665),
.A2(n_667),
.B(n_636),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_688),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_683),
.B(n_28),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_644),
.Y(n_731)
);

OAI21x1_ASAP7_75t_L g732 ( 
.A1(n_643),
.A2(n_106),
.B(n_191),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_682),
.Y(n_733)
);

OA21x2_ASAP7_75t_L g734 ( 
.A1(n_639),
.A2(n_645),
.B(n_656),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_670),
.B(n_29),
.Y(n_735)
);

AOI21xp33_ASAP7_75t_L g736 ( 
.A1(n_654),
.A2(n_686),
.B(n_684),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_684),
.B(n_30),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_686),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_667),
.A2(n_31),
.B(n_32),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_682),
.B(n_31),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_654),
.B(n_32),
.Y(n_741)
);

INVx5_ASAP7_75t_L g742 ( 
.A(n_670),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_698),
.Y(n_743)
);

OAI211xp5_ASAP7_75t_SL g744 ( 
.A1(n_740),
.A2(n_673),
.B(n_651),
.C(n_666),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_705),
.B(n_675),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_709),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_716),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_698),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_692),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_738),
.A2(n_730),
.B1(n_723),
.B2(n_706),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_SL g752 ( 
.A1(n_739),
.A2(n_673),
.B(n_637),
.C(n_655),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_707),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_729),
.B(n_637),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_738),
.A2(n_640),
.B1(n_657),
.B2(n_633),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_705),
.B(n_649),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_730),
.A2(n_720),
.B1(n_733),
.B2(n_737),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_741),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_714),
.B(n_33),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_729),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_735),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_SL g762 ( 
.A(n_717),
.B(n_727),
.C(n_696),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_SL g763 ( 
.A1(n_701),
.A2(n_640),
.B1(n_657),
.B2(n_633),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_697),
.A2(n_674),
.B1(n_677),
.B2(n_637),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_693),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_735),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_710),
.B(n_702),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_735),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_702),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_735),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_L g771 ( 
.A1(n_710),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_710),
.B(n_36),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_692),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_689),
.B(n_655),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_692),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_736),
.A2(n_674),
.B1(n_655),
.B2(n_677),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_SL g777 ( 
.A(n_695),
.B(n_37),
.C(n_38),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_710),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_702),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_713),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_713),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_692),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_700),
.B(n_669),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_721),
.A2(n_674),
.B1(n_677),
.B2(n_42),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_718),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_SL g786 ( 
.A(n_718),
.B(n_40),
.Y(n_786)
);

OAI221xp5_ASAP7_75t_L g787 ( 
.A1(n_715),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.C(n_669),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_718),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_691),
.B(n_45),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_721),
.A2(n_206),
.B1(n_54),
.B2(n_58),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_718),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_690),
.A2(n_52),
.B(n_61),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_742),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_793)
);

OAI221xp5_ASAP7_75t_L g794 ( 
.A1(n_715),
.A2(n_190),
.B1(n_66),
.B2(n_68),
.C(n_69),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_SL g795 ( 
.A(n_690),
.B(n_65),
.C(n_70),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_703),
.A2(n_184),
.B(n_72),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_703),
.A2(n_179),
.B(n_73),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_709),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_691),
.B(n_71),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_691),
.Y(n_800)
);

CKINVDCx11_ASAP7_75t_R g801 ( 
.A(n_725),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_742),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_709),
.Y(n_803)
);

OAI31xp33_ASAP7_75t_L g804 ( 
.A1(n_766),
.A2(n_712),
.A3(n_725),
.B(n_721),
.Y(n_804)
);

OAI211xp5_ASAP7_75t_SL g805 ( 
.A1(n_777),
.A2(n_731),
.B(n_712),
.C(n_719),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_748),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_745),
.B(n_699),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_784),
.A2(n_694),
.B(n_726),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_777),
.B(n_751),
.C(n_795),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_751),
.A2(n_721),
.B1(n_699),
.B2(n_742),
.Y(n_810)
);

AOI222xp33_ASAP7_75t_L g811 ( 
.A1(n_762),
.A2(n_721),
.B1(n_742),
.B2(n_719),
.C1(n_722),
.C2(n_694),
.Y(n_811)
);

AOI222xp33_ASAP7_75t_L g812 ( 
.A1(n_757),
.A2(n_721),
.B1(n_742),
.B2(n_722),
.C1(n_699),
.C2(n_732),
.Y(n_812)
);

OAI22xp33_ASAP7_75t_L g813 ( 
.A1(n_794),
.A2(n_728),
.B1(n_734),
.B2(n_731),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_757),
.A2(n_787),
.B1(n_771),
.B2(n_758),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_771),
.A2(n_734),
.B1(n_731),
.B2(n_708),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_753),
.Y(n_816)
);

OAI211xp5_ASAP7_75t_L g817 ( 
.A1(n_792),
.A2(n_734),
.B(n_732),
.C(n_726),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_786),
.A2(n_700),
.B1(n_724),
.B2(n_711),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_761),
.B(n_768),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_770),
.B(n_708),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_791),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_785),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_774),
.A2(n_754),
.B1(n_784),
.B2(n_778),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_760),
.B(n_708),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_744),
.A2(n_724),
.B1(n_711),
.B2(n_708),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_748),
.B(n_77),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_776),
.A2(n_78),
.B(n_81),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_755),
.B(n_82),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_781),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_769),
.B(n_779),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_755),
.B(n_87),
.Y(n_831)
);

AOI221xp5_ASAP7_75t_L g832 ( 
.A1(n_752),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.C(n_93),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_743),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_749),
.Y(n_834)
);

AOI221xp5_ASAP7_75t_L g835 ( 
.A1(n_795),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_108),
.Y(n_835)
);

AO21x1_ASAP7_75t_L g836 ( 
.A1(n_793),
.A2(n_109),
.B(n_110),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_759),
.B(n_111),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_773),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_785),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_803),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_776),
.A2(n_112),
.B(n_114),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_790),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_842)
);

AOI211xp5_ASAP7_75t_L g843 ( 
.A1(n_793),
.A2(n_122),
.B(n_124),
.C(n_125),
.Y(n_843)
);

AOI211xp5_ASAP7_75t_L g844 ( 
.A1(n_772),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_765),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_747),
.B(n_133),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_782),
.B(n_134),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_747),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_SL g849 ( 
.A1(n_746),
.A2(n_802),
.B1(n_780),
.B2(n_767),
.Y(n_849)
);

AOI222xp33_ASAP7_75t_L g850 ( 
.A1(n_790),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.C1(n_141),
.C2(n_144),
.Y(n_850)
);

AOI21xp33_ASAP7_75t_L g851 ( 
.A1(n_764),
.A2(n_145),
.B(n_149),
.Y(n_851)
);

NOR2x1_ASAP7_75t_L g852 ( 
.A(n_775),
.B(n_151),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_796),
.A2(n_797),
.B1(n_789),
.B2(n_756),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_806),
.B(n_798),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_807),
.B(n_798),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_848),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_820),
.B(n_807),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_840),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_816),
.B(n_763),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_821),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_808),
.B(n_783),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_820),
.B(n_848),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_824),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_808),
.B(n_819),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_840),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_819),
.B(n_783),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_834),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_820),
.B(n_846),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_833),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_833),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_838),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_846),
.B(n_783),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_822),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_815),
.Y(n_874)
);

OR2x2_ASAP7_75t_SL g875 ( 
.A(n_809),
.B(n_788),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_830),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_812),
.B(n_800),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_839),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_823),
.B(n_785),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_839),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_826),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_814),
.A2(n_789),
.B1(n_767),
.B2(n_750),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_823),
.B(n_785),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_837),
.B(n_775),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_827),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_810),
.B(n_756),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_827),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_810),
.B(n_750),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_825),
.B(n_801),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_827),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_814),
.B(n_746),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_882),
.B(n_843),
.C(n_804),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_858),
.Y(n_894)
);

OAI211xp5_ASAP7_75t_L g895 ( 
.A1(n_874),
.A2(n_850),
.B(n_835),
.C(n_829),
.Y(n_895)
);

OAI31xp33_ASAP7_75t_L g896 ( 
.A1(n_883),
.A2(n_845),
.A3(n_805),
.B(n_831),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_874),
.A2(n_831),
.B1(n_828),
.B2(n_842),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_858),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_858),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_869),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_886),
.A2(n_836),
.B(n_813),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_SL g902 ( 
.A(n_885),
.B(n_853),
.C(n_817),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_882),
.A2(n_828),
.B1(n_832),
.B2(n_851),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_854),
.B(n_825),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_871),
.B(n_881),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_879),
.B(n_844),
.C(n_849),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_865),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_865),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_871),
.B(n_811),
.Y(n_909)
);

OAI211xp5_ASAP7_75t_SL g910 ( 
.A1(n_854),
.A2(n_829),
.B(n_847),
.C(n_852),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_869),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_856),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_SL g913 ( 
.A1(n_886),
.A2(n_841),
.B1(n_799),
.B2(n_158),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_857),
.B(n_841),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_875),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_881),
.B(n_855),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_894),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_914),
.B(n_916),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_904),
.B(n_855),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_914),
.B(n_864),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_907),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_907),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_912),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_908),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_914),
.B(n_864),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_912),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_SL g927 ( 
.A(n_909),
.B(n_883),
.C(n_880),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_900),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_905),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_914),
.B(n_864),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_904),
.B(n_855),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_929),
.B(n_919),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_921),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_923),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_926),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_927),
.A2(n_906),
.B1(n_893),
.B2(n_895),
.Y(n_936)
);

NAND4xp25_ASAP7_75t_L g937 ( 
.A(n_918),
.B(n_893),
.C(n_896),
.D(n_901),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_918),
.B(n_860),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_920),
.B(n_915),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_SL g940 ( 
.A1(n_920),
.A2(n_896),
.B(n_910),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_919),
.B(n_881),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_940),
.B(n_931),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_939),
.B(n_930),
.Y(n_943)
);

INVx3_ASAP7_75t_SL g944 ( 
.A(n_939),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_937),
.B(n_931),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_934),
.A2(n_915),
.B(n_936),
.C(n_935),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_938),
.B(n_902),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_936),
.B(n_921),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_932),
.B(n_924),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_933),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_948),
.B(n_941),
.Y(n_951)
);

AOI21xp33_ASAP7_75t_SL g952 ( 
.A1(n_946),
.A2(n_930),
.B(n_925),
.Y(n_952)
);

AOI321xp33_ASAP7_75t_L g953 ( 
.A1(n_942),
.A2(n_915),
.A3(n_903),
.B1(n_891),
.B2(n_877),
.C(n_890),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_950),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_945),
.B(n_925),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_954),
.Y(n_956)
);

NAND2x1_ASAP7_75t_L g957 ( 
.A(n_951),
.B(n_943),
.Y(n_957)
);

OAI32xp33_ASAP7_75t_L g958 ( 
.A1(n_955),
.A2(n_947),
.A3(n_949),
.B1(n_892),
.B2(n_891),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_SL g959 ( 
.A(n_957),
.B(n_944),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_956),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_958),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_956),
.B(n_952),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_960),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_961),
.B(n_962),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_959),
.B(n_943),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_962),
.Y(n_966)
);

NAND4xp25_ASAP7_75t_L g967 ( 
.A(n_959),
.B(n_953),
.C(n_897),
.D(n_860),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_SL g968 ( 
.A(n_961),
.B(n_913),
.C(n_890),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_959),
.B(n_897),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_960),
.Y(n_970)
);

OAI211xp5_ASAP7_75t_SL g971 ( 
.A1(n_964),
.A2(n_922),
.B(n_924),
.C(n_888),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_966),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_969),
.A2(n_922),
.B(n_886),
.Y(n_973)
);

OAI211xp5_ASAP7_75t_L g974 ( 
.A1(n_965),
.A2(n_860),
.B(n_890),
.C(n_873),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_963),
.Y(n_975)
);

AOI222xp33_ASAP7_75t_L g976 ( 
.A1(n_968),
.A2(n_888),
.B1(n_877),
.B2(n_859),
.C1(n_879),
.C2(n_884),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_967),
.A2(n_888),
.B1(n_877),
.B2(n_892),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_975),
.A2(n_970),
.B1(n_884),
.B2(n_859),
.Y(n_978)
);

AOI211xp5_ASAP7_75t_L g979 ( 
.A1(n_972),
.A2(n_880),
.B(n_884),
.C(n_875),
.Y(n_979)
);

AOI31xp33_ASAP7_75t_L g980 ( 
.A1(n_974),
.A2(n_868),
.A3(n_889),
.B(n_872),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_R g981 ( 
.A(n_973),
.B(n_873),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_976),
.B(n_908),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_977),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_971),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_984),
.B(n_878),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_983),
.B(n_878),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_978),
.B(n_889),
.C(n_856),
.Y(n_987)
);

NAND3xp33_ASAP7_75t_L g988 ( 
.A(n_979),
.B(n_878),
.C(n_861),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_982),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_980),
.Y(n_990)
);

AOI222xp33_ASAP7_75t_L g991 ( 
.A1(n_981),
.A2(n_917),
.B1(n_928),
.B2(n_863),
.C1(n_867),
.C2(n_861),
.Y(n_991)
);

NAND4xp75_ASAP7_75t_L g992 ( 
.A(n_978),
.B(n_868),
.C(n_861),
.D(n_872),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_990),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_989),
.A2(n_917),
.B1(n_928),
.B2(n_863),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_985),
.B(n_917),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_SL g996 ( 
.A(n_986),
.B(n_868),
.C(n_872),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_SL g997 ( 
.A(n_988),
.B(n_867),
.C(n_154),
.Y(n_997)
);

XOR2xp5_ASAP7_75t_L g998 ( 
.A(n_985),
.B(n_887),
.Y(n_998)
);

NAND5xp2_ASAP7_75t_L g999 ( 
.A(n_991),
.B(n_866),
.C(n_876),
.D(n_162),
.E(n_166),
.Y(n_999)
);

BUFx4f_ASAP7_75t_SL g1000 ( 
.A(n_993),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_995),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_992),
.Y(n_1002)
);

AOI211xp5_ASAP7_75t_L g1003 ( 
.A1(n_999),
.A2(n_987),
.B(n_887),
.C(n_857),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_L g1004 ( 
.A(n_994),
.B(n_899),
.C(n_898),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1000),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1001),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1002),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_998),
.Y(n_1008)
);

NOR4xp75_ASAP7_75t_L g1009 ( 
.A(n_1008),
.B(n_996),
.C(n_1004),
.D(n_167),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1007),
.A2(n_899),
.B1(n_898),
.B2(n_894),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_SL g1011 ( 
.A(n_1006),
.B(n_911),
.C(n_900),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1010),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1009),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_L g1014 ( 
.A(n_1013),
.B(n_1005),
.C(n_1011),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_1012),
.A2(n_911),
.B(n_857),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_1013),
.A2(n_857),
.B(n_159),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_1016),
.B(n_857),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_1014),
.A2(n_152),
.B(n_168),
.Y(n_1018)
);

AOI322xp5_ASAP7_75t_L g1019 ( 
.A1(n_1018),
.A2(n_1015),
.A3(n_876),
.B1(n_862),
.B2(n_866),
.C1(n_869),
.C2(n_870),
.Y(n_1019)
);

AOI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1019),
.A2(n_1017),
.B1(n_170),
.B2(n_171),
.C(n_172),
.Y(n_1020)
);

AOI211xp5_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_169),
.B(n_175),
.C(n_176),
.Y(n_1021)
);


endmodule