module fake_netlist_6_751_n_1680 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1680);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1680;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_38),
.Y(n_166)
);

BUFx8_ASAP7_75t_SL g167 ( 
.A(n_39),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_11),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_21),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_28),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_39),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_157),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_21),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_64),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_25),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_53),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_49),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_112),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_33),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_127),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_75),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_45),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_80),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_7),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_17),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_45),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_115),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_31),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_52),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_16),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_50),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_26),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_77),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_44),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_54),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_41),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_17),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_106),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_139),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_88),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_96),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_25),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_38),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_153),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_16),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_62),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_105),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_26),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_148),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_28),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_97),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_6),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_124),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_120),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_63),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_131),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_8),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_92),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_116),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_87),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_82),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_3),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_5),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_154),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_123),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_100),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_51),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_132),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_43),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_60),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_31),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_14),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_98),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_24),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_107),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_36),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_32),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_144),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_119),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_67),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_78),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_61),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_70),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_18),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_94),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_47),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_35),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_113),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_13),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_73),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_20),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_0),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_29),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_83),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_33),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_141),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_150),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_22),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_46),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_27),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_167),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_236),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_174),
.B(n_1),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_221),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_287),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_205),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_4),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_241),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_301),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_234),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_212),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_234),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_214),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_160),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_219),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_169),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_159),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_160),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_173),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_173),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_176),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_176),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_224),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_226),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_169),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_170),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_232),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_226),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_251),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_306),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_251),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_242),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_245),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_247),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_273),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_248),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_252),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_273),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_166),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_185),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_200),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_201),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_257),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_215),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_218),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_263),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_174),
.B(n_10),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_203),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_237),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_170),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_240),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_171),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_246),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_277),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_204),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_261),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_207),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_327),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_386),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_337),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_334),
.B(n_260),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_345),
.B(n_168),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_341),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_346),
.B(n_274),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_343),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_354),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_363),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_364),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_325),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_374),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_274),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_338),
.B(n_260),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_322),
.B(n_220),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_358),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_365),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_367),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_R g430 ( 
.A(n_387),
.B(n_389),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_342),
.B(n_220),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_321),
.B(n_379),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_385),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_369),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_368),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_344),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_316),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_319),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_319),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_318),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_320),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_342),
.B(n_269),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_324),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_324),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_356),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_R g453 ( 
.A(n_332),
.B(n_162),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_361),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_357),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_384),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_388),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_326),
.B(n_269),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_348),
.B(n_269),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_384),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_382),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_369),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_436),
.B(n_271),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_462),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

INVx4_ASAP7_75t_SL g466 ( 
.A(n_426),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_397),
.B(n_441),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_439),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_315),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_419),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_317),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_422),
.B(n_271),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_323),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_330),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_418),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_422),
.B(n_277),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_277),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_418),
.B(n_265),
.Y(n_479)
);

INVx6_ASAP7_75t_L g480 ( 
.A(n_426),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_R g481 ( 
.A(n_456),
.B(n_171),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

OAI22xp33_ASAP7_75t_L g484 ( 
.A1(n_399),
.A2(n_281),
.B1(n_328),
.B2(n_210),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_408),
.B(n_333),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_461),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_432),
.B(n_161),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_426),
.B(n_277),
.Y(n_491)
);

NOR2x1p5_ASAP7_75t_L g492 ( 
.A(n_391),
.B(n_180),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_432),
.B(n_163),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_408),
.B(n_350),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_349),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_452),
.B(n_351),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_460),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_401),
.B(n_164),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_442),
.B(n_285),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_401),
.B(n_165),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_431),
.B(n_348),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_398),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_405),
.B(n_352),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_442),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_432),
.B(n_352),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_399),
.A2(n_177),
.B1(n_187),
.B2(n_184),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_396),
.B(n_353),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_413),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_403),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_432),
.B(n_353),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_400),
.B(n_355),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

BUFx8_ASAP7_75t_SL g525 ( 
.A(n_454),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_393),
.B(n_172),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_430),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_406),
.B(n_355),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_446),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_409),
.A2(n_162),
.B1(n_199),
.B2(n_198),
.Y(n_531)
);

BUFx6f_ASAP7_75t_SL g532 ( 
.A(n_410),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_415),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_411),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_427),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_415),
.A2(n_305),
.B1(n_297),
.B2(n_388),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_417),
.A2(n_268),
.B1(n_182),
.B2(n_186),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_360),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_417),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_407),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_428),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_447),
.B(n_285),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

BUFx8_ASAP7_75t_SL g548 ( 
.A(n_429),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_416),
.B(n_360),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_447),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_393),
.B(n_181),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_423),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_420),
.B(n_366),
.C(n_362),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_420),
.A2(n_390),
.B1(n_377),
.B2(n_282),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_447),
.B(n_192),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_421),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_421),
.B(n_362),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_407),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_424),
.B(n_366),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_424),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_447),
.B(n_197),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_425),
.A2(n_229),
.B1(n_243),
.B2(n_231),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_425),
.A2(n_209),
.B1(n_208),
.B2(n_262),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

OAI22x1_ASAP7_75t_L g567 ( 
.A1(n_440),
.A2(n_266),
.B1(n_313),
.B2(n_312),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_434),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_434),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_393),
.B(n_202),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_435),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_435),
.B(n_206),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_457),
.B(n_216),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_437),
.B(n_390),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_444),
.B(n_329),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_414),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_444),
.B(n_223),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_438),
.B(n_329),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_404),
.B(n_225),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_404),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_438),
.B(n_230),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_404),
.B(n_235),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_443),
.B(n_331),
.Y(n_584)
);

BUFx4f_ASAP7_75t_L g585 ( 
.A(n_414),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_443),
.B(n_331),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_414),
.B(n_238),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_414),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_414),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_414),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_448),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_448),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_450),
.B(n_335),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_450),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_450),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_451),
.B(n_244),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_451),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_451),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_401),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_407),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_426),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_436),
.B(n_250),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_436),
.B(n_177),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_467),
.B(n_340),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_608),
.B(n_254),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_488),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_607),
.A2(n_253),
.B1(n_258),
.B2(n_259),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_608),
.B(n_256),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_593),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_264),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_607),
.A2(n_285),
.B1(n_276),
.B2(n_291),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_509),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_467),
.B(n_527),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_593),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_293),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_465),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_296),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_594),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_468),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_463),
.A2(n_266),
.B1(n_313),
.B2(n_312),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_471),
.B(n_178),
.Y(n_626)
);

AO221x1_ASAP7_75t_L g627 ( 
.A1(n_484),
.A2(n_311),
.B1(n_310),
.B2(n_303),
.C(n_280),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_606),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_471),
.B(n_178),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_488),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_532),
.B(n_180),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_475),
.A2(n_463),
.B1(n_479),
.B2(n_480),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_606),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_469),
.B(n_340),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_529),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_475),
.B(n_179),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_529),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_477),
.B(n_179),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_483),
.B(n_183),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_485),
.B(n_183),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_496),
.B(n_184),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_480),
.A2(n_270),
.B1(n_188),
.B2(n_190),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_474),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_543),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_594),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_557),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_519),
.B(n_187),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_519),
.B(n_190),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_497),
.B(n_194),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_503),
.B(n_194),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_472),
.A2(n_285),
.B1(n_191),
.B2(n_278),
.Y(n_653)
);

NAND2x1_ASAP7_75t_L g654 ( 
.A(n_480),
.B(n_335),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_540),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_571),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_466),
.B(n_285),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_507),
.B(n_195),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_523),
.B(n_195),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_584),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_510),
.B(n_196),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_511),
.B(n_196),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_576),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_466),
.B(n_527),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_584),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_495),
.A2(n_189),
.B1(n_191),
.B2(n_278),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_517),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_521),
.B(n_533),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_466),
.B(n_285),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_535),
.B(n_561),
.Y(n_671)
);

NAND2x1p5_ASAP7_75t_L g672 ( 
.A(n_491),
.B(n_336),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_565),
.B(n_198),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_523),
.B(n_199),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_528),
.B(n_233),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_549),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_528),
.B(n_285),
.Y(n_677)
);

NOR2x1p5_ASAP7_75t_L g678 ( 
.A(n_513),
.B(n_486),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_563),
.A2(n_495),
.B1(n_567),
.B2(n_538),
.C(n_302),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_473),
.B(n_233),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_566),
.B(n_267),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_568),
.B(n_267),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_494),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_569),
.B(n_336),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

BUFx5_ASAP7_75t_L g686 ( 
.A(n_493),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_472),
.B(n_603),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_574),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_574),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_603),
.B(n_275),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_574),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_542),
.B(n_189),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

BUFx8_ASAP7_75t_L g694 ( 
.A(n_532),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_515),
.A2(n_295),
.B1(n_308),
.B2(n_289),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_498),
.B(n_502),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_499),
.B(n_292),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_498),
.B(n_294),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_515),
.B(n_339),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_502),
.B(n_294),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_515),
.A2(n_298),
.B1(n_308),
.B2(n_295),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_499),
.B(n_298),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_476),
.B(n_211),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_518),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_531),
.B(n_280),
.Y(n_705)
);

NOR2x1p5_ASAP7_75t_L g706 ( 
.A(n_537),
.B(n_286),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_494),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_558),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_586),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_515),
.B(n_339),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_522),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_516),
.B(n_213),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_536),
.B(n_93),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_476),
.B(n_604),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_598),
.Y(n_715)
);

OAI221xp5_ASAP7_75t_L g716 ( 
.A1(n_538),
.A2(n_217),
.B1(n_227),
.B2(n_228),
.C(n_249),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_522),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_255),
.C(n_307),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_470),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_520),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_553),
.B(n_573),
.C(n_572),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_522),
.A2(n_280),
.B1(n_302),
.B2(n_300),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_522),
.A2(n_307),
.B1(n_300),
.B2(n_299),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_558),
.A2(n_299),
.B(n_290),
.C(n_288),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_494),
.B(n_290),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_494),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_584),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_481),
.A2(n_288),
.B1(n_286),
.B2(n_239),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_464),
.B(n_239),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_560),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_560),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_478),
.B(n_518),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_505),
.B(n_514),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_520),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_487),
.Y(n_735)
);

NOR2x2_ASAP7_75t_L g736 ( 
.A(n_481),
.B(n_12),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_548),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_478),
.B(n_57),
.Y(n_738)
);

NOR2xp67_ASAP7_75t_L g739 ( 
.A(n_552),
.B(n_65),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_501),
.B(n_482),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_R g741 ( 
.A(n_537),
.B(n_56),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_478),
.B(n_68),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_478),
.B(n_158),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_539),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_744)
);

INVx8_ASAP7_75t_L g745 ( 
.A(n_493),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_489),
.B(n_69),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_478),
.B(n_152),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_530),
.B(n_490),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_602),
.B(n_149),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_530),
.B(n_15),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_602),
.B(n_145),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_602),
.B(n_133),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_505),
.B(n_130),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_545),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_514),
.B(n_128),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_500),
.B(n_126),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_585),
.A2(n_125),
.B(n_121),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_548),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_500),
.B(n_117),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_500),
.B(n_109),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_587),
.A2(n_19),
.B(n_24),
.C(n_27),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_524),
.B(n_103),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_595),
.A2(n_29),
.B(n_32),
.C(n_35),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_490),
.B(n_37),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_589),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_597),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_554),
.B(n_95),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_572),
.B(n_37),
.C(n_40),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_714),
.A2(n_585),
.B(n_491),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_687),
.A2(n_544),
.B(n_547),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_655),
.B(n_588),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_632),
.A2(n_547),
.B(n_544),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_644),
.B(n_530),
.Y(n_774)
);

O2A1O1Ixp5_ASAP7_75t_L g775 ( 
.A1(n_610),
.A2(n_613),
.B(n_677),
.C(n_620),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_708),
.A2(n_573),
.B(n_582),
.C(n_556),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_676),
.B(n_555),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_708),
.A2(n_582),
.B(n_562),
.C(n_556),
.Y(n_778)
);

AOI21x1_ASAP7_75t_L g779 ( 
.A1(n_696),
.A2(n_733),
.B(n_670),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_717),
.B(n_492),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_731),
.A2(n_596),
.B(n_597),
.Y(n_781)
);

BUFx4f_ASAP7_75t_L g782 ( 
.A(n_740),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_731),
.B(n_578),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_626),
.A2(n_555),
.B1(n_504),
.B2(n_508),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_642),
.B(n_512),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_570),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_626),
.B(n_525),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_732),
.A2(n_512),
.B(n_544),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_615),
.A2(n_622),
.B(n_630),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_661),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_629),
.B(n_578),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_624),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_629),
.A2(n_493),
.B1(n_578),
.B2(n_562),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_630),
.A2(n_590),
.B(n_591),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_666),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_616),
.A2(n_599),
.B(n_601),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_609),
.B(n_578),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_704),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_666),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_730),
.B(n_578),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_692),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_669),
.A2(n_590),
.B(n_591),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_649),
.B(n_493),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_649),
.B(n_493),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_671),
.A2(n_534),
.B(n_541),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_614),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_650),
.B(n_605),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_650),
.B(n_605),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_758),
.B(n_539),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_619),
.A2(n_534),
.B(n_541),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_704),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_623),
.A2(n_550),
.B(n_524),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_647),
.A2(n_550),
.B(n_583),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_724),
.A2(n_580),
.B(n_526),
.C(n_551),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_659),
.B(n_605),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_688),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_745),
.A2(n_506),
.B(n_546),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_711),
.B(n_577),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_659),
.B(n_577),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_R g820 ( 
.A(n_737),
.B(n_577),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_644),
.A2(n_599),
.B(n_506),
.C(n_546),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_674),
.B(n_554),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_704),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_720),
.B(n_539),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_734),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_674),
.A2(n_581),
.B1(n_554),
.B2(n_600),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_675),
.B(n_600),
.Y(n_827)
);

AO22x1_ASAP7_75t_L g828 ( 
.A1(n_712),
.A2(n_525),
.B1(n_41),
.B2(n_42),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_745),
.A2(n_670),
.B(n_657),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_689),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_712),
.A2(n_592),
.B1(n_559),
.B2(n_43),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_SL g832 ( 
.A1(n_753),
.A2(n_40),
.B(n_42),
.C(n_46),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_642),
.B(n_592),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_719),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_697),
.A2(n_559),
.B(n_49),
.C(n_51),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_702),
.A2(n_48),
.B(n_72),
.C(n_86),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_729),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_745),
.A2(n_90),
.B(n_91),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_657),
.A2(n_48),
.B(n_665),
.Y(n_839)
);

CKINVDCx10_ASAP7_75t_R g840 ( 
.A(n_694),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_704),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_677),
.A2(n_756),
.B(n_767),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_617),
.B(n_618),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_616),
.A2(n_691),
.B(n_636),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_612),
.A2(n_744),
.B1(n_653),
.B2(n_679),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_L g846 ( 
.A(n_702),
.B(n_705),
.C(n_680),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_665),
.A2(n_611),
.B(n_633),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_612),
.A2(n_744),
.B1(n_653),
.B2(n_664),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_721),
.A2(n_765),
.B(n_766),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_634),
.B(n_680),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_668),
.B(n_685),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_711),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_635),
.B(n_637),
.Y(n_853)
);

OAI321xp33_ASAP7_75t_L g854 ( 
.A1(n_625),
.A2(n_754),
.A3(n_728),
.B1(n_768),
.B2(n_716),
.C(n_718),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_725),
.B(n_645),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_725),
.B(n_646),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_628),
.A2(n_678),
.B1(n_660),
.B2(n_648),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_656),
.B(n_721),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_728),
.B(n_693),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_625),
.A2(n_700),
.B(n_698),
.C(n_761),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_699),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_698),
.A2(n_700),
.B(n_763),
.C(n_703),
.Y(n_862)
);

OAI21xp33_ASAP7_75t_L g863 ( 
.A1(n_709),
.A2(n_715),
.B(n_723),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_683),
.B(n_726),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_759),
.A2(n_760),
.B(n_751),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_749),
.A2(n_752),
.B(n_735),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_707),
.A2(n_746),
.B1(n_713),
.B2(n_739),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_690),
.A2(n_695),
.B1(n_701),
.B2(n_638),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_748),
.B(n_662),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_667),
.B(n_750),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_699),
.B(n_710),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_710),
.B(n_741),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_654),
.A2(n_762),
.B(n_753),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_755),
.A2(n_762),
.B(n_738),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_639),
.B(n_651),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_742),
.A2(n_743),
.B(n_747),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_640),
.A2(n_681),
.B(n_682),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_631),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_SL g879 ( 
.A1(n_764),
.A2(n_673),
.B(n_641),
.C(n_663),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_764),
.A2(n_652),
.B(n_658),
.C(n_672),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_672),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_757),
.A2(n_686),
.B(n_643),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_694),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_686),
.A2(n_627),
.B(n_722),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_684),
.A2(n_686),
.B(n_706),
.C(n_741),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_684),
.Y(n_886)
);

NAND2x1_ASAP7_75t_L g887 ( 
.A(n_684),
.B(n_686),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_686),
.B(n_736),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_686),
.A2(n_731),
.B1(n_629),
.B2(n_626),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_684),
.A2(n_626),
.B1(n_629),
.B2(n_607),
.Y(n_890)
);

INVx11_ASAP7_75t_L g891 ( 
.A(n_694),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_708),
.A2(n_463),
.B(n_613),
.C(n_610),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_758),
.B(n_621),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_737),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_626),
.B(n_629),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_731),
.B(n_608),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_708),
.A2(n_632),
.B(n_731),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_L g900 ( 
.A1(n_626),
.A2(n_629),
.B(n_608),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_655),
.B(n_527),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_661),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_655),
.B(n_527),
.Y(n_905)
);

OAI321xp33_ASAP7_75t_L g906 ( 
.A1(n_626),
.A2(n_629),
.A3(n_744),
.B1(n_625),
.B2(n_608),
.C(n_754),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_608),
.Y(n_908)
);

BUFx12f_ASAP7_75t_L g909 ( 
.A(n_694),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_708),
.A2(n_632),
.B(n_731),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_708),
.A2(n_632),
.B(n_731),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_L g914 ( 
.A(n_626),
.B(n_629),
.C(n_608),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_731),
.B(n_608),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_626),
.A2(n_629),
.B(n_608),
.C(n_613),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_621),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_704),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_731),
.B(n_608),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_729),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_696),
.A2(n_733),
.B(n_670),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_661),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_612),
.A2(n_731),
.B1(n_744),
.B2(n_730),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_708),
.A2(n_632),
.B(n_731),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_731),
.B(n_608),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_708),
.A2(n_463),
.B(n_613),
.C(n_610),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_737),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_612),
.A2(n_731),
.B1(n_744),
.B2(n_730),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_612),
.A2(n_731),
.B1(n_744),
.B2(n_730),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_731),
.B(n_608),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_704),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_644),
.B(n_467),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_642),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_612),
.A2(n_731),
.B1(n_744),
.B2(n_730),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_731),
.B(n_608),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_731),
.A2(n_629),
.B1(n_626),
.B2(n_610),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_708),
.A2(n_463),
.B(n_613),
.C(n_610),
.Y(n_940)
);

O2A1O1Ixp5_ASAP7_75t_L g941 ( 
.A1(n_610),
.A2(n_463),
.B(n_613),
.C(n_677),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_626),
.B(n_629),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_661),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_717),
.B(n_688),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_714),
.A2(n_687),
.B(n_632),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_896),
.B(n_943),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_897),
.B(n_908),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_914),
.A2(n_916),
.B1(n_900),
.B2(n_915),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_941),
.A2(n_939),
.B(n_775),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_894),
.A2(n_947),
.B(n_902),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_773),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_845),
.A2(n_906),
.B(n_936),
.C(n_930),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_899),
.A2(n_907),
.B(n_903),
.Y(n_955)
);

AO31x2_ASAP7_75t_L g956 ( 
.A1(n_889),
.A2(n_845),
.A3(n_932),
.B(n_945),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_895),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_805),
.A2(n_866),
.B(n_788),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_934),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_873),
.A2(n_789),
.B(n_847),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_912),
.A2(n_918),
.B(n_913),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_924),
.A2(n_930),
.B(n_929),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_852),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_850),
.B(n_782),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_855),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_798),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_937),
.A2(n_942),
.B(n_797),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_782),
.B(n_774),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_849),
.A2(n_770),
.B(n_813),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_816),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_801),
.B(n_837),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_874),
.A2(n_882),
.B(n_844),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_810),
.A2(n_812),
.B(n_887),
.Y(n_973)
);

OA21x2_ASAP7_75t_L g974 ( 
.A1(n_898),
.A2(n_911),
.B(n_910),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_876),
.A2(n_794),
.B(n_842),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_920),
.B(n_926),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_830),
.Y(n_977)
);

BUFx10_ASAP7_75t_L g978 ( 
.A(n_859),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_921),
.B(n_870),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_856),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_844),
.A2(n_791),
.B(n_807),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_931),
.B(n_938),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_875),
.B(n_846),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_L g984 ( 
.A(n_924),
.B(n_936),
.C(n_929),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_825),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_869),
.B(n_858),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_893),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_892),
.A2(n_927),
.B(n_940),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_798),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_890),
.A2(n_911),
.B1(n_910),
.B2(n_925),
.Y(n_990)
);

AOI21xp33_ASAP7_75t_L g991 ( 
.A1(n_848),
.A2(n_868),
.B(n_860),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_783),
.A2(n_769),
.B(n_925),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_898),
.A2(n_848),
.B(n_854),
.C(n_862),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_808),
.A2(n_819),
.B(n_815),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_822),
.A2(n_827),
.B(n_804),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_SL g996 ( 
.A1(n_787),
.A2(n_831),
.B(n_878),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_834),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_851),
.B(n_771),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_829),
.A2(n_802),
.B(n_865),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_800),
.A2(n_877),
.B(n_803),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_863),
.A2(n_777),
.B(n_843),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_817),
.A2(n_781),
.B(n_796),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_798),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_871),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_786),
.B(n_853),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_806),
.B(n_795),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_SL g1007 ( 
.A1(n_780),
.A2(n_861),
.B(n_864),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_818),
.A2(n_781),
.B(n_796),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_917),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_790),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_826),
.A2(n_884),
.B(n_785),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_784),
.A2(n_778),
.B(n_776),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_814),
.A2(n_821),
.B(n_839),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_835),
.A2(n_880),
.B(n_836),
.C(n_793),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_879),
.A2(n_867),
.B(n_872),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_888),
.A2(n_857),
.B1(n_946),
.B2(n_780),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_799),
.A2(n_904),
.B1(n_923),
.B2(n_944),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_841),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_841),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_852),
.A2(n_881),
.B1(n_935),
.B2(n_811),
.Y(n_1020)
);

OA21x2_ASAP7_75t_L g1021 ( 
.A1(n_885),
.A2(n_838),
.B(n_833),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_886),
.A2(n_946),
.B(n_933),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_905),
.A2(n_933),
.B(n_811),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_841),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_823),
.A2(n_832),
.B(n_901),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_823),
.B(n_919),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_919),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_909),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_792),
.A2(n_824),
.B(n_828),
.Y(n_1029)
);

O2A1O1Ixp5_ASAP7_75t_L g1030 ( 
.A1(n_824),
.A2(n_809),
.B(n_820),
.C(n_893),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_809),
.A2(n_893),
.B(n_928),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_809),
.A2(n_883),
.B(n_891),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_840),
.A2(n_922),
.B(n_779),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_934),
.B(n_850),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_894),
.A2(n_902),
.B(n_899),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_896),
.A2(n_943),
.B(n_900),
.C(n_914),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_916),
.A2(n_889),
.A3(n_943),
.B(n_896),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_916),
.A2(n_914),
.B(n_896),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_807),
.A2(n_815),
.B(n_808),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_896),
.B(n_943),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_916),
.A2(n_914),
.B(n_896),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_807),
.A2(n_815),
.B(n_808),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_934),
.B(n_850),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_916),
.A2(n_914),
.B(n_896),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_935),
.B(n_852),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_896),
.A2(n_943),
.B(n_900),
.C(n_914),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_893),
.B(n_825),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_780),
.B(n_861),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_896),
.B(n_943),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1055)
);

CKINVDCx10_ASAP7_75t_R g1056 ( 
.A(n_840),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_896),
.B(n_943),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_896),
.B(n_943),
.Y(n_1058)
);

AO31x2_ASAP7_75t_L g1059 ( 
.A1(n_916),
.A2(n_889),
.A3(n_943),
.B(n_896),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_773),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_894),
.A2(n_902),
.B(n_899),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_894),
.A2(n_902),
.B(n_899),
.Y(n_1063)
);

NOR2x1_ASAP7_75t_L g1064 ( 
.A(n_914),
.B(n_740),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_916),
.A2(n_914),
.B(n_896),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_896),
.B(n_943),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_917),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_894),
.A2(n_902),
.B(n_899),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_798),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_SL g1070 ( 
.A1(n_916),
.A2(n_817),
.B(n_896),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_801),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_916),
.A2(n_914),
.B(n_896),
.Y(n_1073)
);

AOI222xp33_ASAP7_75t_L g1074 ( 
.A1(n_845),
.A2(n_906),
.B1(n_612),
.B2(n_896),
.C1(n_943),
.C2(n_900),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_798),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_934),
.B(n_850),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_917),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_773),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_916),
.A2(n_889),
.A3(n_943),
.B(n_896),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_L g1081 ( 
.A(n_900),
.B(n_846),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_896),
.A2(n_943),
.B1(n_914),
.B2(n_916),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_779),
.A2(n_922),
.B(n_772),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_935),
.B(n_852),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_896),
.A2(n_943),
.B(n_900),
.C(n_914),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_807),
.A2(n_815),
.B(n_808),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_934),
.B(n_850),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_807),
.A2(n_815),
.B(n_808),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_895),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1070),
.A2(n_972),
.B(n_1002),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1054),
.A2(n_1066),
.B(n_1058),
.C(n_1057),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1054),
.A2(n_1066),
.B1(n_1041),
.B2(n_954),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1089),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_949),
.B(n_976),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_970),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_963),
.Y(n_1096)
);

OR2x6_ASAP7_75t_SL g1097 ( 
.A(n_1082),
.B(n_983),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_982),
.B(n_986),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1034),
.B(n_1046),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1002),
.A2(n_972),
.B(n_952),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1076),
.B(n_1087),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_954),
.A2(n_1036),
.B1(n_1085),
.B2(n_1049),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1060),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1078),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1071),
.B(n_959),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_959),
.B(n_948),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1051),
.B(n_968),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1036),
.A2(n_1049),
.B(n_1085),
.C(n_1038),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1051),
.B(n_964),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_SL g1110 ( 
.A(n_991),
.B(n_1043),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_993),
.A2(n_948),
.B1(n_984),
.B2(n_1073),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_997),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1010),
.Y(n_1113)
);

CKINVDCx8_ASAP7_75t_R g1114 ( 
.A(n_1056),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1047),
.A2(n_1065),
.B(n_962),
.C(n_993),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_L g1116 ( 
.A(n_1001),
.B(n_1064),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1074),
.B(n_950),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1006),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_L g1119 ( 
.A(n_1067),
.B(n_1077),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_971),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_1050),
.B(n_987),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_R g1122 ( 
.A(n_957),
.B(n_985),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_966),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1004),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1004),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_980),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1050),
.B(n_1007),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_990),
.A2(n_980),
.B1(n_965),
.B2(n_974),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1026),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_955),
.A2(n_1035),
.B(n_1061),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1081),
.B(n_974),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_979),
.A2(n_978),
.B1(n_974),
.B2(n_1012),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_978),
.B(n_1031),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1029),
.A2(n_998),
.B1(n_1005),
.B2(n_1016),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_996),
.A2(n_1014),
.B(n_988),
.C(n_1030),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1050),
.B(n_963),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1024),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1027),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1077),
.B(n_1009),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_1048),
.B(n_1084),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1037),
.B(n_1059),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1032),
.B(n_1030),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1048),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_966),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_966),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1037),
.B(n_1059),
.Y(n_1146)
);

AOI21xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1033),
.A2(n_1020),
.B(n_1025),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1019),
.B(n_1022),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_955),
.A2(n_1063),
.B(n_1068),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1037),
.B(n_1080),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_989),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1037),
.B(n_1059),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1003),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1059),
.B(n_1080),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1015),
.A2(n_1017),
.B1(n_951),
.B2(n_992),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1028),
.A2(n_1017),
.B1(n_1019),
.B2(n_1003),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1080),
.B(n_994),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1019),
.B(n_1075),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_1018),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1069),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1015),
.B(n_1069),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_1069),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1075),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1080),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1014),
.A2(n_1023),
.B1(n_1000),
.B2(n_1021),
.Y(n_1166)
);

BUFx2_ASAP7_75t_SL g1167 ( 
.A(n_1023),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_956),
.B(n_1088),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_981),
.A2(n_1008),
.B1(n_1021),
.B2(n_1013),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1021),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_981),
.B(n_994),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_956),
.B(n_967),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_961),
.A2(n_1035),
.B1(n_1068),
.B2(n_1063),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_961),
.A2(n_1061),
.B1(n_967),
.B2(n_969),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_999),
.A2(n_960),
.B(n_958),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_956),
.B(n_1086),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_L g1177 ( 
.A(n_956),
.B(n_1011),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1039),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_975),
.A2(n_1052),
.B(n_1079),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1083),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1044),
.B(n_1072),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1053),
.A2(n_1055),
.B(n_1062),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_L g1184 ( 
.A(n_1040),
.B(n_1045),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_995),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_973),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1070),
.A2(n_1002),
.B(n_972),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1051),
.B(n_968),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1054),
.A2(n_1066),
.B1(n_896),
.B2(n_943),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_983),
.B(n_1034),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1019),
.B(n_935),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1051),
.B(n_968),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1054),
.B(n_1066),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_953),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_993),
.A2(n_916),
.B(n_896),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1070),
.A2(n_1002),
.B(n_972),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_953),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1054),
.B(n_1066),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_977),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1051),
.B(n_968),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1082),
.A2(n_896),
.B(n_943),
.C(n_916),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_985),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1054),
.B(n_1066),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1051),
.B(n_968),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_1082),
.A2(n_896),
.B(n_943),
.C(n_916),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_953),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_993),
.A2(n_943),
.B(n_896),
.Y(n_1207)
);

BUFx8_ASAP7_75t_SL g1208 ( 
.A(n_1028),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1054),
.B(n_782),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_963),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1054),
.A2(n_1066),
.B1(n_1057),
.B2(n_1058),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1054),
.A2(n_1066),
.B1(n_1057),
.B2(n_1058),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_953),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1054),
.B(n_1066),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1034),
.B(n_1046),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_985),
.Y(n_1216)
);

AOI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1074),
.A2(n_943),
.B(n_896),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1070),
.A2(n_972),
.B(n_1002),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1034),
.B(n_1046),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1095),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1127),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1092),
.B(n_1097),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1104),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1120),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1189),
.A2(n_1211),
.B1(n_1212),
.B2(n_1092),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1161),
.B(n_1179),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1211),
.B(n_1212),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1113),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1193),
.A2(n_1203),
.B1(n_1214),
.B2(n_1198),
.Y(n_1229)
);

OAI222xp33_ASAP7_75t_L g1230 ( 
.A1(n_1117),
.A2(n_1102),
.B1(n_1111),
.B2(n_1214),
.C1(n_1203),
.C2(n_1198),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1207),
.A2(n_1110),
.B1(n_1117),
.B2(n_1102),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1103),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1217),
.A2(n_1207),
.B1(n_1111),
.B2(n_1110),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1194),
.Y(n_1234)
);

BUFx8_ASAP7_75t_SL g1235 ( 
.A(n_1208),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1197),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1175),
.A2(n_1180),
.B(n_1090),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1158),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1184),
.A2(n_1183),
.B(n_1171),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1158),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1141),
.B(n_1150),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1182),
.A2(n_1173),
.B(n_1187),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1217),
.A2(n_1142),
.B1(n_1209),
.B2(n_1193),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_1135),
.A2(n_1131),
.B(n_1128),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1206),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1196),
.A2(n_1218),
.B(n_1173),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1213),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1127),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1091),
.B(n_1098),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1182),
.A2(n_1218),
.B(n_1174),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1199),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1134),
.A2(n_1116),
.B1(n_1133),
.B2(n_1132),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1156),
.A2(n_1098),
.B1(n_1094),
.B2(n_1190),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1094),
.A2(n_1195),
.B1(n_1115),
.B2(n_1120),
.Y(n_1254)
);

NAND2x1p5_ASAP7_75t_L g1255 ( 
.A(n_1148),
.B(n_1181),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1114),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1105),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1140),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1099),
.A2(n_1219),
.B1(n_1215),
.B2(n_1128),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1139),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1185),
.A2(n_1101),
.B1(n_1165),
.B2(n_1106),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1121),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1146),
.A2(n_1121),
.B1(n_1109),
.B2(n_1200),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1201),
.A2(n_1205),
.B(n_1108),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1122),
.A2(n_1192),
.B1(n_1204),
.B2(n_1188),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_SL g1266 ( 
.A(n_1202),
.Y(n_1266)
);

INVx4_ASAP7_75t_SL g1267 ( 
.A(n_1140),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1216),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1126),
.A2(n_1125),
.B1(n_1124),
.B2(n_1121),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1112),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1100),
.A2(n_1172),
.B(n_1176),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1119),
.Y(n_1272)
);

INVx11_ASAP7_75t_L g1273 ( 
.A(n_1159),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1162),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1172),
.A2(n_1176),
.B(n_1157),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1093),
.Y(n_1276)
);

INVx4_ASAP7_75t_SL g1277 ( 
.A(n_1140),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1107),
.A2(n_1188),
.B1(n_1204),
.B2(n_1192),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1129),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1138),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1107),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1118),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1200),
.A2(n_1136),
.B1(n_1126),
.B2(n_1148),
.Y(n_1283)
);

CKINVDCx16_ASAP7_75t_R g1284 ( 
.A(n_1136),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1137),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1155),
.A2(n_1131),
.B1(n_1152),
.B2(n_1150),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1167),
.A2(n_1096),
.B1(n_1143),
.B2(n_1210),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1096),
.A2(n_1143),
.B1(n_1210),
.B2(n_1157),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1141),
.A2(n_1154),
.B1(n_1152),
.B2(n_1168),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1151),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1164),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1160),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1181),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1154),
.B(n_1153),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1177),
.A2(n_1123),
.B1(n_1144),
.B2(n_1153),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1163),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1169),
.A2(n_1145),
.B1(n_1186),
.B2(n_1123),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1123),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1147),
.B(n_1144),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1191),
.A2(n_943),
.B(n_896),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1130),
.A2(n_1149),
.B(n_952),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1095),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1092),
.B(n_1038),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1207),
.A2(n_943),
.B(n_896),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1161),
.B(n_1178),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1114),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1162),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1093),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1183),
.A2(n_1180),
.B(n_975),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1217),
.A2(n_943),
.B1(n_896),
.B2(n_1054),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1162),
.Y(n_1312)
);

AOI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1180),
.A2(n_1184),
.B(n_1183),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1180),
.A2(n_1184),
.B(n_1183),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1105),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1217),
.A2(n_943),
.B1(n_896),
.B2(n_1054),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1095),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1095),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1141),
.B(n_1150),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1224),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1227),
.B(n_1229),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1279),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1221),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1246),
.A2(n_1264),
.B(n_1244),
.Y(n_1324)
);

CKINVDCx11_ASAP7_75t_R g1325 ( 
.A(n_1307),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_SL g1326 ( 
.A(n_1307),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1246),
.A2(n_1310),
.B(n_1313),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1275),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1294),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1241),
.B(n_1319),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1294),
.B(n_1304),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1241),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1300),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1258),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1225),
.B(n_1304),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1315),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1289),
.B(n_1286),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1271),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1311),
.A2(n_1316),
.B1(n_1231),
.B2(n_1233),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1222),
.B(n_1243),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1222),
.B(n_1254),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1259),
.B(n_1305),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1257),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1292),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1291),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1242),
.A2(n_1250),
.B(n_1305),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1244),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1302),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1261),
.B(n_1249),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1296),
.B(n_1221),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1282),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1267),
.B(n_1277),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1255),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1252),
.B(n_1269),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1302),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1296),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1296),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1314),
.A2(n_1239),
.B(n_1306),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1237),
.A2(n_1301),
.B(n_1230),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1258),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1248),
.Y(n_1361)
);

OR2x2_ASAP7_75t_SL g1362 ( 
.A(n_1284),
.B(n_1228),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1232),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1295),
.A2(n_1226),
.B(n_1287),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1293),
.A2(n_1245),
.B(n_1247),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1234),
.A2(n_1236),
.B(n_1280),
.Y(n_1366)
);

AO21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1298),
.A2(n_1283),
.B(n_1263),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1262),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1288),
.A2(n_1253),
.B(n_1299),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1270),
.Y(n_1370)
);

AO21x1_ASAP7_75t_L g1371 ( 
.A1(n_1220),
.A2(n_1318),
.B(n_1317),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1309),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1223),
.B(n_1303),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1330),
.B(n_1251),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1358),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1331),
.B(n_1267),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1331),
.B(n_1277),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1365),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1332),
.B(n_1260),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1330),
.B(n_1312),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1324),
.B(n_1277),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1324),
.B(n_1277),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1365),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1332),
.B(n_1285),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1343),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1324),
.B(n_1297),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1328),
.B(n_1274),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1348),
.B(n_1312),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1329),
.B(n_1238),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1344),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1329),
.B(n_1238),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1335),
.B(n_1272),
.Y(n_1392)
);

OAI31xp33_ASAP7_75t_L g1393 ( 
.A1(n_1339),
.A2(n_1281),
.A3(n_1308),
.B(n_1268),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1355),
.B(n_1240),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1321),
.B(n_1240),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_1308),
.Y(n_1396)
);

BUFx2_ASAP7_75t_SL g1397 ( 
.A(n_1352),
.Y(n_1397)
);

BUFx4f_ASAP7_75t_SL g1398 ( 
.A(n_1343),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1341),
.B(n_1290),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1400)
);

OAI21xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1393),
.A2(n_1369),
.B(n_1337),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1392),
.A2(n_1265),
.B1(n_1354),
.B2(n_1349),
.C(n_1369),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1387),
.B(n_1354),
.C(n_1336),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1396),
.B(n_1356),
.Y(n_1404)
);

AND2x2_ASAP7_75t_SL g1405 ( 
.A(n_1381),
.B(n_1352),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1385),
.B(n_1320),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1399),
.A2(n_1337),
.B(n_1349),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1385),
.B(n_1320),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1380),
.B(n_1322),
.Y(n_1409)
);

OAI22x1_ASAP7_75t_SL g1410 ( 
.A1(n_1398),
.A2(n_1256),
.B1(n_1372),
.B2(n_1290),
.Y(n_1410)
);

NAND4xp25_ASAP7_75t_L g1411 ( 
.A(n_1379),
.B(n_1340),
.C(n_1342),
.D(n_1322),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1380),
.B(n_1345),
.Y(n_1412)
);

NAND4xp25_ASAP7_75t_SL g1413 ( 
.A(n_1379),
.B(n_1364),
.C(n_1341),
.D(n_1340),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1394),
.B(n_1357),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1390),
.B(n_1368),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1376),
.A2(n_1364),
.B(n_1360),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1394),
.B(n_1333),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1398),
.B(n_1235),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1394),
.B(n_1388),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1388),
.B(n_1333),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1389),
.B(n_1333),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1387),
.B(n_1347),
.C(n_1366),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1387),
.B(n_1347),
.C(n_1366),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1399),
.A2(n_1362),
.B1(n_1350),
.B2(n_1278),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1389),
.B(n_1333),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1390),
.B(n_1361),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1395),
.B(n_1361),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1395),
.B(n_1351),
.Y(n_1428)
);

NAND3xp33_ASAP7_75t_SL g1429 ( 
.A(n_1374),
.B(n_1371),
.C(n_1256),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1383),
.A2(n_1327),
.B(n_1358),
.Y(n_1430)
);

NAND4xp25_ASAP7_75t_L g1431 ( 
.A(n_1384),
.B(n_1373),
.C(n_1370),
.D(n_1363),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1376),
.A2(n_1362),
.B1(n_1350),
.B2(n_1352),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1381),
.A2(n_1360),
.B(n_1353),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1391),
.B(n_1346),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1391),
.B(n_1346),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1391),
.B(n_1346),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1384),
.B(n_1370),
.C(n_1373),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1386),
.B(n_1346),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1386),
.B(n_1359),
.Y(n_1439)
);

AND2x2_ASAP7_75t_SL g1440 ( 
.A(n_1405),
.B(n_1381),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1438),
.B(n_1382),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1434),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1405),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1435),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1435),
.B(n_1382),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1436),
.B(n_1439),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1436),
.B(n_1382),
.Y(n_1447)
);

AND2x4_ASAP7_75t_SL g1448 ( 
.A(n_1421),
.B(n_1376),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1437),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1422),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1430),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1437),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1419),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1433),
.B(n_1397),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1422),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1423),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1430),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1405),
.B(n_1417),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1421),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1423),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1410),
.B(n_1326),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1414),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1414),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1415),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1426),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1409),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1431),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1427),
.B(n_1378),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1428),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1458),
.B(n_1425),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1455),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1458),
.B(n_1425),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1443),
.B(n_1420),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1455),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1464),
.B(n_1407),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1458),
.B(n_1433),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1450),
.A2(n_1400),
.B(n_1407),
.C(n_1401),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1462),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1454),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1440),
.B(n_1404),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1457),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1448),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1406),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1461),
.B(n_1418),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1457),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1464),
.B(n_1408),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1440),
.B(n_1404),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1462),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1466),
.B(n_1410),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1450),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1443),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1456),
.B(n_1411),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1463),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1460),
.B(n_1411),
.Y(n_1496)
);

AND2x4_ASAP7_75t_SL g1497 ( 
.A(n_1454),
.B(n_1377),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1463),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1449),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1457),
.Y(n_1501)
);

NAND2x2_ASAP7_75t_L g1502 ( 
.A(n_1459),
.B(n_1323),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1440),
.B(n_1375),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1449),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1453),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1451),
.Y(n_1506)
);

OAI21xp33_ASAP7_75t_L g1507 ( 
.A1(n_1491),
.A2(n_1460),
.B(n_1413),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1472),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1484),
.B(n_1468),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1477),
.B(n_1454),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1472),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1475),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1475),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1506),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1479),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1484),
.B(n_1468),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1492),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1506),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1506),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1479),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1489),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1493),
.B(n_1452),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1489),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1476),
.B(n_1452),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1493),
.B(n_1465),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1495),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1477),
.B(n_1454),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1481),
.B(n_1454),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1482),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1465),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1466),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1495),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1470),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_1488),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1502),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1480),
.A2(n_1401),
.B1(n_1416),
.B2(n_1402),
.Y(n_1537)
);

NAND2x1p5_ASAP7_75t_L g1538 ( 
.A(n_1492),
.B(n_1334),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1498),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1498),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1480),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1494),
.B(n_1470),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1480),
.B(n_1448),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1488),
.B(n_1441),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

INVxp67_ASAP7_75t_SL g1547 ( 
.A(n_1499),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1480),
.A2(n_1416),
.B1(n_1432),
.B2(n_1429),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1469),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1524),
.Y(n_1550)
);

CKINVDCx16_ASAP7_75t_R g1551 ( 
.A(n_1515),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1530),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1526),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1544),
.B(n_1497),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1524),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1544),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1523),
.B(n_1500),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1544),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1561)
);

CKINVDCx16_ASAP7_75t_R g1562 ( 
.A(n_1515),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1525),
.B(n_1504),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1542),
.Y(n_1564)
);

NAND2x1_ASAP7_75t_L g1565 ( 
.A(n_1515),
.B(n_1483),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1545),
.B(n_1503),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1518),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1545),
.B(n_1529),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.B(n_1504),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1515),
.B(n_1510),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_1537),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1507),
.A2(n_1497),
.B1(n_1474),
.B2(n_1483),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1532),
.A2(n_1474),
.B1(n_1502),
.B2(n_1424),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1532),
.A2(n_1474),
.B1(n_1502),
.B2(n_1485),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1516),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1547),
.A2(n_1487),
.B(n_1473),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1510),
.B(n_1471),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1528),
.B(n_1471),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1521),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1522),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1528),
.B(n_1473),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1542),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1509),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1517),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1571),
.A2(n_1531),
.B(n_1534),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1571),
.A2(n_1543),
.B(n_1511),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1567),
.B(n_1508),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1567),
.B(n_1325),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1550),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1536),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1564),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1550),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1564),
.Y(n_1594)
);

AND2x2_ASAP7_75t_SL g1595 ( 
.A(n_1551),
.B(n_1548),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1584),
.A2(n_1512),
.B(n_1513),
.C(n_1536),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1584),
.B(n_1549),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1585),
.A2(n_1538),
.B(n_1549),
.C(n_1514),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1557),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_SL g1601 ( 
.A(n_1565),
.B(n_1266),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1558),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1585),
.B(n_1527),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1558),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1560),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1572),
.A2(n_1538),
.B(n_1533),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1551),
.A2(n_1359),
.B1(n_1367),
.B2(n_1541),
.Y(n_1608)
);

AOI322xp5_ASAP7_75t_L g1609 ( 
.A1(n_1562),
.A2(n_1444),
.A3(n_1442),
.B1(n_1446),
.B2(n_1441),
.C1(n_1445),
.C2(n_1447),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1562),
.B(n_1235),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1610),
.B(n_1568),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1610),
.B(n_1560),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1587),
.A2(n_1576),
.B1(n_1565),
.B2(n_1574),
.C(n_1555),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1602),
.B(n_1568),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1589),
.B(n_1555),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1593),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1597),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1600),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1604),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1606),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1605),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1586),
.B(n_1596),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1588),
.B(n_1569),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_L g1626 ( 
.A(n_1601),
.B(n_1570),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1591),
.B(n_1570),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1595),
.A2(n_1570),
.B1(n_1556),
.B2(n_1569),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1563),
.Y(n_1629)
);

OAI21xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1624),
.A2(n_1595),
.B(n_1609),
.Y(n_1630)
);

AOI222xp33_ASAP7_75t_L g1631 ( 
.A1(n_1614),
.A2(n_1576),
.B1(n_1607),
.B2(n_1603),
.C1(n_1608),
.C2(n_1563),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1621),
.A2(n_1601),
.B1(n_1569),
.B2(n_1556),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_SL g1633 ( 
.A(n_1616),
.B(n_1599),
.C(n_1580),
.Y(n_1633)
);

AOI21xp33_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1583),
.B(n_1564),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1612),
.B(n_1594),
.C(n_1592),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1623),
.A2(n_1608),
.B1(n_1583),
.B2(n_1592),
.C(n_1594),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1620),
.A2(n_1573),
.B1(n_1554),
.B2(n_1552),
.C(n_1580),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1625),
.A2(n_1581),
.B1(n_1575),
.B2(n_1559),
.C(n_1552),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1626),
.A2(n_1559),
.B(n_1581),
.Y(n_1639)
);

OAI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1628),
.A2(n_1554),
.B(n_1552),
.Y(n_1640)
);

XOR2xp5_ASAP7_75t_L g1641 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1634),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1639),
.B(n_1615),
.Y(n_1643)
);

AOI211xp5_ASAP7_75t_L g1644 ( 
.A1(n_1630),
.A2(n_1626),
.B(n_1611),
.C(n_1627),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1635),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1640),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1637),
.B(n_1622),
.Y(n_1648)
);

AOI22x1_ASAP7_75t_SL g1649 ( 
.A1(n_1631),
.A2(n_1613),
.B1(n_1619),
.B2(n_1618),
.Y(n_1649)
);

OAI211xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1644),
.A2(n_1636),
.B(n_1638),
.C(n_1617),
.Y(n_1650)
);

NAND4xp25_ASAP7_75t_L g1651 ( 
.A(n_1647),
.B(n_1629),
.C(n_1556),
.D(n_1554),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1645),
.A2(n_1648),
.B1(n_1642),
.B2(n_1646),
.C(n_1641),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1649),
.B(n_1578),
.C(n_1553),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1579),
.C(n_1577),
.Y(n_1654)
);

AOI31xp33_ASAP7_75t_L g1655 ( 
.A1(n_1652),
.A2(n_1538),
.A3(n_1556),
.B(n_1579),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_L g1656 ( 
.A(n_1653),
.B(n_1561),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1650),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1654),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1654),
.B(n_1577),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1654),
.B(n_1582),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1657),
.B(n_1578),
.C(n_1553),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_R g1662 ( 
.A(n_1658),
.B(n_1309),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1578),
.C(n_1553),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1656),
.B(n_1582),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1659),
.B(n_1660),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1664),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1665),
.Y(n_1667)
);

NOR2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1662),
.B(n_1661),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1666),
.A2(n_1663),
.B1(n_1561),
.B2(n_1514),
.Y(n_1669)
);

NAND4xp25_ASAP7_75t_L g1670 ( 
.A(n_1669),
.B(n_1667),
.C(n_1668),
.D(n_1561),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1668),
.B1(n_1561),
.B2(n_1566),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1670),
.A2(n_1566),
.B1(n_1519),
.B2(n_1520),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1671),
.A2(n_1566),
.B1(n_1520),
.B2(n_1519),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1672),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1673),
.B(n_1540),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1674),
.A2(n_1266),
.B1(n_1546),
.B2(n_1539),
.C(n_1482),
.Y(n_1676)
);

XNOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1675),
.B(n_1276),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1676),
.B1(n_1276),
.B2(n_1266),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1501),
.B1(n_1486),
.B2(n_1482),
.C(n_1474),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1276),
.B(n_1273),
.C(n_1486),
.Y(n_1680)
);


endmodule