module fake_jpeg_18472_n_50 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_16),
.B1(n_19),
.B2(n_15),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_9),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_20),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_33),
.B(n_32),
.Y(n_39)
);

AND2x4_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_26),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_25),
.C(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_37),
.B(n_39),
.Y(n_42)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B(n_38),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_2),
.B(n_3),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_3),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_4),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_6),
.C(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_4),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_5),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_5),
.Y(n_50)
);


endmodule