module fake_jpeg_12582_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_55),
.B(n_56),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_1),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_63),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_2),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_104),
.Y(n_140)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_84),
.Y(n_154)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_87),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_20),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_47),
.B1(n_20),
.B2(n_32),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_107),
.A2(n_142),
.B1(n_143),
.B2(n_154),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_25),
.B1(n_50),
.B2(n_28),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_118),
.A2(n_148),
.B1(n_153),
.B2(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_127),
.B(n_136),
.Y(n_181)
);

AND2x4_ASAP7_75t_SL g130 ( 
.A(n_84),
.B(n_49),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_90),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_42),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_70),
.B(n_42),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_144),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_49),
.B1(n_38),
.B2(n_47),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_79),
.A2(n_49),
.B1(n_38),
.B2(n_47),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_40),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_88),
.A2(n_32),
.B1(n_39),
.B2(n_50),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_40),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_38),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_91),
.A2(n_45),
.B1(n_39),
.B2(n_32),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_94),
.A2(n_105),
.B1(n_104),
.B2(n_100),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_58),
.A2(n_45),
.B1(n_38),
.B2(n_49),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_35),
.B1(n_87),
.B2(n_73),
.Y(n_212)
);

HAxp5_ASAP7_75t_SL g166 ( 
.A(n_75),
.B(n_49),
.CON(n_166),
.SN(n_166)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_38),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_65),
.B(n_52),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_99),
.Y(n_179)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_171),
.Y(n_231)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_27),
.B1(n_52),
.B2(n_51),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_120),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_178),
.A2(n_149),
.B(n_128),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_3),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_197),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_117),
.A2(n_27),
.B1(n_51),
.B2(n_36),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_107),
.A2(n_77),
.B1(n_60),
.B2(n_74),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_185),
.A2(n_188),
.B1(n_191),
.B2(n_223),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_186),
.B(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_187),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_143),
.B1(n_125),
.B2(n_63),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_99),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_193),
.B(n_195),
.Y(n_276)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_83),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_49),
.C(n_38),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_215),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_140),
.B(n_137),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_202),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_108),
.B(n_103),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_203),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_117),
.A2(n_36),
.B1(n_66),
.B2(n_62),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_222),
.B1(n_226),
.B2(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_113),
.B(n_2),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_229),
.B1(n_152),
.B2(n_116),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_145),
.A2(n_96),
.B(n_35),
.C(n_83),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_72),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_131),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_138),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_225),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_126),
.A2(n_59),
.B1(n_96),
.B2(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_218),
.Y(n_258)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_128),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_227),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_110),
.A2(n_155),
.B1(n_115),
.B2(n_146),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_109),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_230),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_248),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_180),
.A2(n_152),
.B1(n_156),
.B2(n_129),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_269),
.B1(n_223),
.B2(n_206),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_253),
.A2(n_170),
.B(n_192),
.Y(n_311)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_215),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_264),
.Y(n_309)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

INVx11_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_215),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_188),
.A2(n_116),
.B1(n_109),
.B2(n_122),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_279),
.B1(n_200),
.B2(n_212),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_149),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_268),
.B(n_280),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_200),
.A2(n_160),
.B1(n_5),
.B2(n_6),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_205),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_224),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_180),
.A2(n_160),
.B1(n_5),
.B2(n_6),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_173),
.B(n_196),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_283),
.B(n_10),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_173),
.C(n_190),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_284),
.B(n_257),
.C(n_254),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_293),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_286),
.A2(n_307),
.B1(n_308),
.B2(n_326),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_235),
.B(n_171),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_289),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_196),
.B1(n_227),
.B2(n_220),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_264),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_213),
.B1(n_171),
.B2(n_199),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_292),
.A2(n_303),
.B1(n_236),
.B2(n_252),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_258),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_234),
.A2(n_201),
.B(n_210),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_296),
.A2(n_260),
.B(n_281),
.Y(n_357)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_232),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_314),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_211),
.C(n_197),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_300),
.C(n_304),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_172),
.C(n_230),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_182),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_306),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_271),
.A2(n_235),
.B1(n_239),
.B2(n_248),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_231),
.B(n_198),
.C(n_208),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_261),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_175),
.B1(n_225),
.B2(n_226),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_244),
.A2(n_194),
.B1(n_219),
.B2(n_227),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_313),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_309),
.B(n_305),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_231),
.B(n_216),
.C(n_222),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_317),
.C(n_331),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_214),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_237),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_189),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_318),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_265),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_319),
.A2(n_322),
.B1(n_277),
.B2(n_273),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_253),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_249),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_326)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_327),
.A2(n_328),
.B(n_11),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_17),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_10),
.C(n_11),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_287),
.A2(n_271),
.B(n_245),
.C(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

AOI32xp33_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_301),
.A3(n_313),
.B1(n_293),
.B2(n_306),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_339),
.A2(n_349),
.B(n_351),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_245),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_348),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_346),
.A2(n_354),
.B1(n_368),
.B2(n_316),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_242),
.B(n_273),
.Y(n_349)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_286),
.A2(n_236),
.B1(n_238),
.B2(n_262),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_289),
.A2(n_238),
.B(n_275),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

OAI32xp33_ASAP7_75t_L g356 ( 
.A1(n_288),
.A2(n_256),
.A3(n_263),
.B1(n_240),
.B2(n_272),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_257),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_364),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_288),
.A2(n_281),
.B1(n_255),
.B2(n_256),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_361),
.A2(n_315),
.B1(n_329),
.B2(n_318),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_305),
.A2(n_240),
.B(n_272),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_363),
.B(n_361),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_302),
.A2(n_300),
.B1(n_307),
.B2(n_308),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_295),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_371),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_289),
.A2(n_243),
.B1(n_256),
.B2(n_263),
.Y(n_372)
);

XNOR2x2_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_304),
.Y(n_382)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_374),
.A2(n_395),
.B(n_402),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_368),
.A2(n_317),
.B1(n_322),
.B2(n_312),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_377),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_387),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_382),
.A2(n_407),
.B(n_337),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_351),
.A2(n_326),
.B1(n_328),
.B2(n_284),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_383),
.A2(n_386),
.B1(n_397),
.B2(n_399),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_355),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_343),
.A2(n_342),
.B1(n_369),
.B2(n_357),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_352),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_315),
.B1(n_320),
.B2(n_325),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_347),
.A2(n_346),
.B1(n_354),
.B2(n_349),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_346),
.A2(n_330),
.B1(n_294),
.B2(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_332),
.A2(n_323),
.B1(n_324),
.B2(n_331),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_394),
.A2(n_406),
.B1(n_372),
.B2(n_360),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_343),
.A2(n_243),
.B1(n_295),
.B2(n_282),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_348),
.A2(n_282),
.B1(n_254),
.B2(n_260),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_260),
.B1(n_12),
.B2(n_13),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_400),
.A2(n_336),
.B1(n_337),
.B2(n_365),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_338),
.B(n_11),
.Y(n_401)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_401),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_SL g402 ( 
.A1(n_339),
.A2(n_12),
.B(n_13),
.Y(n_402)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_366),
.A2(n_12),
.A3(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_405),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_17),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_14),
.B1(n_15),
.B2(n_360),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_409),
.A2(n_379),
.B(n_375),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_333),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_420),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_333),
.C(n_345),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_425),
.C(n_428),
.Y(n_446)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_413),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_397),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_416),
.B(n_417),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_359),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_350),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_418),
.B(n_427),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_419),
.A2(n_399),
.B1(n_380),
.B2(n_400),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_364),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_404),
.B(n_367),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_423),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_356),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_396),
.A2(n_363),
.B(n_336),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_407),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_382),
.B(n_384),
.C(n_379),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_401),
.B(n_362),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_340),
.C(n_344),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_389),
.B1(n_393),
.B2(n_388),
.Y(n_450)
);

MAJx2_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_396),
.C(n_383),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_373),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_435),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_375),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_406),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_438),
.A2(n_436),
.B(n_422),
.Y(n_481)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_440),
.B(n_430),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_411),
.A2(n_391),
.B1(n_374),
.B2(n_395),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_443),
.A2(n_450),
.B1(n_437),
.B2(n_419),
.Y(n_469)
);

MAJx2_ASAP7_75t_L g482 ( 
.A(n_444),
.B(n_463),
.C(n_433),
.Y(n_482)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_390),
.C(n_394),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_452),
.C(n_423),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_449),
.A2(n_454),
.B1(n_429),
.B2(n_411),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_420),
.C(n_425),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_414),
.A2(n_385),
.B1(n_381),
.B2(n_358),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_426),
.Y(n_455)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_455),
.Y(n_477)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_459),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_405),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_408),
.Y(n_467)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_428),
.B(n_398),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_468),
.Y(n_491)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_414),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_469),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_421),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_475),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_424),
.B1(n_435),
.B2(n_422),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_473),
.Y(n_494)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_417),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_436),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_481),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_483),
.C(n_484),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_433),
.C(n_434),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_441),
.B(n_365),
.C(n_358),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_483),
.B(n_457),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_489),
.Y(n_512)
);

NOR2x1_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_459),
.Y(n_486)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_486),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_484),
.B(n_438),
.C(n_440),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_SL g490 ( 
.A(n_478),
.B(n_463),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_498),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_476),
.A2(n_438),
.B1(n_444),
.B2(n_456),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_496),
.A2(n_449),
.B1(n_479),
.B2(n_453),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_454),
.C(n_456),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_445),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_442),
.C(n_458),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_500),
.B(n_462),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_482),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_505),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_497),
.A2(n_473),
.B(n_469),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_508),
.B(n_501),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_471),
.C(n_451),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_509),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_506),
.B(n_507),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_335),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_494),
.A2(n_480),
.B(n_451),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_335),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_461),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_511),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_505),
.A2(n_493),
.B1(n_492),
.B2(n_497),
.Y(n_515)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

AOI21x1_ASAP7_75t_SL g524 ( 
.A1(n_517),
.A2(n_503),
.B(n_514),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_488),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_486),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_498),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_513),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_524),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_SL g525 ( 
.A1(n_517),
.A2(n_496),
.B(n_502),
.C(n_508),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_520),
.C(n_521),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_528),
.B(n_516),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_529),
.B(n_530),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_531),
.A2(n_527),
.B(n_526),
.C(n_521),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_532),
.A2(n_520),
.B(n_518),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_534),
.A2(n_533),
.B1(n_464),
.B2(n_472),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_477),
.B(n_515),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_403),
.B(n_495),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_495),
.Y(n_538)
);


endmodule