module fake_jpeg_24757_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_24),
.B1(n_35),
.B2(n_17),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_61),
.B(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_28),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_24),
.B1(n_35),
.B2(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_30),
.Y(n_97)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_24),
.B1(n_23),
.B2(n_34),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_34),
.B1(n_47),
.B2(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_23),
.B1(n_34),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_77),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_48),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_48),
.C(n_42),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_83),
.B1(n_102),
.B2(n_110),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_23),
.B1(n_20),
.B2(n_29),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_87),
.B1(n_105),
.B2(n_45),
.Y(n_116)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_84),
.B(n_94),
.Y(n_132)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_29),
.B1(n_36),
.B2(n_48),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_93),
.B(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_44),
.B1(n_48),
.B2(n_42),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_48),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_38),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_33),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_32),
.B1(n_18),
.B2(n_27),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_38),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_41),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_128),
.B1(n_141),
.B2(n_101),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_55),
.B1(n_25),
.B2(n_27),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_98),
.B1(n_94),
.B2(n_84),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_125),
.C(n_134),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_48),
.C(n_42),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_59),
.B1(n_25),
.B2(n_33),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_138),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_59),
.B1(n_19),
.B2(n_21),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_86),
.B1(n_103),
.B2(n_108),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_42),
.C(n_41),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_138),
.B(n_129),
.Y(n_175)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_106),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_97),
.A2(n_41),
.B(n_39),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_37),
.B(n_39),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_170),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_149),
.A2(n_151),
.B1(n_154),
.B2(n_176),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_98),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g201 ( 
.A(n_150),
.B(n_157),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_95),
.B1(n_75),
.B2(n_114),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_95),
.B(n_85),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_152),
.A2(n_172),
.B(n_1),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_87),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_171),
.C(n_142),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_122),
.B1(n_128),
.B2(n_116),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_81),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_164),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_166),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_82),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_112),
.B1(n_104),
.B2(n_91),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_119),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_104),
.B1(n_90),
.B2(n_78),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_109),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_100),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_92),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_37),
.C(n_38),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_177),
.B1(n_121),
.B2(n_120),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_109),
.B1(n_39),
.B2(n_37),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_37),
.B1(n_21),
.B2(n_19),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_181),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_33),
.A3(n_19),
.B1(n_21),
.B2(n_31),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_188),
.C(n_202),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_187),
.B1(n_189),
.B2(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_121),
.B1(n_118),
.B2(n_127),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_130),
.C(n_121),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_127),
.B1(n_120),
.B2(n_31),
.Y(n_189)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_31),
.B1(n_89),
.B2(n_76),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_209),
.B1(n_5),
.B2(n_8),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_31),
.B(n_1),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_8),
.B(n_9),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_0),
.C(n_1),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_152),
.B1(n_157),
.B2(n_149),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_8),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_177),
.B1(n_146),
.B2(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_222),
.B1(n_235),
.B2(n_200),
.Y(n_251)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_203),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_158),
.B1(n_151),
.B2(n_157),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_223),
.B1(n_180),
.B2(n_183),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_153),
.B1(n_167),
.B2(n_168),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_147),
.C(n_159),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_228),
.C(n_232),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_11),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_202),
.C(n_209),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_5),
.C(n_6),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_180),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_208),
.B1(n_210),
.B2(n_186),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_5),
.C(n_7),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

OA21x2_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_201),
.B(n_207),
.Y(n_244)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_191),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_245),
.A2(n_260),
.B1(n_211),
.B2(n_234),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_192),
.C(n_179),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_252),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_192),
.C(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_237),
.B1(n_228),
.B2(n_214),
.Y(n_281)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_201),
.C(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_259),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_190),
.CI(n_193),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_190),
.C(n_191),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_181),
.B1(n_178),
.B2(n_199),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_253),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_223),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_276),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_266),
.B(n_239),
.Y(n_292)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_280),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_215),
.B1(n_226),
.B2(n_213),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_273),
.B1(n_281),
.B2(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_254),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_215),
.B1(n_221),
.B2(n_216),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_221),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_235),
.B(n_218),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_252),
.B(n_245),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_232),
.Y(n_280)
);

OA21x2_ASAP7_75t_SL g282 ( 
.A1(n_279),
.A2(n_259),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_261),
.C(n_246),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_286),
.C(n_287),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_249),
.C(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_293),
.C(n_297),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_269),
.B1(n_274),
.B2(n_277),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_9),
.B(n_12),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_242),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_265),
.B1(n_276),
.B2(n_280),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_241),
.C(n_9),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_281),
.B(n_264),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_296),
.C(n_283),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_309),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_293),
.B1(n_286),
.B2(n_288),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_291),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_290),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_291),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_296),
.C(n_14),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_309),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_301),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_320),
.A2(n_321),
.B(n_307),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_308),
.B(n_301),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_326),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_302),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_304),
.B(n_300),
.C(n_307),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_325),
.A2(n_298),
.B(n_317),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_330),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_323),
.B(n_332),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_329),
.C(n_319),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_320),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_15),
.Y(n_337)
);


endmodule