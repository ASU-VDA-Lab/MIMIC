module fake_jpeg_21683_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx11_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_5),
.B(n_4),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_3),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_6),
.C(n_10),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_13),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_13),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_6),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_7),
.B1(n_24),
.B2(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.C(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_29),
.B1(n_17),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_16),
.A2(n_7),
.B1(n_9),
.B2(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.C(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_33),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_40),
.B(n_29),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_27),
.B(n_30),
.C(n_37),
.D(n_36),
.Y(n_44)
);


endmodule