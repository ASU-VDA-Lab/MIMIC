module fake_netlist_5_770_n_88 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_88);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_88;

wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_15),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

OAI22x1_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_14),
.B1(n_4),
.B2(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_2),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_3),
.B1(n_9),
.B2(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AO32x2_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_31),
.A3(n_28),
.B1(n_33),
.B2(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_26),
.B(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_34),
.B(n_21),
.C(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_42),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_43),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_40),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NAND2x1_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_53),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_41),
.B1(n_21),
.B2(n_30),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI221xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_28),
.B1(n_55),
.B2(n_38),
.C(n_29),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_25),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_29),
.B1(n_31),
.B2(n_24),
.C(n_27),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_32),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_65),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_32),
.B(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_32),
.Y(n_79)
);

AOI211xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_32),
.B(n_20),
.C(n_22),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_75),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_80),
.B1(n_79),
.B2(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

OAI22x1_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_83),
.B1(n_77),
.B2(n_22),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_20),
.B(n_22),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_22),
.B(n_86),
.Y(n_88)
);


endmodule