module fake_netlist_5_289_n_1938 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1938);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1938;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_74),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_176),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_149),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_78),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_67),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_30),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_30),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_87),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_0),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_34),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_72),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_66),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_106),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_68),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_128),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_57),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_73),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_132),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_13),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_29),
.Y(n_218)
);

BUFx8_ASAP7_75t_SL g219 ( 
.A(n_156),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_90),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_28),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_42),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_21),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_104),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_108),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_3),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_138),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_81),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_51),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_165),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_21),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_9),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_62),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_70),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_99),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_94),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_39),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_65),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_24),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_31),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_118),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_55),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_25),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_158),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_79),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_26),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_46),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_38),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_177),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_33),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_61),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_129),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_174),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_33),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_12),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_47),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_96),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_83),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_54),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_39),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_9),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_120),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_71),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_140),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_14),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_17),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_85),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_48),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_60),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_146),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_6),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_112),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_141),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_114),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_103),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_139),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_180),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_167),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_16),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_168),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_7),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_119),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_10),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_101),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_23),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_105),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_122),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_109),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_163),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_20),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_178),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_157),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_31),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_89),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_20),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_97),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_53),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_46),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_124),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_15),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_86),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_54),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_121),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_123),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_2),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_12),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_37),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_115),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_117),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_82),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_61),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_102),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_5),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_91),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_53),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_162),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_113),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_154),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_18),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_56),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_77),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_60),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_150),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_57),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_14),
.Y(n_346)
);

BUFx8_ASAP7_75t_SL g347 ( 
.A(n_172),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_136),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_18),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_1),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_45),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_130),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_164),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_137),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_40),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_133),
.Y(n_356)
);

CKINVDCx6p67_ASAP7_75t_R g357 ( 
.A(n_80),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_48),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_37),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_44),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_281),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_208),
.B(n_179),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_261),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_257),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_218),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_190),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_261),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_221),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_298),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_226),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_2),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_261),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_227),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_228),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_261),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_238),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_231),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_235),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_236),
.Y(n_382)
);

INVx4_ASAP7_75t_R g383 ( 
.A(n_183),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_329),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_270),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_219),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_261),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_293),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_261),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_181),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_247),
.B(n_3),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_182),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_242),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_246),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_191),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_261),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_213),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_250),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_255),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_261),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_283),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_264),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_295),
.Y(n_404)
);

BUFx6f_ASAP7_75t_SL g405 ( 
.A(n_183),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_258),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_283),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_273),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_278),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_212),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_283),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_284),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_283),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_283),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_287),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_215),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_193),
.B(n_4),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_283),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_302),
.B(n_4),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_283),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_191),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_220),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_225),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_283),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_286),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_286),
.B(n_7),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_289),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_286),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_286),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_286),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_286),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_229),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_230),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_286),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_299),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_233),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_286),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_186),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_234),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_305),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_214),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_302),
.B(n_8),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_214),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_315),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_318),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_214),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_214),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_322),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_383),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_444),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_427),
.A2(n_256),
.B(n_247),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_419),
.B(n_214),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_396),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_328),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_373),
.B(n_208),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_373),
.B(n_186),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_364),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_276),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_369),
.A2(n_304),
.B(n_192),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_374),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_365),
.B(n_328),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_377),
.B(n_320),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_363),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_380),
.B(n_276),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_363),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_371),
.B(n_320),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_363),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_363),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_413),
.B(n_304),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_414),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_422),
.B(n_197),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_417),
.B(n_208),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_425),
.B(n_320),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_384),
.B(n_320),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_363),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_361),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_429),
.Y(n_496)
);

BUFx8_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_430),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_435),
.B(n_320),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_366),
.B(n_339),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_184),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_392),
.B(n_339),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_391),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_393),
.B(n_339),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_366),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_370),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_370),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_375),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_375),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_416),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_376),
.B(n_339),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_376),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_379),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_379),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_381),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_381),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_403),
.B(n_208),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_362),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_382),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_382),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_523),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_459),
.A2(n_199),
.B1(n_292),
.B2(n_280),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_423),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_451),
.B(n_398),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_450),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_196),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_495),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_470),
.B(n_399),
.C(n_395),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_488),
.Y(n_544)
);

OAI22x1_ASAP7_75t_L g545 ( 
.A1(n_457),
.A2(n_271),
.B1(n_359),
.B2(n_355),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_510),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_502),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_452),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_503),
.B(n_195),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_452),
.Y(n_553)
);

AND3x2_ASAP7_75t_L g554 ( 
.A(n_458),
.B(n_268),
.C(n_256),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_395),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_456),
.A2(n_202),
.B(n_200),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_495),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_453),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_509),
.B(n_424),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_464),
.B(n_399),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_509),
.B(n_433),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_488),
.A2(n_339),
.B1(n_345),
.B2(n_313),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_463),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_464),
.B(n_400),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_461),
.B(n_206),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_482),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_488),
.A2(n_345),
.B1(n_313),
.B2(n_268),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_467),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_451),
.B(n_400),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_515),
.B(n_406),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_473),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_487),
.B(n_404),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_451),
.B(n_406),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_482),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_507),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_474),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_487),
.B(n_408),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_434),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_507),
.B(n_408),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_482),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_490),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_474),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_475),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_507),
.B(n_409),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_467),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_475),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_519),
.B(n_409),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_515),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_519),
.B(n_412),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_467),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_490),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_477),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_461),
.B(n_210),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_476),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_456),
.A2(n_266),
.B1(n_360),
.B2(n_358),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_511),
.B(n_437),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_484),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_484),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_496),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_496),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_477),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_486),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_486),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_519),
.B(n_412),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_462),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_515),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_501),
.B(n_415),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_471),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_489),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_489),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_498),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_498),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_494),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_512),
.B(n_386),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_494),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_462),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_487),
.B(n_415),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_470),
.B(n_436),
.C(n_428),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_494),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_461),
.B(n_211),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_477),
.B(n_208),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_494),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_494),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_465),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_522),
.B(n_428),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_471),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_465),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_466),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_516),
.B(n_440),
.Y(n_643)
);

INVx11_ASAP7_75t_L g644 ( 
.A(n_497),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_510),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_480),
.B(n_436),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_466),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_491),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_468),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_454),
.A2(n_260),
.B1(n_223),
.B2(n_232),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_441),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_465),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_454),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_501),
.B(n_441),
.Y(n_655)
);

AND3x2_ASAP7_75t_L g656 ( 
.A(n_458),
.B(n_237),
.C(n_224),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_477),
.Y(n_657)
);

AO21x2_ASAP7_75t_L g658 ( 
.A1(n_491),
.A2(n_243),
.B(n_241),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_454),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_454),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_454),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_481),
.B(n_252),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_502),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_517),
.B(n_445),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_461),
.B(n_269),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_503),
.B(n_282),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_468),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_502),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_481),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_517),
.B(n_445),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_480),
.B(n_492),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_502),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_510),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_502),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_500),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_460),
.A2(n_310),
.B1(n_217),
.B2(n_240),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_481),
.B(n_288),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_492),
.B(n_446),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_485),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_668),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_557),
.B(n_478),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_574),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_SL g684 ( 
.A(n_574),
.B(n_481),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_544),
.B(n_519),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_576),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_544),
.B(n_506),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_668),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_667),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_671),
.B(n_506),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_596),
.B(n_508),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_668),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_667),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_576),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_528),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_596),
.B(n_508),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_678),
.B(n_508),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_667),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_552),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_671),
.B(n_506),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_672),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_621),
.B(n_506),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_534),
.B(n_503),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_620),
.B(n_527),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_457),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_672),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_574),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_582),
.B(n_520),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_639),
.B(n_506),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_551),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_649),
.B(n_506),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_663),
.B(n_519),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_663),
.B(n_519),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_663),
.B(n_519),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_531),
.B(n_513),
.C(n_524),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_571),
.A2(n_566),
.B1(n_675),
.B2(n_649),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_655),
.B(n_527),
.Y(n_718)
);

BUFx6f_ASAP7_75t_SL g719 ( 
.A(n_552),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_534),
.B(n_520),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_675),
.B(n_506),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_SL g722 ( 
.A(n_540),
.B(n_527),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_663),
.B(n_527),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_546),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_579),
.B(n_520),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_680),
.A2(n_651),
.B1(n_661),
.B2(n_558),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_680),
.B(n_526),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_582),
.B(n_526),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_619),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_574),
.B(n_601),
.Y(n_730)
);

BUFx8_ASAP7_75t_L g731 ( 
.A(n_557),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_564),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_564),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_530),
.B(n_524),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_530),
.B(n_524),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_645),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_543),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_553),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_674),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_574),
.B(n_527),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_619),
.A2(n_527),
.B1(n_524),
.B2(n_512),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_587),
.A2(n_525),
.B1(n_518),
.B2(n_522),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_534),
.B(n_505),
.Y(n_743)
);

BUFx4f_ASAP7_75t_L g744 ( 
.A(n_552),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_539),
.B(n_527),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_553),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_574),
.B(n_479),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_652),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_592),
.B(n_518),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_543),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_555),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_601),
.B(n_479),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_601),
.B(n_479),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_568),
.B(n_478),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_679),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_539),
.B(n_512),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_542),
.B(n_512),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_SL g758 ( 
.A(n_559),
.B(n_512),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_542),
.B(n_522),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_679),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_572),
.B(n_522),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_572),
.B(n_522),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_577),
.B(n_522),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_543),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_577),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_555),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_578),
.B(n_522),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_578),
.B(n_522),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_664),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_561),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_561),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_583),
.B(n_522),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_583),
.B(n_590),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_601),
.B(n_479),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_590),
.B(n_591),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_533),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_591),
.B(n_460),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_594),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_594),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_568),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_605),
.B(n_460),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_605),
.B(n_460),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_647),
.B(n_513),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_647),
.B(n_670),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_608),
.B(n_460),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_541),
.B(n_389),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_460),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_533),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_631),
.B(n_595),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_601),
.B(n_479),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_597),
.B(n_446),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_610),
.B(n_460),
.Y(n_792)
);

INVx8_ASAP7_75t_L g793 ( 
.A(n_552),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_610),
.B(n_460),
.Y(n_794)
);

BUFx8_ASAP7_75t_L g795 ( 
.A(n_534),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_611),
.B(n_460),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_611),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_615),
.B(n_485),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_617),
.B(n_449),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_584),
.A2(n_385),
.B1(n_388),
.B2(n_378),
.Y(n_800)
);

O2A1O1Ixp5_ASAP7_75t_L g801 ( 
.A1(n_661),
.A2(n_485),
.B(n_504),
.C(n_478),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_615),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_533),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_563),
.B(n_449),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_616),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_538),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_616),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_601),
.B(n_481),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_622),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_538),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_607),
.B(n_481),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_538),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_622),
.B(n_485),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_630),
.B(n_521),
.C(n_514),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_623),
.B(n_624),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_623),
.B(n_485),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_624),
.B(n_505),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_627),
.B(n_497),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_625),
.B(n_481),
.Y(n_819)
);

INVx8_ASAP7_75t_L g820 ( 
.A(n_552),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_550),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_550),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_L g823 ( 
.A(n_565),
.B(n_609),
.C(n_586),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_625),
.B(n_483),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_580),
.B(n_222),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_643),
.B(n_514),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_618),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_554),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_607),
.B(n_483),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_661),
.B(n_483),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_673),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_618),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_529),
.B(n_514),
.Y(n_833)
);

AO22x2_ASAP7_75t_L g834 ( 
.A1(n_654),
.A2(n_660),
.B1(n_659),
.B2(n_569),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_607),
.B(n_483),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_629),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_545),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_549),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_569),
.B(n_483),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_569),
.B(n_483),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_545),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_629),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_641),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_558),
.A2(n_245),
.B1(n_335),
.B2(n_272),
.Y(n_844)
);

AOI221xp5_ASAP7_75t_L g845 ( 
.A1(n_529),
.A2(n_251),
.B1(n_346),
.B2(n_359),
.C(n_201),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_641),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_569),
.B(n_602),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_548),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_784),
.A2(n_606),
.B(n_660),
.C(n_659),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_737),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_717),
.A2(n_549),
.B1(n_654),
.B2(n_660),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_795),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_784),
.A2(n_638),
.B(n_504),
.C(n_648),
.Y(n_853)
);

NOR2x1_ASAP7_75t_L g854 ( 
.A(n_741),
.B(n_521),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_838),
.B(n_607),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_747),
.A2(n_562),
.B(n_547),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_682),
.B(n_521),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_695),
.B(n_367),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_747),
.A2(n_562),
.B(n_547),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_752),
.A2(n_562),
.B(n_547),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_748),
.B(n_368),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_717),
.A2(n_549),
.B1(n_654),
.B2(n_660),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_848),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_752),
.A2(n_562),
.B(n_547),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_697),
.B(n_548),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_L g866 ( 
.A(n_724),
.B(n_602),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_697),
.B(n_691),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_754),
.B(n_372),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_753),
.A2(n_598),
.B(n_573),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_795),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_753),
.A2(n_598),
.B(n_573),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_691),
.B(n_548),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_774),
.A2(n_598),
.B(n_573),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_696),
.B(n_604),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_726),
.A2(n_659),
.B(n_654),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_769),
.B(n_532),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_774),
.A2(n_598),
.B(n_573),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_790),
.A2(n_657),
.B(n_614),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_604),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_790),
.A2(n_657),
.B(n_614),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_727),
.B(n_604),
.Y(n_881)
);

BUFx8_ASAP7_75t_L g882 ( 
.A(n_831),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_789),
.A2(n_602),
.B1(n_633),
.B2(n_665),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_736),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_690),
.A2(n_659),
.B(n_633),
.C(n_665),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_700),
.B(n_708),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_783),
.B(n_602),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_708),
.B(n_728),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_737),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_743),
.B(n_666),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_808),
.A2(n_657),
.B(n_614),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_702),
.A2(n_709),
.B(n_657),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_749),
.A2(n_728),
.B(n_685),
.C(n_783),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_749),
.B(n_633),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_683),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_804),
.B(n_633),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_839),
.A2(n_614),
.B(n_607),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_840),
.A2(n_614),
.B(n_607),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_765),
.B(n_778),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_L g900 ( 
.A1(n_825),
.A2(n_201),
.B(n_194),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_683),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_750),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_847),
.A2(n_669),
.B(n_614),
.Y(n_903)
);

CKINVDCx8_ASAP7_75t_R g904 ( 
.A(n_793),
.Y(n_904)
);

INVx11_ASAP7_75t_L g905 ( 
.A(n_731),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_789),
.A2(n_665),
.B1(n_549),
.B2(n_575),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_686),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_681),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_740),
.A2(n_669),
.B(n_640),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_740),
.A2(n_669),
.B(n_640),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_683),
.A2(n_669),
.B(n_640),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_683),
.A2(n_669),
.B(n_640),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_826),
.B(n_665),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_685),
.A2(n_650),
.B(n_648),
.C(n_632),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_793),
.B(n_666),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_779),
.B(n_628),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_797),
.B(n_628),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_802),
.B(n_628),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_707),
.A2(n_669),
.B(n_653),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_707),
.A2(n_730),
.B(n_721),
.Y(n_920)
);

BUFx8_ASAP7_75t_SL g921 ( 
.A(n_833),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_707),
.A2(n_653),
.B(n_637),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_800),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_726),
.A2(n_711),
.B1(n_687),
.B2(n_729),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_688),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_725),
.B(n_628),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_705),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_732),
.B(n_626),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_733),
.B(n_656),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_684),
.A2(n_829),
.B(n_811),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_694),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_692),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_805),
.B(n_558),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_807),
.B(n_650),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_707),
.A2(n_653),
.B(n_637),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_750),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_773),
.A2(n_626),
.B(n_632),
.C(n_666),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_809),
.B(n_635),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_701),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_704),
.A2(n_294),
.B(n_291),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_635),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_706),
.Y(n_942)
);

AND2x2_ASAP7_75t_SL g943 ( 
.A(n_823),
.B(n_300),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_730),
.A2(n_653),
.B(n_637),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_739),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_713),
.A2(n_637),
.B(n_593),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_720),
.A2(n_666),
.B1(n_658),
.B2(n_677),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_815),
.B(n_635),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_734),
.B(n_636),
.Y(n_949)
);

NOR2x1_ASAP7_75t_L g950 ( 
.A(n_786),
.B(n_666),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_713),
.A2(n_593),
.B(n_585),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_755),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_689),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_780),
.B(n_825),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_735),
.B(n_636),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_689),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_720),
.B(n_636),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_714),
.A2(n_593),
.B(n_585),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_764),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_845),
.A2(n_303),
.B(n_249),
.C(n_317),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_714),
.A2(n_593),
.B(n_585),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_715),
.A2(n_593),
.B(n_585),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_791),
.B(n_253),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_791),
.A2(n_203),
.B(n_194),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_799),
.A2(n_267),
.B(n_244),
.C(n_341),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_799),
.A2(n_326),
.B(n_349),
.C(n_323),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_756),
.B(n_556),
.Y(n_967)
);

NOR2x1_ASAP7_75t_L g968 ( 
.A(n_818),
.B(n_658),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_693),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_764),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_757),
.B(n_556),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_760),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_837),
.B(n_263),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_745),
.B(n_556),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_832),
.B(n_556),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_L g976 ( 
.A(n_716),
.B(n_308),
.C(n_209),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_715),
.A2(n_593),
.B(n_585),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_723),
.A2(n_642),
.B(n_585),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_723),
.A2(n_646),
.B(n_642),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_560),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_843),
.B(n_560),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_843),
.B(n_560),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_L g983 ( 
.A(n_841),
.B(n_758),
.C(n_814),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_846),
.B(n_560),
.Y(n_984)
);

AO21x1_ASAP7_75t_L g985 ( 
.A1(n_718),
.A2(n_306),
.B(n_307),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_801),
.A2(n_588),
.B(n_600),
.Y(n_986)
);

AO21x1_ASAP7_75t_L g987 ( 
.A1(n_759),
.A2(n_309),
.B(n_312),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_811),
.A2(n_646),
.B(n_642),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_742),
.B(n_483),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_SL g990 ( 
.A1(n_777),
.A2(n_332),
.B(n_353),
.C(n_354),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_761),
.A2(n_600),
.B(n_599),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_829),
.A2(n_646),
.B(n_642),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_835),
.A2(n_646),
.B(n_642),
.Y(n_993)
);

NOR2x1_ASAP7_75t_R g994 ( 
.A(n_828),
.B(n_203),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_835),
.A2(n_642),
.B(n_646),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_744),
.B(n_838),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_846),
.B(n_603),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_798),
.A2(n_816),
.B(n_813),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_698),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_731),
.Y(n_1000)
);

AO21x1_ASAP7_75t_L g1001 ( 
.A1(n_762),
.A2(n_589),
.B(n_567),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_817),
.B(n_827),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_836),
.B(n_603),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_819),
.A2(n_646),
.B(n_589),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_824),
.A2(n_612),
.B(n_570),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_763),
.A2(n_612),
.B(n_570),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_848),
.B(n_658),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_842),
.B(n_603),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_710),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_767),
.A2(n_567),
.B(n_588),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_710),
.Y(n_1011)
);

OAI321xp33_ASAP7_75t_L g1012 ( 
.A1(n_844),
.A2(n_676),
.A3(n_301),
.B1(n_295),
.B2(n_271),
.C(n_350),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_744),
.B(n_581),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_699),
.B(n_719),
.Y(n_1014)
);

BUFx4f_ASAP7_75t_L g1015 ( 
.A(n_793),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_768),
.A2(n_600),
.B(n_581),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_698),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_834),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_743),
.B(n_331),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_712),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_844),
.B(n_603),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_703),
.B(n_295),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_SL g1023 ( 
.A(n_699),
.B(n_497),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_703),
.A2(n_677),
.B1(n_662),
.B2(n_493),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_834),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_772),
.A2(n_599),
.B(n_588),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_781),
.A2(n_581),
.B(n_599),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_782),
.A2(n_787),
.B(n_785),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_719),
.B(n_644),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_792),
.A2(n_613),
.B(n_535),
.C(n_536),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_712),
.B(n_613),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_738),
.B(n_613),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_722),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_794),
.A2(n_613),
.B(n_536),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_738),
.B(n_535),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_796),
.A2(n_535),
.B(n_536),
.Y(n_1036)
);

OR2x6_ASAP7_75t_SL g1037 ( 
.A(n_746),
.B(n_331),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_954),
.B(n_820),
.Y(n_1038)
);

AO21x1_ASAP7_75t_L g1039 ( 
.A1(n_893),
.A2(n_770),
.B(n_746),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_892),
.A2(n_834),
.B(n_751),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_1015),
.B(n_751),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_953),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_963),
.A2(n_861),
.B(n_927),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_963),
.B(n_766),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_858),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_998),
.A2(n_770),
.B(n_771),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_960),
.A2(n_771),
.B(n_766),
.C(n_822),
.Y(n_1047)
);

INVx3_ASAP7_75t_SL g1048 ( 
.A(n_884),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_908),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_895),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_886),
.A2(n_806),
.B(n_788),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_956),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_849),
.A2(n_776),
.B(n_788),
.C(n_803),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_868),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_888),
.B(n_830),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_867),
.B(n_830),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_890),
.B(n_821),
.Y(n_1057)
);

OAI21xp33_ASAP7_75t_SL g1058 ( 
.A1(n_894),
.A2(n_822),
.B(n_821),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_907),
.Y(n_1059)
);

CKINVDCx12_ASAP7_75t_R g1060 ( 
.A(n_857),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_907),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_875),
.A2(n_803),
.B(n_812),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_861),
.B(n_820),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_887),
.B(n_830),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1002),
.B(n_830),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_891),
.A2(n_820),
.B(n_830),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_858),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_896),
.B(n_943),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_1029),
.B(n_239),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_876),
.B(n_644),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_931),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_L g1072 ( 
.A1(n_940),
.A2(n_812),
.B(n_810),
.C(n_806),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1022),
.B(n_301),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_872),
.A2(n_776),
.B(n_810),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1002),
.B(n_535),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_926),
.B(n_536),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_926),
.B(n_537),
.Y(n_1077)
);

INVx3_ASAP7_75t_SL g1078 ( 
.A(n_852),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_L g1079 ( 
.A(n_964),
.B(n_325),
.C(n_327),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_895),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_913),
.B(n_537),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_856),
.A2(n_537),
.B(n_493),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_883),
.A2(n_493),
.B1(n_357),
.B2(n_189),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_874),
.A2(n_537),
.B(n_248),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_853),
.A2(n_185),
.B(n_189),
.C(n_198),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_943),
.A2(n_321),
.B1(n_254),
.B2(n_259),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_876),
.A2(n_185),
.B(n_198),
.C(n_204),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_931),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_865),
.B(n_634),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_969),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_973),
.B(n_301),
.Y(n_1091)
);

BUFx2_ASAP7_75t_SL g1092 ( 
.A(n_866),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_923),
.B(n_340),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_895),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_906),
.A2(n_493),
.B1(n_357),
.B2(n_204),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_890),
.B(n_497),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_976),
.A2(n_334),
.B(n_207),
.C(n_330),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_879),
.A2(n_262),
.B(n_265),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_973),
.B(n_340),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_R g1100 ( 
.A(n_904),
.B(n_497),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_899),
.B(n_634),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_851),
.A2(n_274),
.B(n_275),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_L g1103 ( 
.A(n_959),
.B(n_277),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_945),
.B(n_928),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_999),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1017),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_882),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_960),
.A2(n_343),
.B(n_350),
.C(n_351),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_985),
.A2(n_677),
.B(n_662),
.C(n_634),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1000),
.A2(n_343),
.B1(n_351),
.B2(n_355),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_933),
.A2(n_677),
.B(n_662),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1020),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_854),
.B(n_959),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_966),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_849),
.A2(n_677),
.B(n_662),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_945),
.A2(n_493),
.B1(n_205),
.B2(n_334),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_900),
.B(n_970),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_862),
.A2(n_279),
.B(n_285),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_882),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_1023),
.B(n_205),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_928),
.B(n_634),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1014),
.A2(n_207),
.B1(n_356),
.B2(n_352),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_970),
.B(n_330),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_924),
.A2(n_290),
.B(n_296),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_976),
.B(n_338),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_885),
.A2(n_297),
.B(n_311),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_881),
.B(n_634),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1015),
.B(n_342),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_952),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_921),
.B(n_338),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_925),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_983),
.B(n_850),
.Y(n_1132)
);

AOI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_1019),
.A2(n_337),
.B(n_352),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_921),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_932),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_SL g1136 ( 
.A1(n_989),
.A2(n_677),
.B(n_662),
.C(n_634),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_895),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_972),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1037),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_852),
.B(n_342),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_983),
.A2(n_314),
.B1(n_316),
.B2(n_319),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1018),
.A2(n_493),
.B1(n_336),
.B2(n_337),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1018),
.A2(n_1025),
.B1(n_1033),
.B2(n_1021),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_937),
.A2(n_348),
.B(n_336),
.C(n_344),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_850),
.B(n_634),
.Y(n_1145)
);

NAND2x1p5_ASAP7_75t_L g1146 ( 
.A(n_901),
.B(n_677),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_863),
.B(n_662),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_859),
.A2(n_324),
.B(n_356),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_885),
.A2(n_989),
.B(n_920),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_901),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_967),
.A2(n_348),
.B(n_344),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1009),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_965),
.A2(n_16),
.B(n_19),
.Y(n_1153)
);

BUFx2_ASAP7_75t_R g1154 ( 
.A(n_870),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_915),
.B(n_134),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1012),
.A2(n_662),
.B(n_22),
.C(n_23),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_863),
.B(n_19),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_905),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_994),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_860),
.A2(n_170),
.B(n_169),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_966),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_864),
.A2(n_166),
.B(n_153),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1011),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_889),
.B(n_148),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_SL g1165 ( 
.A(n_870),
.B(n_147),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_965),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_929),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_996),
.A2(n_144),
.B1(n_143),
.B2(n_142),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1014),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1029),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_889),
.B(n_902),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_902),
.B(n_27),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_936),
.B(n_127),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1025),
.B(n_32),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_SL g1175 ( 
.A1(n_1030),
.A2(n_116),
.B(n_100),
.C(n_98),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_936),
.B(n_88),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_916),
.A2(n_84),
.B1(n_76),
.B2(n_75),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_934),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_901),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_947),
.A2(n_914),
.B(n_968),
.C(n_1028),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_915),
.B(n_63),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_1001),
.A2(n_32),
.B(n_35),
.C(n_36),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_915),
.B(n_35),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_996),
.B(n_36),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_939),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1027),
.A2(n_38),
.B(n_40),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_971),
.A2(n_42),
.B(n_43),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_922),
.A2(n_43),
.B(n_44),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_942),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_R g1190 ( 
.A(n_901),
.B(n_59),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_950),
.B(n_957),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_935),
.A2(n_45),
.B(n_49),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_974),
.A2(n_49),
.B(n_50),
.Y(n_1193)
);

BUFx2_ASAP7_75t_SL g1194 ( 
.A(n_1013),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_903),
.A2(n_52),
.B(n_56),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_930),
.B(n_52),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1180),
.A2(n_873),
.B(n_877),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1149),
.A2(n_871),
.B(n_869),
.Y(n_1198)
);

OAI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1093),
.A2(n_1013),
.B1(n_1007),
.B2(n_917),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1049),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1043),
.B(n_918),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_SL g1202 ( 
.A(n_1100),
.B(n_948),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1149),
.A2(n_880),
.B(n_878),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1050),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1054),
.B(n_941),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1104),
.A2(n_919),
.B(n_912),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1178),
.B(n_938),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1156),
.A2(n_955),
.B(n_949),
.C(n_1003),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1039),
.A2(n_987),
.A3(n_910),
.B(n_909),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1044),
.B(n_1032),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1046),
.A2(n_911),
.B(n_944),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1048),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1067),
.B(n_855),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1046),
.A2(n_1040),
.B(n_1066),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1040),
.A2(n_986),
.B(n_898),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1099),
.B(n_1008),
.Y(n_1216)
);

AOI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1117),
.A2(n_981),
.B(n_980),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1065),
.A2(n_897),
.B(n_946),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1056),
.A2(n_991),
.B(n_1006),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1085),
.A2(n_1026),
.A3(n_1016),
.B(n_1010),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1061),
.B(n_982),
.Y(n_1221)
);

INVx3_ASAP7_75t_SL g1222 ( 
.A(n_1158),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1144),
.A2(n_1005),
.A3(n_1034),
.B(n_1036),
.Y(n_1223)
);

AOI221x1_ASAP7_75t_L g1224 ( 
.A1(n_1153),
.A2(n_1004),
.B1(n_1031),
.B2(n_984),
.C(n_997),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1055),
.A2(n_975),
.B(n_1035),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1075),
.A2(n_978),
.B(n_979),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1167),
.Y(n_1227)
);

OAI21xp33_ASAP7_75t_L g1228 ( 
.A1(n_1091),
.A2(n_1024),
.B(n_855),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1108),
.A2(n_977),
.B(n_962),
.C(n_951),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1132),
.A2(n_990),
.B(n_961),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1071),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1129),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_1084),
.A2(n_990),
.B(n_958),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1143),
.A2(n_988),
.A3(n_992),
.B(n_993),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1084),
.A2(n_995),
.A3(n_58),
.B(n_59),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1150),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1070),
.B(n_1063),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1138),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1073),
.B(n_1123),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1184),
.B(n_1088),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1152),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1111),
.A2(n_1074),
.B(n_1062),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1076),
.A2(n_1077),
.B(n_1089),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1068),
.B(n_1059),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1184),
.B(n_1170),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1074),
.A2(n_1062),
.B(n_1051),
.Y(n_1246)
);

AO21x1_ASAP7_75t_L g1247 ( 
.A1(n_1195),
.A2(n_1188),
.B(n_1192),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1078),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1119),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1045),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1051),
.A2(n_1191),
.B(n_1127),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1082),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1126),
.A2(n_1195),
.A3(n_1095),
.B(n_1192),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1115),
.A2(n_1072),
.B(n_1047),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1064),
.A2(n_1113),
.B(n_1081),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_SL g1256 ( 
.A1(n_1175),
.A2(n_1164),
.B(n_1176),
.C(n_1173),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1121),
.A2(n_1101),
.B(n_1150),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1169),
.B(n_1185),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1154),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1166),
.A2(n_1114),
.B1(n_1161),
.B2(n_1187),
.C(n_1193),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1126),
.A2(n_1188),
.A3(n_1124),
.B(n_1083),
.Y(n_1261)
);

OAI22x1_ASAP7_75t_L g1262 ( 
.A1(n_1174),
.A2(n_1139),
.B1(n_1183),
.B2(n_1125),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1057),
.B(n_1189),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1133),
.A2(n_1097),
.B(n_1087),
.C(n_1079),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1130),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1042),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1157),
.A2(n_1172),
.B(n_1038),
.C(n_1147),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1124),
.A2(n_1118),
.B(n_1102),
.C(n_1151),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1057),
.A2(n_1194),
.B1(n_1135),
.B2(n_1131),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1140),
.B(n_1120),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1102),
.A2(n_1118),
.B(n_1098),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1171),
.B(n_1163),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1150),
.A2(n_1162),
.B(n_1160),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_R g1274 ( 
.A(n_1060),
.B(n_1107),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1098),
.A2(n_1151),
.B(n_1148),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1112),
.B(n_1105),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1052),
.B(n_1106),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1086),
.A2(n_1141),
.B(n_1187),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1122),
.B(n_1128),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1165),
.A2(n_1183),
.B1(n_1096),
.B2(n_1155),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1090),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1150),
.A2(n_1145),
.B(n_1136),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1177),
.A2(n_1109),
.B(n_1041),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1134),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1159),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1190),
.B(n_1069),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1155),
.A2(n_1181),
.B(n_1168),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1094),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1050),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1155),
.B(n_1181),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1193),
.A2(n_1182),
.B(n_1142),
.C(n_1116),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1050),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1181),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1186),
.A2(n_1041),
.B(n_1146),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1080),
.B(n_1179),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_SL g1296 ( 
.A1(n_1094),
.A2(n_1137),
.B(n_1196),
.C(n_1146),
.Y(n_1296)
);

AOI221x1_ASAP7_75t_L g1297 ( 
.A1(n_1110),
.A2(n_1137),
.B1(n_1092),
.B2(n_1080),
.C(n_1179),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1103),
.A2(n_823),
.B(n_963),
.C(n_784),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1155),
.B(n_1181),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1099),
.A2(n_963),
.B1(n_823),
.B2(n_943),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_784),
.B(n_893),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1099),
.A2(n_784),
.B(n_963),
.C(n_789),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1049),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1180),
.A2(n_892),
.B(n_709),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1180),
.A2(n_892),
.B(n_709),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1178),
.B(n_784),
.Y(n_1307)
);

BUFx10_ASAP7_75t_L g1308 ( 
.A(n_1130),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1048),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1119),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1043),
.B(n_963),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1104),
.A2(n_784),
.B1(n_963),
.B2(n_888),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1048),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1119),
.Y(n_1316)
);

INVx3_ASAP7_75t_SL g1317 ( 
.A(n_1048),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1039),
.A2(n_1180),
.A3(n_987),
.B(n_1001),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1049),
.Y(n_1319)
);

OAI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1099),
.A2(n_963),
.B(n_784),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1039),
.A2(n_1180),
.A3(n_987),
.B(n_1001),
.Y(n_1321)
);

AO32x2_ASAP7_75t_L g1322 ( 
.A1(n_1143),
.A2(n_924),
.A3(n_1095),
.B1(n_1083),
.B2(n_1142),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1049),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1061),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1178),
.B(n_784),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_SL g1326 ( 
.A1(n_1188),
.A2(n_1192),
.B(n_1195),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1099),
.A2(n_963),
.B1(n_784),
.B2(n_823),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1049),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1150),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1178),
.B(n_784),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_L g1331 ( 
.A(n_1099),
.B(n_823),
.C(n_784),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1057),
.B(n_890),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1180),
.A2(n_892),
.B(n_709),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1049),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1155),
.B(n_1181),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1048),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1180),
.A2(n_784),
.B(n_893),
.Y(n_1338)
);

O2A1O1Ixp5_ASAP7_75t_L g1339 ( 
.A1(n_1124),
.A2(n_784),
.B(n_818),
.C(n_963),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1043),
.A2(n_823),
.B(n_963),
.C(n_784),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1057),
.B(n_890),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1180),
.A2(n_784),
.B(n_893),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1057),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1180),
.A2(n_892),
.B(n_709),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1046),
.A2(n_1111),
.B(n_1074),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1061),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1054),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1048),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1178),
.B(n_784),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1040),
.A2(n_1149),
.B(n_1111),
.Y(n_1352)
);

BUFx4_ASAP7_75t_SL g1353 ( 
.A(n_1107),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1180),
.A2(n_784),
.B(n_893),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1178),
.B(n_784),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1099),
.A2(n_784),
.B(n_963),
.C(n_789),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1048),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1180),
.A2(n_892),
.B(n_709),
.Y(n_1358)
);

INVx6_ASAP7_75t_L g1359 ( 
.A(n_1236),
.Y(n_1359)
);

INVx6_ASAP7_75t_L g1360 ( 
.A(n_1236),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1310),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1311),
.A2(n_1300),
.B1(n_1320),
.B2(n_1327),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1200),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1327),
.A2(n_1237),
.B1(n_1270),
.B2(n_1314),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1316),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1331),
.A2(n_1354),
.B1(n_1344),
.B2(n_1338),
.Y(n_1366)
);

CKINVDCx6p67_ASAP7_75t_R g1367 ( 
.A(n_1317),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1331),
.A2(n_1336),
.B1(n_1299),
.B2(n_1280),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1329),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1329),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1320),
.A2(n_1341),
.B(n_1279),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1302),
.A2(n_1356),
.B1(n_1325),
.B2(n_1330),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1232),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1238),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1304),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1319),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1249),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1301),
.A2(n_1278),
.B1(n_1216),
.B2(n_1299),
.Y(n_1378)
);

CKINVDCx12_ASAP7_75t_R g1379 ( 
.A(n_1299),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1323),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1278),
.A2(n_1336),
.B1(n_1290),
.B2(n_1307),
.Y(n_1381)
);

BUFx5_ASAP7_75t_L g1382 ( 
.A(n_1288),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1328),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1335),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1204),
.Y(n_1385)
);

INVx8_ASAP7_75t_L g1386 ( 
.A(n_1204),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1336),
.A2(n_1290),
.B1(n_1355),
.B2(n_1351),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1262),
.A2(n_1280),
.B1(n_1239),
.B2(n_1205),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1349),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1212),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1244),
.A2(n_1227),
.B1(n_1298),
.B2(n_1207),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1241),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1245),
.A2(n_1228),
.B1(n_1286),
.B2(n_1202),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1281),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1324),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1293),
.A2(n_1308),
.B1(n_1265),
.B2(n_1240),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1293),
.A2(n_1308),
.B1(n_1265),
.B2(n_1326),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1272),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1348),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1250),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1276),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1201),
.A2(n_1213),
.B1(n_1258),
.B2(n_1269),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1247),
.A2(n_1228),
.B1(n_1271),
.B2(n_1210),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1199),
.A2(n_1345),
.B1(n_1221),
.B2(n_1263),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1333),
.B(n_1343),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1222),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1289),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1277),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1333),
.B(n_1343),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1287),
.A2(n_1259),
.B1(n_1357),
.B2(n_1316),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1231),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1315),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1284),
.Y(n_1414)
);

CKINVDCx11_ASAP7_75t_R g1415 ( 
.A(n_1353),
.Y(n_1415)
);

OAI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1297),
.A2(n_1248),
.B1(n_1350),
.B2(n_1337),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1274),
.A2(n_1275),
.B1(n_1197),
.B2(n_1215),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1285),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1295),
.A2(n_1292),
.B1(n_1339),
.B2(n_1264),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1235),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1217),
.A2(n_1358),
.B1(n_1346),
.B2(n_1334),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1318),
.Y(n_1422)
);

BUFx2_ASAP7_75t_SL g1423 ( 
.A(n_1294),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1255),
.A2(n_1224),
.B1(n_1306),
.B2(n_1305),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1296),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1243),
.A2(n_1230),
.B1(n_1283),
.B2(n_1214),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1352),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1246),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1242),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1260),
.A2(n_1268),
.B1(n_1256),
.B2(n_1267),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1260),
.B(n_1322),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1291),
.A2(n_1273),
.B(n_1229),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1322),
.A2(n_1254),
.B1(n_1208),
.B2(n_1252),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1318),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1257),
.A2(n_1282),
.B1(n_1251),
.B2(n_1206),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1321),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1218),
.A2(n_1225),
.B1(n_1198),
.B2(n_1219),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1321),
.B(n_1253),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1303),
.B(n_1347),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1322),
.A2(n_1261),
.B1(n_1253),
.B2(n_1321),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1312),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1233),
.A2(n_1203),
.B1(n_1211),
.B2(n_1226),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1234),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1233),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1313),
.A2(n_1342),
.B1(n_1340),
.B2(n_1332),
.Y(n_1445)
);

BUFx12f_ASAP7_75t_L g1446 ( 
.A(n_1209),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1261),
.A2(n_1253),
.B1(n_1223),
.B2(n_1220),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1209),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1261),
.A2(n_963),
.B1(n_1320),
.B2(n_1311),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1220),
.A2(n_1327),
.B1(n_963),
.B2(n_1331),
.Y(n_1450)
);

BUFx8_ASAP7_75t_L g1451 ( 
.A(n_1223),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1223),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1220),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1248),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1266),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1300),
.A2(n_963),
.B1(n_1311),
.B2(n_1327),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1200),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1249),
.Y(n_1459)
);

CKINVDCx6p67_ASAP7_75t_R g1460 ( 
.A(n_1317),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1248),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1245),
.B(n_1240),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1300),
.A2(n_1327),
.B1(n_963),
.B2(n_1311),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1349),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1300),
.A2(n_963),
.B1(n_1311),
.B2(n_1327),
.Y(n_1465)
);

BUFx8_ASAP7_75t_L g1466 ( 
.A(n_1249),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1266),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1320),
.A2(n_1311),
.B1(n_963),
.B2(n_1300),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1320),
.A2(n_1311),
.B1(n_963),
.B2(n_1300),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1200),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1349),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1320),
.A2(n_1311),
.B1(n_963),
.B2(n_1300),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1324),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1200),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1310),
.Y(n_1475)
);

CKINVDCx11_ASAP7_75t_R g1476 ( 
.A(n_1310),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1320),
.A2(n_1311),
.B1(n_963),
.B2(n_1300),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1357),
.Y(n_1478)
);

BUFx2_ASAP7_75t_SL g1479 ( 
.A(n_1357),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1200),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1357),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1482)
);

INVx6_ASAP7_75t_L g1483 ( 
.A(n_1236),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1327),
.A2(n_963),
.B1(n_1331),
.B2(n_1311),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1245),
.B(n_1240),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1310),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1320),
.A2(n_963),
.B1(n_1311),
.B2(n_1300),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1300),
.A2(n_1327),
.B1(n_963),
.B2(n_1311),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1349),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1311),
.A2(n_963),
.B1(n_823),
.B2(n_1300),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1357),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1327),
.A2(n_963),
.B1(n_1331),
.B2(n_1311),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1320),
.A2(n_1311),
.B1(n_963),
.B2(n_1300),
.Y(n_1495)
);

BUFx8_ASAP7_75t_SL g1496 ( 
.A(n_1249),
.Y(n_1496)
);

BUFx4f_ASAP7_75t_SL g1497 ( 
.A(n_1249),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1311),
.A2(n_963),
.B1(n_1331),
.B2(n_784),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1427),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1431),
.B(n_1366),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1420),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1456),
.A2(n_1465),
.B1(n_1489),
.B2(n_1463),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1482),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1425),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1395),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1438),
.B(n_1452),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1491),
.A2(n_1493),
.B1(n_1484),
.B2(n_1488),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1366),
.B(n_1449),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1434),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1436),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1399),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1462),
.B(n_1485),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1487),
.B(n_1494),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1435),
.A2(n_1439),
.B(n_1445),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1378),
.B(n_1448),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1378),
.B(n_1362),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1468),
.A2(n_1469),
.B1(n_1495),
.B2(n_1472),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1439),
.A2(n_1445),
.B(n_1437),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1422),
.B(n_1404),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1422),
.B(n_1404),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1443),
.Y(n_1521)
);

INVx6_ASAP7_75t_L g1522 ( 
.A(n_1408),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1424),
.A2(n_1432),
.B(n_1430),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1444),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1440),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1373),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1442),
.A2(n_1426),
.B(n_1421),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1364),
.A2(n_1372),
.B(n_1402),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1371),
.B(n_1416),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1426),
.A2(n_1421),
.B(n_1447),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1428),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1399),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1429),
.B(n_1441),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1389),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_SL g1535 ( 
.A(n_1459),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1446),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1405),
.A2(n_1381),
.B(n_1477),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1451),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1374),
.B(n_1380),
.Y(n_1539)
);

NOR2xp67_ASAP7_75t_R g1540 ( 
.A(n_1365),
.B(n_1486),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1451),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1498),
.A2(n_1493),
.B(n_1484),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1473),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1363),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1359),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1392),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1382),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1391),
.B(n_1450),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1382),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1405),
.A2(n_1381),
.B(n_1387),
.Y(n_1550)
);

INVxp33_ASAP7_75t_L g1551 ( 
.A(n_1471),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1398),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1382),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1382),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1424),
.A2(n_1450),
.B(n_1368),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1473),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1401),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1375),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1453),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1468),
.B(n_1469),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1359),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1376),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1383),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1384),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1472),
.A2(n_1477),
.B(n_1495),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1457),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1417),
.A2(n_1433),
.B(n_1419),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1470),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1474),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1480),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1394),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1423),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1433),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1359),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1417),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1368),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1409),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1455),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1467),
.Y(n_1579)
);

AO31x2_ASAP7_75t_L g1580 ( 
.A1(n_1385),
.A2(n_1410),
.A3(n_1406),
.B(n_1416),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1464),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1379),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1397),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1397),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1360),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1387),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1388),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1393),
.A2(n_1388),
.B(n_1411),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1411),
.Y(n_1589)
);

CKINVDCx11_ASAP7_75t_R g1590 ( 
.A(n_1415),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1396),
.A2(n_1483),
.B(n_1369),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1370),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1361),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1370),
.Y(n_1594)
);

INVx5_ASAP7_75t_L g1595 ( 
.A(n_1483),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1490),
.B(n_1396),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1412),
.Y(n_1597)
);

NAND4xp25_ASAP7_75t_L g1598 ( 
.A(n_1529),
.B(n_1492),
.C(n_1481),
.D(n_1478),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1513),
.B(n_1454),
.Y(n_1599)
);

OAI211xp5_ASAP7_75t_L g1600 ( 
.A1(n_1529),
.A2(n_1414),
.B(n_1476),
.C(n_1461),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1500),
.B(n_1479),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1542),
.A2(n_1567),
.B(n_1518),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1519),
.B(n_1520),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1511),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1506),
.B(n_1367),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1538),
.B(n_1408),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1557),
.B(n_1413),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1590),
.Y(n_1608)
);

CKINVDCx6p67_ASAP7_75t_R g1609 ( 
.A(n_1504),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1519),
.B(n_1408),
.Y(n_1610)
);

INVx4_ASAP7_75t_L g1611 ( 
.A(n_1595),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1502),
.A2(n_1418),
.B1(n_1413),
.B2(n_1403),
.C(n_1475),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1503),
.B(n_1400),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1520),
.B(n_1403),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1551),
.B(n_1390),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1507),
.A2(n_1460),
.B1(n_1497),
.B2(n_1407),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1515),
.B(n_1390),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1507),
.A2(n_1528),
.B(n_1517),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1528),
.A2(n_1386),
.B1(n_1497),
.B2(n_1459),
.C(n_1466),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1541),
.B(n_1536),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1506),
.B(n_1386),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1536),
.B(n_1386),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1568),
.B(n_1377),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1568),
.B(n_1466),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1548),
.B(n_1501),
.Y(n_1626)
);

BUFx12f_ASAP7_75t_L g1627 ( 
.A(n_1593),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1589),
.A2(n_1576),
.B1(n_1596),
.B2(n_1560),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1569),
.B(n_1555),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_SL g1630 ( 
.A1(n_1548),
.A2(n_1572),
.B(n_1589),
.C(n_1525),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1516),
.B(n_1532),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1555),
.B(n_1508),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1516),
.A2(n_1588),
.B(n_1508),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1544),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1556),
.B(n_1577),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1576),
.A2(n_1587),
.B1(n_1582),
.B2(n_1565),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1534),
.B(n_1597),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1577),
.B(n_1539),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1565),
.A2(n_1586),
.B1(n_1587),
.B2(n_1575),
.Y(n_1639)
);

AO22x2_ASAP7_75t_L g1640 ( 
.A1(n_1525),
.A2(n_1584),
.B1(n_1583),
.B2(n_1573),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1555),
.B(n_1524),
.Y(n_1641)
);

AOI22x1_ASAP7_75t_SL g1642 ( 
.A1(n_1559),
.A2(n_1582),
.B1(n_1584),
.B2(n_1583),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1533),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1530),
.A2(n_1527),
.B(n_1514),
.Y(n_1644)
);

OA21x2_ASAP7_75t_L g1645 ( 
.A1(n_1530),
.A2(n_1527),
.B(n_1514),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1588),
.A2(n_1550),
.B(n_1565),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1558),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1596),
.A2(n_1524),
.B1(n_1559),
.B2(n_1504),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1512),
.B(n_1581),
.Y(n_1649)
);

AO32x2_ASAP7_75t_L g1650 ( 
.A1(n_1543),
.A2(n_1573),
.A3(n_1580),
.B1(n_1510),
.B2(n_1509),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1550),
.A2(n_1565),
.B(n_1591),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1531),
.B(n_1586),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_R g1653 ( 
.A(n_1559),
.B(n_1574),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1523),
.A2(n_1572),
.B(n_1504),
.C(n_1543),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1595),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_SL g1656 ( 
.A(n_1523),
.B(n_1595),
.Y(n_1656)
);

OR2x6_ASAP7_75t_L g1657 ( 
.A(n_1518),
.B(n_1591),
.Y(n_1657)
);

NAND2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1595),
.B(n_1559),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1562),
.B(n_1563),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1618),
.A2(n_1537),
.B1(n_1512),
.B2(n_1535),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1603),
.B(n_1523),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1598),
.B(n_1595),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1632),
.B(n_1499),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1611),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1603),
.B(n_1553),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1616),
.A2(n_1537),
.B1(n_1595),
.B2(n_1574),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1658),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1631),
.B(n_1505),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1632),
.B(n_1549),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1600),
.B(n_1505),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1634),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1641),
.B(n_1553),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1643),
.B(n_1533),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1604),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1629),
.B(n_1521),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1629),
.B(n_1521),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1619),
.A2(n_1537),
.B1(n_1594),
.B2(n_1592),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1610),
.B(n_1554),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1647),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1610),
.B(n_1547),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1626),
.B(n_1580),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1636),
.B(n_1564),
.Y(n_1683)
);

AOI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1612),
.A2(n_1540),
.B1(n_1571),
.B2(n_1579),
.C1(n_1578),
.C2(n_1566),
.Y(n_1684)
);

OR2x6_ASAP7_75t_SL g1685 ( 
.A(n_1648),
.B(n_1566),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1640),
.A2(n_1570),
.B1(n_1546),
.B2(n_1526),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1643),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1635),
.B(n_1580),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1614),
.B(n_1638),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1652),
.B(n_1580),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1614),
.B(n_1640),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1660),
.A2(n_1633),
.B(n_1654),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1651),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1650),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1661),
.B(n_1650),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1661),
.B(n_1650),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1672),
.B(n_1650),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1676),
.B(n_1646),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1688),
.B(n_1659),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1660),
.A2(n_1602),
.B1(n_1628),
.B2(n_1640),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1676),
.B(n_1644),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1678),
.A2(n_1639),
.B1(n_1599),
.B2(n_1605),
.C(n_1625),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1680),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1677),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1686),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1663),
.B(n_1659),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1687),
.Y(n_1708)
);

AND2x2_ASAP7_75t_SL g1709 ( 
.A(n_1662),
.B(n_1645),
.Y(n_1709)
);

OAI31xp33_ASAP7_75t_L g1710 ( 
.A1(n_1666),
.A2(n_1630),
.A3(n_1601),
.B(n_1605),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1687),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1678),
.A2(n_1602),
.B(n_1656),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1691),
.B(n_1617),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1684),
.B(n_1637),
.C(n_1613),
.D(n_1649),
.Y(n_1714)
);

INVxp33_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1686),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1664),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1683),
.A2(n_1608),
.B1(n_1642),
.B2(n_1627),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1665),
.B(n_1657),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1716),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1699),
.B(n_1690),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1713),
.B(n_1675),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1703),
.A2(n_1685),
.B1(n_1609),
.B2(n_1658),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1705),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1716),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1720),
.B(n_1673),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1716),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1668),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1720),
.B(n_1673),
.Y(n_1730)
);

BUFx2_ASAP7_75t_SL g1731 ( 
.A(n_1718),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1716),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1705),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1718),
.B(n_1667),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1699),
.B(n_1690),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1689),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1679),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1720),
.B(n_1673),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1696),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1696),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1692),
.B(n_1657),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1699),
.B(n_1682),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1715),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1693),
.B(n_1679),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1719),
.B(n_1710),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1708),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1693),
.B(n_1681),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1696),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1708),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1704),
.Y(n_1752)
);

INVxp33_ASAP7_75t_L g1753 ( 
.A(n_1719),
.Y(n_1753)
);

NOR2x1p5_ASAP7_75t_L g1754 ( 
.A(n_1714),
.B(n_1608),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1698),
.B(n_1687),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1706),
.B(n_1717),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1704),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1756),
.B(n_1706),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1742),
.B(n_1734),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1744),
.B(n_1715),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1746),
.A2(n_1692),
.B1(n_1701),
.B2(n_1710),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1742),
.B(n_1694),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1734),
.B(n_1694),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1755),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1733),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1756),
.B(n_1717),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1725),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1743),
.B(n_1702),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1723),
.B(n_1701),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1733),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1739),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1739),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1740),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1755),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1740),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1721),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1729),
.B(n_1714),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1743),
.B(n_1722),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1734),
.B(n_1694),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1754),
.B(n_1601),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1734),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1745),
.Y(n_1782)
);

NOR2xp67_ASAP7_75t_L g1783 ( 
.A(n_1724),
.B(n_1627),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1727),
.B(n_1698),
.Y(n_1784)
);

INVxp33_ASAP7_75t_L g1785 ( 
.A(n_1753),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1750),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1754),
.A2(n_1703),
.B1(n_1685),
.B2(n_1709),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1750),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1752),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1752),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1757),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1745),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1721),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1722),
.B(n_1735),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1731),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1726),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1726),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1728),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1759),
.B(n_1741),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1759),
.B(n_1741),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1760),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1780),
.Y(n_1804)
);

OAI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1761),
.A2(n_1741),
.B(n_1709),
.Y(n_1805)
);

NAND2x1_ASAP7_75t_L g1806 ( 
.A(n_1781),
.B(n_1741),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1758),
.B(n_1735),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1771),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1763),
.B(n_1779),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1748),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1785),
.B(n_1748),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1763),
.B(n_1741),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1779),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1767),
.B(n_1749),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1781),
.B(n_1731),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1787),
.A2(n_1662),
.B1(n_1712),
.B2(n_1709),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1784),
.B(n_1727),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1769),
.B(n_1749),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1784),
.B(n_1730),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1771),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1758),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

NAND4xp75_ASAP7_75t_L g1823 ( 
.A(n_1783),
.B(n_1709),
.C(n_1624),
.D(n_1623),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1782),
.B(n_1794),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1766),
.B(n_1778),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1772),
.Y(n_1826)
);

OAI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1766),
.A2(n_1684),
.B(n_1682),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1764),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1793),
.B(n_1737),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1797),
.B(n_1730),
.Y(n_1830)
);

OAI211xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1765),
.A2(n_1607),
.B(n_1615),
.C(n_1728),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1778),
.B(n_1620),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1762),
.B(n_1738),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1765),
.B(n_1738),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1773),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1773),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1803),
.B(n_1770),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1821),
.B(n_1770),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1808),
.Y(n_1839)
);

OAI222xp33_ASAP7_75t_L g1840 ( 
.A1(n_1816),
.A2(n_1796),
.B1(n_1764),
.B2(n_1774),
.C1(n_1768),
.C2(n_1762),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1805),
.A2(n_1712),
.B1(n_1653),
.B2(n_1774),
.Y(n_1841)
);

NOR2xp67_ASAP7_75t_SL g1842 ( 
.A(n_1823),
.B(n_1718),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1808),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1811),
.B(n_1796),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1823),
.A2(n_1609),
.B1(n_1697),
.B2(n_1695),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_L g1846 ( 
.A(n_1827),
.B(n_1718),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1810),
.B(n_1695),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1809),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1801),
.A2(n_1623),
.B(n_1624),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1820),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1820),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1822),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1822),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1825),
.B(n_1718),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1826),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1804),
.B(n_1824),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1824),
.B(n_1809),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1831),
.A2(n_1786),
.B1(n_1775),
.B2(n_1790),
.C(n_1788),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1815),
.B(n_1775),
.Y(n_1859)
);

O2A1O1Ixp5_ASAP7_75t_L g1860 ( 
.A1(n_1806),
.A2(n_1791),
.B(n_1788),
.C(n_1789),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1826),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1806),
.A2(n_1768),
.B1(n_1791),
.B2(n_1789),
.C(n_1790),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1839),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1843),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_SL g1865 ( 
.A(n_1860),
.B(n_1825),
.C(n_1815),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1850),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1856),
.B(n_1813),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1851),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1852),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1841),
.A2(n_1857),
.B1(n_1845),
.B2(n_1848),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1848),
.B(n_1813),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1859),
.B(n_1817),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1859),
.Y(n_1873)
);

OAI21xp33_ASAP7_75t_L g1874 ( 
.A1(n_1844),
.A2(n_1846),
.B(n_1837),
.Y(n_1874)
);

AOI21xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1862),
.A2(n_1807),
.B(n_1814),
.Y(n_1875)
);

NAND2x1_ASAP7_75t_L g1876 ( 
.A(n_1842),
.B(n_1801),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1846),
.A2(n_1818),
.B1(n_1812),
.B2(n_1802),
.Y(n_1877)
);

NOR3xp33_ASAP7_75t_SL g1878 ( 
.A(n_1840),
.B(n_1830),
.C(n_1834),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1842),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1838),
.B(n_1817),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1853),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1858),
.A2(n_1828),
.B1(n_1835),
.B2(n_1836),
.C(n_1802),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1867),
.B(n_1849),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1874),
.B(n_1832),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1873),
.B(n_1819),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1871),
.Y(n_1886)
);

OAI211xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1878),
.A2(n_1854),
.B(n_1855),
.C(n_1861),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1872),
.B(n_1819),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1877),
.B(n_1833),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1865),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1876),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1863),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1864),
.B(n_1854),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1865),
.A2(n_1812),
.B1(n_1828),
.B2(n_1712),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1890),
.B(n_1882),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1886),
.B(n_1875),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1886),
.B(n_1880),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1891),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1885),
.Y(n_1899)
);

NAND3xp33_ASAP7_75t_L g1900 ( 
.A(n_1887),
.B(n_1877),
.C(n_1879),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1894),
.B(n_1893),
.Y(n_1901)
);

NAND3xp33_ASAP7_75t_L g1902 ( 
.A(n_1883),
.B(n_1879),
.C(n_1884),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1888),
.B(n_1870),
.Y(n_1903)
);

NOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1893),
.B(n_1866),
.Y(n_1904)
);

OAI22xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1895),
.A2(n_1892),
.B1(n_1881),
.B2(n_1869),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1900),
.A2(n_1889),
.B1(n_1868),
.B2(n_1807),
.C(n_1847),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1902),
.A2(n_1836),
.B1(n_1835),
.B2(n_1833),
.C(n_1792),
.Y(n_1907)
);

AOI211xp5_ASAP7_75t_L g1908 ( 
.A1(n_1896),
.A2(n_1718),
.B(n_1829),
.C(n_1620),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1901),
.A2(n_1792),
.B(n_1776),
.Y(n_1909)
);

NOR3xp33_ASAP7_75t_L g1910 ( 
.A(n_1903),
.B(n_1617),
.C(n_1620),
.Y(n_1910)
);

OAI211xp5_ASAP7_75t_L g1911 ( 
.A1(n_1904),
.A2(n_1718),
.B(n_1799),
.C(n_1798),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1906),
.A2(n_1897),
.B(n_1898),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1910),
.A2(n_1899),
.B1(n_1718),
.B2(n_1606),
.Y(n_1913)
);

AOI21xp33_ASAP7_75t_L g1914 ( 
.A1(n_1905),
.A2(n_1795),
.B(n_1776),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1909),
.A2(n_1907),
.B1(n_1908),
.B2(n_1911),
.C(n_1800),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1905),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1910),
.A2(n_1606),
.B1(n_1712),
.B2(n_1795),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1905),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1916),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1918),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1912),
.B(n_1798),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1913),
.B(n_1799),
.Y(n_1922)
);

XOR2x2_ASAP7_75t_L g1923 ( 
.A(n_1915),
.B(n_1606),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1919),
.A2(n_1914),
.B1(n_1917),
.B2(n_1800),
.C(n_1751),
.Y(n_1924)
);

NAND3x1_ASAP7_75t_L g1925 ( 
.A(n_1921),
.B(n_1708),
.C(n_1732),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_SL g1926 ( 
.A(n_1920),
.B(n_1611),
.C(n_1655),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1925),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1927),
.Y(n_1928)
);

AO22x2_ASAP7_75t_SL g1929 ( 
.A1(n_1928),
.A2(n_1923),
.B1(n_1924),
.B2(n_1926),
.Y(n_1929)
);

NOR2xp67_ASAP7_75t_L g1930 ( 
.A(n_1928),
.B(n_1922),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_1929),
.Y(n_1931)
);

NAND2xp67_ASAP7_75t_L g1932 ( 
.A(n_1930),
.B(n_1621),
.Y(n_1932)
);

OAI21xp33_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1751),
.B(n_1747),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1931),
.B(n_1622),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1934),
.A2(n_1747),
.B(n_1622),
.Y(n_1935)
);

XNOR2xp5_ASAP7_75t_L g1936 ( 
.A(n_1935),
.B(n_1622),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_R g1937 ( 
.A1(n_1936),
.A2(n_1522),
.B1(n_1732),
.B2(n_1711),
.C(n_1712),
.Y(n_1937)
);

AOI211xp5_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1585),
.B(n_1545),
.C(n_1561),
.Y(n_1938)
);


endmodule