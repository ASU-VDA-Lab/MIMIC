module fake_jpeg_166_n_682 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_682);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_682;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_7),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_63),
.Y(n_209)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_11),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_67),
.B(n_73),
.Y(n_151)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_68),
.Y(n_149)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_69),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_70),
.B(n_81),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_78),
.B(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_83),
.B(n_85),
.Y(n_168)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_91),
.B(n_92),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_29),
.B(n_10),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_97),
.B(n_100),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_98),
.Y(n_163)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_48),
.Y(n_102)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_102),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_114),
.Y(n_136)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_36),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_121),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_21),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_120),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_28),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_49),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_125),
.B(n_34),
.Y(n_203)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_28),
.Y(n_128)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_45),
.C(n_49),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_143),
.B(n_59),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_59),
.B1(n_39),
.B2(n_20),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_150),
.A2(n_191),
.B1(n_61),
.B2(n_142),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_38),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_153),
.B(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_165),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_62),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_167),
.B(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_39),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_172),
.B(n_180),
.Y(n_258)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_178),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_120),
.B(n_19),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_103),
.A2(n_37),
.B1(n_56),
.B2(n_54),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_183),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_68),
.B(n_37),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_189),
.B(n_203),
.Y(n_293)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_200),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_107),
.A2(n_20),
.B1(n_31),
.B2(n_54),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_131),
.B(n_34),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_204),
.B(n_213),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_38),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_205),
.B(n_212),
.Y(n_270)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_66),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_116),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_63),
.B(n_33),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_115),
.B(n_41),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_109),
.B(n_33),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_71),
.B(n_41),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_220),
.Y(n_242)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_104),
.Y(n_218)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_122),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_128),
.B(n_19),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_151),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_108),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_88),
.Y(n_247)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_224),
.B(n_243),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_192),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_142),
.A2(n_127),
.B1(n_113),
.B2(n_31),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_227),
.Y(n_361)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_228),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_229),
.A2(n_268),
.B1(n_296),
.B2(n_135),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_230),
.B(n_236),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_123),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_234),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_179),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_181),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_257),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_240),
.A2(n_175),
.B1(n_171),
.B2(n_154),
.Y(n_316)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

INVx4_ASAP7_75t_SL g342 ( 
.A(n_244),
.Y(n_342)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_245),
.Y(n_353)
);

CKINVDCx12_ASAP7_75t_R g246 ( 
.A(n_178),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_246),
.B(n_248),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_156),
.B(n_90),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_158),
.A2(n_64),
.B1(n_76),
.B2(n_75),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_253),
.A2(n_262),
.B1(n_264),
.B2(n_278),
.Y(n_325)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_142),
.Y(n_256)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_176),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_136),
.Y(n_259)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_259),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_132),
.B(n_44),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_283),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_191),
.A2(n_77),
.B1(n_79),
.B2(n_82),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_263),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_150),
.A2(n_98),
.B1(n_89),
.B2(n_129),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_133),
.B(n_124),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_267),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_144),
.B(n_146),
.Y(n_267)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_277),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_185),
.B(n_113),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_271),
.B(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_196),
.Y(n_272)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_183),
.A2(n_25),
.B1(n_56),
.B2(n_53),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_275),
.A2(n_106),
.B(n_112),
.Y(n_339)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_160),
.Y(n_276)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_168),
.B(n_53),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_210),
.A2(n_26),
.B1(n_98),
.B2(n_89),
.Y(n_278)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_137),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_160),
.Y(n_280)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_159),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_286),
.Y(n_331)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_152),
.B(n_0),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

AO22x1_ASAP7_75t_SL g285 ( 
.A1(n_194),
.A2(n_127),
.B1(n_84),
.B2(n_86),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_285),
.B(n_295),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_195),
.B(n_13),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_134),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_290),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_137),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_288),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_139),
.B(n_141),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_138),
.C(n_145),
.Y(n_348)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_148),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_147),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_292),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_140),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_208),
.B(n_0),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_148),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_149),
.B(n_13),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_300),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_186),
.B(n_0),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_209),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_149),
.B(n_13),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_224),
.A2(n_134),
.B1(n_193),
.B2(n_201),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_306),
.A2(n_328),
.B1(n_296),
.B2(n_288),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_224),
.A2(n_264),
.B(n_271),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_308),
.A2(n_282),
.B(n_241),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_316),
.A2(n_285),
.B1(n_234),
.B2(n_272),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_260),
.A2(n_193),
.B1(n_201),
.B2(n_154),
.Y(n_318)
);

OAI22x1_ASAP7_75t_L g403 ( 
.A1(n_318),
.A2(n_344),
.B1(n_351),
.B2(n_135),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_249),
.Y(n_393)
);

AO22x2_ASAP7_75t_SL g323 ( 
.A1(n_262),
.A2(n_171),
.B1(n_177),
.B2(n_184),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_285),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_258),
.A2(n_177),
.B1(n_184),
.B2(n_207),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_299),
.A2(n_207),
.B1(n_211),
.B2(n_219),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_337),
.A2(n_349),
.B1(n_325),
.B2(n_307),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g382 ( 
.A1(n_339),
.A2(n_346),
.B(n_234),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_243),
.B(n_209),
.C(n_211),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_289),
.C(n_255),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_235),
.B(n_169),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_343),
.B(n_358),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_240),
.A2(n_202),
.B1(n_155),
.B2(n_169),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_145),
.B1(n_138),
.B2(n_155),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_219),
.B1(n_173),
.B2(n_187),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_275),
.A2(n_202),
.B1(n_175),
.B2(n_80),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_242),
.A2(n_94),
.B(n_178),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_355),
.A2(n_265),
.B(n_271),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_94),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_363),
.Y(n_415)
);

INVx13_ASAP7_75t_L g364 ( 
.A(n_353),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_364),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_303),
.B(n_257),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_313),
.B(n_239),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_366),
.B(n_367),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_313),
.B(n_270),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_335),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_368),
.B(n_369),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_324),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_283),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_370),
.B(n_375),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_232),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_371),
.B(n_383),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_377),
.B1(n_381),
.B2(n_328),
.Y(n_418)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_374),
.A2(n_391),
.B(n_392),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_238),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_382),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_350),
.A2(n_274),
.B1(n_287),
.B2(n_289),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_360),
.B(n_233),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_334),
.B(n_265),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_387),
.Y(n_436)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_273),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_386),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_334),
.B(n_350),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_269),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_390),
.Y(n_444)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_348),
.C(n_306),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_252),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_308),
.B(n_244),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_338),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_304),
.B(n_226),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_397),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_304),
.B(n_226),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_310),
.B(n_254),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_401),
.Y(n_423)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_399),
.A2(n_400),
.B1(n_403),
.B2(n_404),
.Y(n_435)
);

BUFx12_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_310),
.B(n_284),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_361),
.A2(n_276),
.B1(n_263),
.B2(n_223),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_402),
.A2(n_405),
.B(n_406),
.Y(n_427)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_358),
.B(n_245),
.Y(n_406)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_302),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_407),
.A2(n_354),
.B(n_251),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_297),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_408),
.A2(n_409),
.B(n_357),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_302),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_362),
.B(n_393),
.C(n_370),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_424),
.C(n_428),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_412),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_387),
.A2(n_325),
.B1(n_337),
.B2(n_349),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_417),
.B1(n_425),
.B2(n_431),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_416),
.B(n_445),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_375),
.A2(n_323),
.B1(n_338),
.B2(n_361),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_443),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_339),
.B(n_355),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_422),
.A2(n_374),
.B(n_384),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_362),
.A2(n_323),
.B1(n_346),
.B2(n_332),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_372),
.A2(n_359),
.B1(n_319),
.B2(n_314),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_426),
.A2(n_442),
.B1(n_415),
.B2(n_435),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_314),
.C(n_333),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_376),
.A2(n_359),
.B1(n_231),
.B2(n_290),
.Y(n_431)
);

AO22x1_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_319),
.B1(n_336),
.B2(n_345),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_434),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_381),
.A2(n_231),
.B1(n_279),
.B2(n_280),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_363),
.A2(n_319),
.B1(n_330),
.B2(n_315),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_392),
.A2(n_333),
.B(n_321),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g445 ( 
.A(n_390),
.B(n_345),
.C(n_301),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_395),
.A2(n_352),
.B1(n_347),
.B2(n_330),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_403),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_392),
.A2(n_321),
.B(n_309),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_L g453 ( 
.A1(n_450),
.A2(n_422),
.B(n_410),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_429),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_L g503 ( 
.A(n_452),
.B(n_454),
.C(n_467),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_453),
.A2(n_468),
.B(n_432),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_420),
.B(n_367),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_425),
.B1(n_417),
.B2(n_431),
.Y(n_488)
);

OAI22x1_ASAP7_75t_SL g457 ( 
.A1(n_442),
.A2(n_380),
.B1(n_408),
.B2(n_363),
.Y(n_457)
);

AOI22x1_ASAP7_75t_L g491 ( 
.A1(n_457),
.A2(n_448),
.B1(n_432),
.B2(n_443),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_444),
.B(n_366),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_458),
.B(n_459),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_444),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_462),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_382),
.Y(n_463)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_463),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_383),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_464),
.B(n_482),
.Y(n_506)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_465),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_420),
.B(n_441),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_440),
.A2(n_380),
.B1(n_363),
.B2(n_369),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_469),
.A2(n_460),
.B1(n_463),
.B2(n_468),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_412),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_473),
.Y(n_509)
);

OAI32xp33_ASAP7_75t_L g472 ( 
.A1(n_436),
.A2(n_401),
.A3(n_377),
.B1(n_405),
.B2(n_379),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_472),
.A2(n_450),
.B(n_448),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_428),
.C(n_416),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_479),
.C(n_419),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_423),
.B(n_398),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_477),
.Y(n_514)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_480),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_424),
.B(n_397),
.C(n_394),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_404),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_439),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_484),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_436),
.B(n_399),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_449),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_433),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_446),
.B(n_409),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_486),
.B(n_487),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_446),
.B(n_406),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_488),
.A2(n_489),
.B1(n_491),
.B2(n_498),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_461),
.A2(n_448),
.B1(n_413),
.B2(n_418),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_463),
.A2(n_410),
.B(n_437),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_490),
.A2(n_501),
.B(n_487),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_414),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_493),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_451),
.B(n_414),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_482),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_499),
.C(n_500),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_424),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_495),
.B(n_505),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_467),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_486),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_464),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_502),
.B(n_516),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_504),
.A2(n_511),
.B1(n_515),
.B2(n_462),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_445),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_461),
.A2(n_380),
.B1(n_427),
.B2(n_445),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_507),
.A2(n_510),
.B1(n_457),
.B2(n_460),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_483),
.A2(n_427),
.B1(n_402),
.B2(n_447),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_452),
.A2(n_433),
.B1(n_419),
.B2(n_430),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_322),
.C(n_327),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_466),
.B(n_434),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_513),
.B(n_505),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_454),
.Y(n_516)
);

A2O1A1O1Ixp25_ASAP7_75t_L g519 ( 
.A1(n_477),
.A2(n_407),
.B(n_447),
.C(n_430),
.D(n_301),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_519),
.A2(n_521),
.B(n_465),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_483),
.A2(n_385),
.B(n_354),
.Y(n_521)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_524),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_525),
.A2(n_528),
.B1(n_552),
.B2(n_521),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_489),
.A2(n_483),
.B1(n_476),
.B2(n_484),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_526),
.A2(n_540),
.B1(n_549),
.B2(n_541),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_466),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_527),
.B(n_532),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_485),
.B1(n_456),
.B2(n_471),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_531),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_480),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g560 ( 
.A(n_534),
.B(n_535),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_497),
.B(n_475),
.Y(n_536)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_536),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_478),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_537),
.B(n_518),
.Y(n_563)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_538),
.Y(n_567)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_496),
.Y(n_539)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_488),
.A2(n_458),
.B1(n_470),
.B2(n_473),
.Y(n_540)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_495),
.B(n_455),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_542),
.B(n_546),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_472),
.Y(n_543)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_543),
.Y(n_577)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_496),
.Y(n_544)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_544),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_481),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_545),
.B(n_551),
.Y(n_566)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_520),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_547),
.B(n_548),
.Y(n_580)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_503),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_517),
.A2(n_396),
.B1(n_378),
.B2(n_373),
.Y(n_549)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_510),
.A2(n_352),
.B1(n_342),
.B2(n_309),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_553),
.B(n_554),
.C(n_501),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_513),
.B(n_322),
.C(n_292),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_523),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_555),
.Y(n_568)
);

FAx1_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_491),
.CI(n_490),
.CON(n_558),
.SN(n_558)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_559),
.B(n_562),
.Y(n_603)
);

XNOR2x1_ASAP7_75t_SL g562 ( 
.A(n_535),
.B(n_518),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_527),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_565),
.A2(n_567),
.B1(n_582),
.B2(n_558),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_543),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_569),
.B(n_572),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_533),
.B(n_542),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_SL g600 ( 
.A(n_570),
.B(n_571),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_533),
.B(n_514),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_545),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_530),
.B(n_514),
.C(n_498),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_578),
.C(n_560),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_529),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_400),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_530),
.B(n_491),
.C(n_522),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_581),
.A2(n_536),
.B1(n_554),
.B2(n_532),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_540),
.A2(n_509),
.B1(n_522),
.B2(n_342),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_584),
.A2(n_553),
.B1(n_268),
.B2(n_327),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_SL g617 ( 
.A(n_585),
.B(n_584),
.Y(n_617)
);

AO221x1_ASAP7_75t_L g586 ( 
.A1(n_581),
.A2(n_528),
.B1(n_525),
.B2(n_552),
.C(n_549),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_586),
.B(n_594),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_587),
.B(n_571),
.Y(n_612)
);

AOI321xp33_ASAP7_75t_L g588 ( 
.A1(n_558),
.A2(n_556),
.A3(n_550),
.B1(n_526),
.B2(n_537),
.C(n_509),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g620 ( 
.A1(n_588),
.A2(n_568),
.B(n_583),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_589),
.A2(n_592),
.B1(n_601),
.B2(n_565),
.Y(n_615)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_580),
.Y(n_591)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_591),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_567),
.A2(n_305),
.B1(n_228),
.B2(n_291),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_593),
.A2(n_597),
.B1(n_607),
.B2(n_582),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_305),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_573),
.B(n_237),
.C(n_250),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_596),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_564),
.B(n_259),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_579),
.Y(n_598)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_598),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_573),
.B(n_297),
.C(n_400),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_604),
.C(n_608),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_577),
.A2(n_173),
.B1(n_187),
.B2(n_256),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_559),
.B(n_297),
.C(n_400),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_364),
.Y(n_605)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_605),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_578),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_606),
.B(n_574),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_570),
.B(n_297),
.C(n_197),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_SL g633 ( 
.A(n_610),
.B(n_617),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_612),
.B(n_616),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_560),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_613),
.B(n_627),
.Y(n_644)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_614),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_615),
.A2(n_588),
.B1(n_8),
.B2(n_12),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_603),
.B(n_563),
.C(n_566),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_557),
.C(n_561),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_618),
.B(n_625),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_589),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_619),
.B(n_595),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_620),
.A2(n_602),
.B(n_590),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_583),
.C(n_576),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_585),
.B(n_197),
.C(n_162),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_626),
.B(n_599),
.C(n_600),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_590),
.A2(n_197),
.B1(n_35),
.B2(n_10),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_8),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_628),
.B(n_625),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_629),
.A2(n_645),
.B(n_6),
.Y(n_650)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_631),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_624),
.B(n_601),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_632),
.B(n_638),
.Y(n_649)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_634),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_618),
.A2(n_616),
.B(n_615),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_636),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_609),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_621),
.B(n_593),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_639),
.B(n_643),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_640),
.B(n_641),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_612),
.B(n_604),
.C(n_608),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_642),
.A2(n_622),
.B1(n_628),
.B2(n_613),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_623),
.B(n_8),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_617),
.A2(n_6),
.B(n_16),
.Y(n_645)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_646),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_636),
.B(n_611),
.C(n_626),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_647),
.B(n_648),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_SL g648 ( 
.A1(n_630),
.A2(n_627),
.B(n_611),
.C(n_2),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_650),
.A2(n_657),
.B(n_644),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_630),
.B(n_635),
.C(n_641),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_651),
.B(n_654),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_17),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_653),
.A2(n_14),
.B(n_17),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_637),
.B(n_0),
.C(n_1),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_658),
.A2(n_629),
.B(n_640),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_660),
.A2(n_661),
.B(n_665),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_656),
.A2(n_645),
.B(n_644),
.Y(n_661)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_662),
.Y(n_670)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_663),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_652),
.B(n_633),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_651),
.B(n_649),
.C(n_647),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_666),
.B(n_633),
.Y(n_668)
);

NOR4xp25_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_667),
.C(n_659),
.D(n_648),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_664),
.B(n_655),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_669),
.A2(n_671),
.B(n_648),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_665),
.A2(n_648),
.B(n_654),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_674),
.B(n_675),
.C(n_673),
.Y(n_678)
);

AOI322xp5_ASAP7_75t_L g676 ( 
.A1(n_670),
.A2(n_15),
.A3(n_17),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_2),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_676),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_678),
.A2(n_672),
.B1(n_17),
.B2(n_4),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_679),
.A2(n_677),
.B(n_2),
.Y(n_680)
);

XOR2xp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_2),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_681),
.B(n_3),
.Y(n_682)
);


endmodule