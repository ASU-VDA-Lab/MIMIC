module fake_jpeg_24281_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_10),
.B(n_8),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_3),
.C(n_4),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_14),
.B1(n_15),
.B2(n_24),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_5),
.B1(n_7),
.B2(n_13),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_10),
.B1(n_11),
.B2(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_20),
.Y(n_41)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_35),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_8),
.B1(n_19),
.B2(n_21),
.Y(n_32)
);

OAI32xp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_9),
.A3(n_14),
.B1(n_15),
.B2(n_7),
.Y(n_34)
);

XNOR2x2_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_22),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_40),
.C(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_24),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_34),
.B1(n_26),
.B2(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_35),
.C(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_43),
.C(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_40),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_27),
.A3(n_33),
.B1(n_37),
.B2(n_39),
.C1(n_42),
.C2(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_33),
.Y(n_54)
);


endmodule