module real_aes_7979_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_86), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g449 ( .A(n_0), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_1), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_2), .A2(n_143), .B(n_146), .C(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_3), .A2(n_171), .B(n_172), .Y(n_170) );
INVx1_ASAP7_75t_L g501 ( .A(n_4), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_5), .B(n_182), .Y(n_181) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_6), .A2(n_171), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g143 ( .A(n_7), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g246 ( .A(n_8), .Y(n_246) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_9), .B(n_41), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_10), .A2(n_270), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_11), .B(n_155), .Y(n_223) );
INVx1_ASAP7_75t_L g483 ( .A(n_12), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_13), .B(n_176), .Y(n_534) );
INVx1_ASAP7_75t_L g135 ( .A(n_14), .Y(n_135) );
INVx1_ASAP7_75t_L g546 ( .A(n_15), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_16), .A2(n_190), .B(n_231), .C(n_233), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_17), .B(n_182), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_18), .B(n_472), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_19), .B(n_171), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_20), .B(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_21), .A2(n_176), .B(n_207), .C(n_210), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_22), .B(n_182), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_23), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_24), .A2(n_209), .B(n_233), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_25), .B(n_155), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g137 ( .A(n_26), .Y(n_137) );
INVx1_ASAP7_75t_L g188 ( .A(n_27), .Y(n_188) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_29), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_30), .B(n_155), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_31), .Y(n_452) );
INVx1_ASAP7_75t_L g275 ( .A(n_32), .Y(n_275) );
INVx1_ASAP7_75t_L g491 ( .A(n_33), .Y(n_491) );
INVx2_ASAP7_75t_L g141 ( .A(n_34), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_35), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_36), .A2(n_176), .B(n_177), .C(n_179), .Y(n_175) );
INVxp67_ASAP7_75t_L g276 ( .A(n_37), .Y(n_276) );
CKINVDCx14_ASAP7_75t_R g173 ( .A(n_38), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_39), .A2(n_146), .B(n_187), .C(n_194), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_143), .B(n_146), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_41), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g490 ( .A(n_42), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_43), .A2(n_49), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_43), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_44), .A2(n_62), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_44), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_45), .A2(n_157), .B(n_244), .C(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_46), .B(n_155), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_47), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_48), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_49), .Y(n_443) );
INVx1_ASAP7_75t_L g205 ( .A(n_50), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_51), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_52), .B(n_171), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_53), .A2(n_146), .B1(n_210), .B2(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_54), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_55), .Y(n_498) );
CKINVDCx14_ASAP7_75t_R g242 ( .A(n_56), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_57), .A2(n_179), .B(n_244), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_58), .Y(n_526) );
INVx1_ASAP7_75t_L g480 ( .A(n_59), .Y(n_480) );
INVx1_ASAP7_75t_L g144 ( .A(n_60), .Y(n_144) );
INVx1_ASAP7_75t_L g134 ( .A(n_61), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_62), .Y(n_744) );
INVx1_ASAP7_75t_SL g178 ( .A(n_63), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_65), .B(n_182), .Y(n_212) );
INVx1_ASAP7_75t_L g150 ( .A(n_66), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_67), .A2(n_179), .B(n_472), .C(n_473), .Y(n_471) );
INVxp67_ASAP7_75t_L g474 ( .A(n_68), .Y(n_474) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_70), .A2(n_171), .B(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_71), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_72), .A2(n_171), .B(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_73), .Y(n_494) );
INVx1_ASAP7_75t_L g520 ( .A(n_74), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_75), .A2(n_270), .B(n_271), .Y(n_269) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_76), .Y(n_185) );
INVx1_ASAP7_75t_L g229 ( .A(n_77), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_78), .A2(n_143), .B(n_146), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_79), .A2(n_171), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g232 ( .A(n_80), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_81), .B(n_189), .Y(n_514) );
INVx2_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
INVx1_ASAP7_75t_L g222 ( .A(n_83), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_84), .B(n_472), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_85), .A2(n_143), .B(n_146), .C(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g446 ( .A(n_86), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g458 ( .A(n_86), .Y(n_458) );
OR2x2_ASAP7_75t_L g741 ( .A(n_86), .B(n_448), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_87), .A2(n_146), .B(n_149), .C(n_159), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_88), .B(n_164), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_89), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_90), .A2(n_143), .B(n_146), .C(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_91), .Y(n_538) );
INVx1_ASAP7_75t_L g470 ( .A(n_92), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_93), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_94), .B(n_189), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_95), .A2(n_102), .B1(n_113), .B2(n_754), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_96), .B(n_130), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_97), .B(n_130), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g208 ( .A(n_99), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_100), .A2(n_171), .B(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_105), .Y(n_755) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_453), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g753 ( .A(n_117), .Y(n_753) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_445), .B(n_451), .Y(n_119) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_442), .Y(n_120) );
INVx3_ASAP7_75t_L g742 ( .A(n_121), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_121), .A2(n_456), .B1(n_740), .B2(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_397), .Y(n_121) );
NOR4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_334), .C(n_368), .D(n_384), .Y(n_122) );
NAND4xp25_ASAP7_75t_SL g123 ( .A(n_124), .B(n_260), .C(n_298), .D(n_314), .Y(n_123) );
AOI222xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_197), .B1(n_235), .B2(n_248), .C1(n_253), .C2(n_259), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI31xp33_ASAP7_75t_L g430 ( .A1(n_126), .A2(n_431), .A3(n_432), .B(n_434), .Y(n_430) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_165), .Y(n_126) );
AND2x2_ASAP7_75t_L g405 ( .A(n_127), .B(n_167), .Y(n_405) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_SL g252 ( .A(n_128), .Y(n_252) );
AND2x2_ASAP7_75t_L g259 ( .A(n_128), .B(n_183), .Y(n_259) );
AND2x2_ASAP7_75t_L g319 ( .A(n_128), .B(n_168), .Y(n_319) );
AO21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_161), .Y(n_128) );
INVx3_ASAP7_75t_L g182 ( .A(n_129), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_129), .B(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_129), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_SL g516 ( .A(n_129), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_130), .A2(n_468), .B(n_475), .Y(n_467) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g268 ( .A(n_131), .Y(n_268) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_132), .B(n_133), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_145), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_138), .A2(n_164), .B(n_185), .C(n_186), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_138), .A2(n_219), .B(n_220), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_138), .A2(n_160), .B1(n_488), .B2(n_492), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_138), .A2(n_498), .B(n_499), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_138), .A2(n_520), .B(n_521), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
AND2x4_ASAP7_75t_L g171 ( .A(n_139), .B(n_143), .Y(n_171) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
INVx3_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
INVx1_ASAP7_75t_L g472 ( .A(n_142), .Y(n_472) );
INVx4_ASAP7_75t_SL g160 ( .A(n_143), .Y(n_160) );
BUFx3_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
INVx5_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_154), .C(n_156), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_156), .B(n_222), .C(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_152), .A2(n_153), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g209 ( .A(n_153), .Y(n_209) );
INVx4_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx2_ASAP7_75t_L g244 ( .A(n_155), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_156), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_156), .A2(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g233 ( .A(n_158), .Y(n_233) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_160), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g204 ( .A1(n_160), .A2(n_174), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_SL g228 ( .A1(n_160), .A2(n_174), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_160), .A2(n_174), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_160), .A2(n_174), .B(n_272), .C(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_160), .A2(n_174), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_160), .A2(n_174), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_160), .A2(n_174), .B(n_543), .C(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx1_ASAP7_75t_L g278 ( .A(n_163), .Y(n_278) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_163), .A2(n_530), .B(n_537), .Y(n_529) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_164), .A2(n_240), .B(n_247), .Y(n_239) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_164), .A2(n_541), .B(n_547), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_165), .B(n_349), .Y(n_348) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_166), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_166), .B(n_263), .Y(n_309) );
AND2x2_ASAP7_75t_L g402 ( .A(n_166), .B(n_342), .Y(n_402) );
OAI321xp33_ASAP7_75t_L g436 ( .A1(n_166), .A2(n_252), .A3(n_409), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_166), .B(n_238), .C(n_349), .D(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_183), .Y(n_166) );
AND2x2_ASAP7_75t_L g304 ( .A(n_167), .B(n_250), .Y(n_304) );
AND2x2_ASAP7_75t_L g323 ( .A(n_167), .B(n_252), .Y(n_323) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g251 ( .A(n_168), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g279 ( .A(n_168), .B(n_183), .Y(n_279) );
AND2x2_ASAP7_75t_L g365 ( .A(n_168), .B(n_250), .Y(n_365) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_181), .Y(n_168) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_203), .B(n_212), .Y(n_202) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_169), .A2(n_227), .B(n_234), .Y(n_226) );
BUFx2_ASAP7_75t_L g270 ( .A(n_171), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_176), .B(n_178), .Y(n_177) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_180), .Y(n_535) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_182), .A2(n_478), .B(n_484), .Y(n_477) );
INVx3_ASAP7_75t_SL g250 ( .A(n_183), .Y(n_250) );
AND2x2_ASAP7_75t_L g297 ( .A(n_183), .B(n_284), .Y(n_297) );
OR2x2_ASAP7_75t_L g330 ( .A(n_183), .B(n_252), .Y(n_330) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_183), .Y(n_337) );
AND2x2_ASAP7_75t_L g366 ( .A(n_183), .B(n_251), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_183), .B(n_339), .Y(n_381) );
AND2x2_ASAP7_75t_L g413 ( .A(n_183), .B(n_405), .Y(n_413) );
AND2x2_ASAP7_75t_L g422 ( .A(n_183), .B(n_264), .Y(n_422) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_195), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .C(n_192), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g274 ( .A1(n_189), .A2(n_209), .B1(n_275), .B2(n_276), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_189), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
INVx5_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_190), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_190), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_190), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_193), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
INVx1_ASAP7_75t_SL g390 ( .A(n_199), .Y(n_390) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g255 ( .A(n_200), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g237 ( .A(n_201), .B(n_215), .Y(n_237) );
AND2x2_ASAP7_75t_L g326 ( .A(n_201), .B(n_239), .Y(n_326) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g296 ( .A(n_202), .B(n_226), .Y(n_296) );
OR2x2_ASAP7_75t_L g307 ( .A(n_202), .B(n_239), .Y(n_307) );
AND2x2_ASAP7_75t_L g333 ( .A(n_202), .B(n_239), .Y(n_333) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_202), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_209), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_209), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g503 ( .A(n_210), .Y(n_503) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_213), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_213), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g306 ( .A(n_214), .B(n_307), .Y(n_306) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_214), .A2(n_296), .A3(n_302), .B1(n_333), .B2(n_383), .C1(n_393), .C2(n_395), .Y(n_392) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_215), .B(n_238), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_215), .B(n_239), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_215), .B(n_256), .Y(n_313) );
AND2x2_ASAP7_75t_L g367 ( .A(n_215), .B(n_333), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_215), .Y(n_371) );
AND2x2_ASAP7_75t_L g383 ( .A(n_215), .B(n_226), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_215), .B(n_255), .Y(n_415) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g280 ( .A(n_216), .B(n_226), .Y(n_280) );
BUFx3_ASAP7_75t_L g294 ( .A(n_216), .Y(n_294) );
AND3x2_ASAP7_75t_L g376 ( .A(n_216), .B(n_356), .C(n_377), .Y(n_376) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_217), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_217), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_217), .B(n_538), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g236 ( .A(n_226), .B(n_237), .C(n_238), .Y(n_236) );
INVx1_ASAP7_75t_SL g256 ( .A(n_226), .Y(n_256) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_226), .Y(n_361) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g355 ( .A(n_237), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g362 ( .A(n_237), .Y(n_362) );
AND2x2_ASAP7_75t_L g400 ( .A(n_238), .B(n_378), .Y(n_400) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx3_ASAP7_75t_L g281 ( .A(n_239), .Y(n_281) );
AND2x2_ASAP7_75t_L g356 ( .A(n_239), .B(n_256), .Y(n_356) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OR2x2_ASAP7_75t_L g300 ( .A(n_250), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g419 ( .A(n_250), .B(n_319), .Y(n_419) );
AND2x2_ASAP7_75t_L g433 ( .A(n_250), .B(n_252), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_251), .B(n_264), .Y(n_374) );
AND2x2_ASAP7_75t_L g421 ( .A(n_251), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g284 ( .A(n_252), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_264), .Y(n_301) );
INVx1_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
AND2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_264), .Y(n_342) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_254), .A2(n_385), .B1(n_389), .B2(n_391), .C(n_392), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_255), .B(n_257), .Y(n_254) );
AND2x2_ASAP7_75t_L g288 ( .A(n_255), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_258), .B(n_295), .Y(n_438) );
AOI322xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_280), .A3(n_281), .B1(n_282), .B2(n_288), .C1(n_290), .C2(n_297), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_279), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_263), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_263), .B(n_329), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_263), .A2(n_279), .B(n_353), .C(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_263), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_263), .B(n_323), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_263), .B(n_405), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_263), .B(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_264), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_264), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g394 ( .A(n_264), .B(n_281), .Y(n_394) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_269), .B(n_277), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_266), .A2(n_286), .B(n_287), .Y(n_285) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_266), .A2(n_519), .B(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AOI21xp5_ASAP7_75t_SL g510 ( .A1(n_267), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_268), .A2(n_487), .B(n_493), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_268), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_268), .A2(n_497), .B(n_504), .Y(n_496) );
INVx1_ASAP7_75t_L g286 ( .A(n_269), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_277), .Y(n_287) );
INVx1_ASAP7_75t_L g369 ( .A(n_279), .Y(n_369) );
OAI31xp33_ASAP7_75t_L g379 ( .A1(n_279), .A2(n_304), .A3(n_380), .B(n_382), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_279), .B(n_285), .Y(n_431) );
INVx1_ASAP7_75t_SL g292 ( .A(n_280), .Y(n_292) );
AND2x2_ASAP7_75t_L g325 ( .A(n_280), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g406 ( .A(n_280), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g291 ( .A(n_281), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
AND2x2_ASAP7_75t_L g343 ( .A(n_281), .B(n_296), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_281), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g435 ( .A(n_281), .B(n_383), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_283), .B(n_353), .Y(n_426) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g340 ( .A(n_285), .Y(n_340) );
NAND2xp33_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
OAI211xp5_ASAP7_75t_SL g334 ( .A1(n_292), .A2(n_335), .B(n_341), .C(n_357), .Y(n_334) );
OR2x2_ASAP7_75t_L g409 ( .A(n_292), .B(n_390), .Y(n_409) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_294), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_294), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g315 ( .A(n_296), .B(n_316), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B(n_305), .C(n_308), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g349 ( .A(n_301), .Y(n_349) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_304), .B(n_342), .Y(n_347) );
INVx1_ASAP7_75t_L g353 ( .A(n_304), .Y(n_353) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g312 ( .A(n_307), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g345 ( .A(n_307), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g407 ( .A(n_307), .Y(n_407) );
AOI21xp33_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_310), .B(n_312), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_310), .A2(n_321), .B(n_324), .Y(n_320) );
AOI211xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_320), .C(n_327), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_315), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_318), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g331 ( .A(n_319), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g386 ( .A1(n_321), .A2(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_326), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g351 ( .A(n_326), .Y(n_351) );
AOI21xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_331), .B(n_332), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g382 ( .A(n_333), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_339), .B(n_365), .Y(n_391) );
AND2x2_ASAP7_75t_L g404 ( .A(n_339), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g418 ( .A(n_339), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g428 ( .A(n_339), .B(n_366), .Y(n_428) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_344), .C(n_352), .Y(n_341) );
INVx1_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_348), .B2(n_350), .Y(n_344) );
OR2x2_ASAP7_75t_L g350 ( .A(n_346), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_346), .B(n_407), .Y(n_429) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g423 ( .A(n_356), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_363), .B1(n_366), .B2(n_367), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g441 ( .A(n_361), .Y(n_441) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g387 ( .A(n_365), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B(n_372), .C(n_379), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_387), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR5xp2_ASAP7_75t_L g397 ( .A(n_398), .B(n_416), .C(n_424), .D(n_430), .E(n_436), .Y(n_397) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_401), .B(n_403), .C(n_410), .Y(n_398) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B(n_408), .Y(n_403) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_413), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_423), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g439 ( .A(n_419), .Y(n_439) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B(n_429), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_446), .B(n_452), .Y(n_451) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_447), .B(n_458), .Y(n_750) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g457 ( .A(n_448), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_451), .A2(n_454), .B(n_752), .Y(n_453) );
OAI222xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_743), .B1(n_746), .B2(n_748), .C1(n_749), .C2(n_751), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_459), .B1(n_740), .B2(n_742), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g747 ( .A(n_459), .Y(n_747) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND4x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_658), .C(n_705), .D(n_725), .Y(n_460) );
NOR3xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_588), .C(n_613), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_506), .B(n_548), .C(n_578), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_485), .Y(n_464) );
INVx3_ASAP7_75t_SL g630 ( .A(n_465), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_465), .B(n_561), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_465), .B(n_495), .Y(n_711) );
AND2x2_ASAP7_75t_L g734 ( .A(n_465), .B(n_600), .Y(n_734) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g552 ( .A(n_467), .B(n_477), .Y(n_552) );
INVx3_ASAP7_75t_L g565 ( .A(n_467), .Y(n_565) );
AND2x2_ASAP7_75t_L g570 ( .A(n_467), .B(n_476), .Y(n_570) );
OR2x2_ASAP7_75t_L g621 ( .A(n_467), .B(n_562), .Y(n_621) );
BUFx2_ASAP7_75t_L g641 ( .A(n_467), .Y(n_641) );
AND2x2_ASAP7_75t_L g651 ( .A(n_467), .B(n_562), .Y(n_651) );
AND2x2_ASAP7_75t_L g657 ( .A(n_467), .B(n_486), .Y(n_657) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_477), .B(n_562), .Y(n_576) );
INVx2_ASAP7_75t_L g586 ( .A(n_477), .Y(n_586) );
AND2x2_ASAP7_75t_L g599 ( .A(n_477), .B(n_565), .Y(n_599) );
OR2x2_ASAP7_75t_L g610 ( .A(n_477), .B(n_562), .Y(n_610) );
AND2x2_ASAP7_75t_SL g656 ( .A(n_477), .B(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g668 ( .A(n_477), .Y(n_668) );
AND2x2_ASAP7_75t_L g714 ( .A(n_477), .B(n_486), .Y(n_714) );
INVx3_ASAP7_75t_SL g587 ( .A(n_485), .Y(n_587) );
OR2x2_ASAP7_75t_L g640 ( .A(n_485), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
INVx3_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
AND2x2_ASAP7_75t_L g629 ( .A(n_486), .B(n_496), .Y(n_629) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_486), .Y(n_697) );
AOI33xp33_ASAP7_75t_L g701 ( .A1(n_486), .A2(n_630), .A3(n_637), .B1(n_646), .B2(n_702), .B3(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g550 ( .A(n_495), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_495), .B(n_565), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_495), .B(n_625), .C(n_627), .Y(n_624) );
AND2x2_ASAP7_75t_L g650 ( .A(n_495), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_495), .B(n_657), .Y(n_660) );
AND2x2_ASAP7_75t_L g713 ( .A(n_495), .B(n_714), .Y(n_713) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g569 ( .A(n_496), .Y(n_569) );
OR2x2_ASAP7_75t_L g663 ( .A(n_496), .B(n_562), .Y(n_663) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_527), .Y(n_506) );
AOI32xp33_ASAP7_75t_L g614 ( .A1(n_507), .A2(n_615), .A3(n_617), .B1(n_619), .B2(n_622), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g687 ( .A(n_507), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g717 ( .A(n_507), .Y(n_717) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g649 ( .A(n_508), .B(n_633), .Y(n_649) );
AND2x2_ASAP7_75t_L g669 ( .A(n_508), .B(n_595), .Y(n_669) );
AND2x2_ASAP7_75t_L g737 ( .A(n_508), .B(n_655), .Y(n_737) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
INVx3_ASAP7_75t_L g558 ( .A(n_509), .Y(n_558) );
AND2x2_ASAP7_75t_L g572 ( .A(n_509), .B(n_556), .Y(n_572) );
OR2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_555), .Y(n_577) );
INVx1_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
AND2x2_ASAP7_75t_L g592 ( .A(n_509), .B(n_566), .Y(n_592) );
AND2x2_ASAP7_75t_L g594 ( .A(n_509), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_509), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g647 ( .A(n_509), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_509), .B(n_732), .Y(n_731) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx2_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
AND2x2_ASAP7_75t_L g602 ( .A(n_518), .B(n_528), .Y(n_602) );
AND2x2_ASAP7_75t_L g612 ( .A(n_518), .B(n_540), .Y(n_612) );
INVx2_ASAP7_75t_L g732 ( .A(n_527), .Y(n_732) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_528), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
AND2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g633 ( .A(n_528), .B(n_596), .Y(n_633) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g581 ( .A(n_529), .Y(n_581) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g646 ( .A(n_529), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_529), .B(n_556), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g557 ( .A(n_539), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_539), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g655 ( .A(n_539), .Y(n_655) );
INVx1_ASAP7_75t_L g688 ( .A(n_539), .Y(n_688) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g566 ( .A(n_540), .B(n_556), .Y(n_566) );
INVx1_ASAP7_75t_L g596 ( .A(n_540), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_553), .B1(n_559), .B2(n_566), .C(n_567), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_550), .B(n_570), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_550), .B(n_633), .Y(n_710) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_552), .B(n_600), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_552), .B(n_561), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_552), .B(n_575), .Y(n_704) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
AND2x2_ASAP7_75t_L g601 ( .A(n_557), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g679 ( .A(n_557), .Y(n_679) );
AND2x2_ASAP7_75t_L g611 ( .A(n_558), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_558), .B(n_581), .Y(n_627) );
AND2x2_ASAP7_75t_L g691 ( .A(n_558), .B(n_617), .Y(n_691) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g600 ( .A(n_562), .B(n_569), .Y(n_600) );
AND2x2_ASAP7_75t_L g696 ( .A(n_563), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_565), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_566), .B(n_573), .Y(n_661) );
AND2x2_ASAP7_75t_L g681 ( .A(n_566), .B(n_581), .Y(n_681) );
AND2x2_ASAP7_75t_L g702 ( .A(n_566), .B(n_646), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .A3(n_573), .B1(n_574), .B2(n_577), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_SL g575 ( .A(n_569), .Y(n_575) );
NAND2x1_ASAP7_75t_L g616 ( .A(n_569), .B(n_599), .Y(n_616) );
OR2x2_ASAP7_75t_L g620 ( .A(n_569), .B(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_569), .B(n_668), .Y(n_721) );
INVx1_ASAP7_75t_L g589 ( .A(n_570), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g707 ( .A1(n_571), .A2(n_662), .B1(n_708), .B2(n_711), .C(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g579 ( .A(n_572), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g622 ( .A(n_572), .B(n_595), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_572), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g700 ( .A(n_572), .B(n_633), .Y(n_700) );
INVxp67_ASAP7_75t_L g636 ( .A(n_573), .Y(n_636) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g706 ( .A(n_575), .B(n_693), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_575), .B(n_656), .Y(n_729) );
INVx1_ASAP7_75t_L g604 ( .A(n_577), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_577), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g722 ( .A(n_577), .B(n_723), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_582), .B(n_585), .Y(n_578) );
AND2x2_ASAP7_75t_L g591 ( .A(n_580), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g675 ( .A(n_584), .B(n_595), .Y(n_675) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AND2x2_ASAP7_75t_L g693 ( .A(n_586), .B(n_651), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_586), .B(n_650), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_587), .B(n_599), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_593), .C(n_603), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_624), .B1(n_628), .B2(n_631), .C(n_634), .Y(n_623) );
AOI31xp33_ASAP7_75t_L g718 ( .A1(n_589), .A2(n_719), .A3(n_720), .B(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B1(n_599), .B2(n_601), .Y(n_593) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g719 ( .A(n_599), .Y(n_719) );
INVx1_ASAP7_75t_L g682 ( .A(n_600), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g725 ( .A1(n_602), .A2(n_726), .B(n_728), .C(n_730), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_607), .B2(n_611), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_608), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_610), .A2(n_644), .B1(n_663), .B2(n_699), .C(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g694 ( .A(n_611), .Y(n_694) );
INVx1_ASAP7_75t_L g648 ( .A(n_612), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_614), .B(n_623), .C(n_638), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_615), .A2(n_665), .B(n_669), .Y(n_664) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_617), .B(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g724 ( .A(n_618), .Y(n_724) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g662 ( .A(n_625), .B(n_645), .Y(n_662) );
INVx1_ASAP7_75t_L g637 ( .A(n_626), .Y(n_637) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g635 ( .A(n_629), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_629), .B(n_667), .Y(n_666) );
NOR4xp25_ASAP7_75t_L g634 ( .A(n_630), .B(n_635), .C(n_636), .D(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_643), .B1(n_649), .B2(n_650), .C1(n_652), .C2(n_656), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g736 ( .A(n_640), .Y(n_736) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_652), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_657), .A2(n_713), .B(n_715), .Y(n_712) );
NOR4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_670), .C(n_683), .D(n_698), .Y(n_658) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .C(n_664), .Y(n_659) );
INVx1_ASAP7_75t_L g739 ( .A(n_660), .Y(n_739) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_667), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
OAI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_676), .B2(n_677), .C1(n_680), .C2(n_682), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_675), .A2(n_706), .B(n_707), .C(n_718), .Y(n_705) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OAI222xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_689), .B1(n_690), .B2(n_692), .C1(n_694), .C2(n_695), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_700), .A2(n_703), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI211xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_733), .B(n_735), .C(n_738), .Y(n_730) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g748 ( .A(n_743), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
endmodule