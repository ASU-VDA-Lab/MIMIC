module fake_jpeg_19923_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_9),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_SL g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_78),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_73),
.B(n_59),
.C(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_61),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_73),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_67),
.B(n_48),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_101),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_0),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_64),
.B1(n_66),
.B2(n_50),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_114),
.B1(n_116),
.B2(n_119),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_68),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_123),
.C(n_1),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_57),
.B1(n_68),
.B2(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_45),
.B1(n_49),
.B2(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_121),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_55),
.B1(n_69),
.B2(n_56),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_74),
.B1(n_62),
.B2(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_60),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_75),
.C(n_65),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_136),
.B1(n_132),
.B2(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_130),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_113),
.C(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_1),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_2),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_3),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_28),
.B(n_7),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_6),
.B1(n_10),
.B2(n_16),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_136),
.C(n_23),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_149),
.B1(n_17),
.B2(n_25),
.Y(n_152)
);

AO21x2_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_43),
.B(n_24),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_151),
.C(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_149),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_142),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_146),
.B(n_138),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_30),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_32),
.Y(n_164)
);


endmodule