module real_aes_2290_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_796, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_796;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g227 ( .A(n_0), .B(n_149), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_1), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_2), .B(n_155), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_3), .B(n_145), .Y(n_504) );
INVx1_ASAP7_75t_L g142 ( .A(n_4), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_5), .B(n_155), .Y(n_168) );
NAND2xp33_ASAP7_75t_SL g219 ( .A(n_6), .B(n_153), .Y(n_219) );
INVx1_ASAP7_75t_L g200 ( .A(n_7), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_8), .A2(n_42), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_8), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g791 ( .A(n_9), .Y(n_791) );
AND2x2_ASAP7_75t_L g166 ( .A(n_10), .B(n_159), .Y(n_166) );
AND2x2_ASAP7_75t_L g506 ( .A(n_11), .B(n_193), .Y(n_506) );
AND2x2_ASAP7_75t_L g514 ( .A(n_12), .B(n_216), .Y(n_514) );
INVx2_ASAP7_75t_L g160 ( .A(n_13), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_14), .B(n_145), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_15), .Y(n_114) );
AND3x1_ASAP7_75t_L g788 ( .A(n_15), .B(n_36), .C(n_789), .Y(n_788) );
AOI221x1_ASAP7_75t_L g213 ( .A1(n_16), .A2(n_137), .B1(n_214), .B2(n_216), .C(n_218), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_17), .B(n_155), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_18), .B(n_155), .Y(n_487) );
INVx1_ASAP7_75t_L g118 ( .A(n_19), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_20), .A2(n_90), .B1(n_155), .B2(n_201), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_21), .A2(n_137), .B(n_170), .Y(n_169) );
AOI221xp5_ASAP7_75t_SL g180 ( .A1(n_22), .A2(n_37), .B1(n_137), .B2(n_155), .C(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_23), .B(n_149), .Y(n_171) );
AOI22xp5_ASAP7_75t_SL g779 ( .A1(n_24), .A2(n_78), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_24), .Y(n_781) );
OR2x2_ASAP7_75t_L g161 ( .A(n_25), .B(n_89), .Y(n_161) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_25), .A2(n_89), .B(n_160), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_26), .B(n_145), .Y(n_192) );
INVxp67_ASAP7_75t_L g212 ( .A(n_27), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_28), .Y(n_120) );
AND2x2_ASAP7_75t_L g243 ( .A(n_29), .B(n_158), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_30), .A2(n_137), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_31), .A2(n_216), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_32), .B(n_145), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_33), .A2(n_137), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_34), .B(n_145), .Y(n_473) );
AND2x2_ASAP7_75t_L g138 ( .A(n_35), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g153 ( .A(n_35), .B(n_142), .Y(n_153) );
INVx1_ASAP7_75t_L g208 ( .A(n_35), .Y(n_208) );
OR2x6_ASAP7_75t_L g116 ( .A(n_36), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_38), .B(n_155), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_39), .A2(n_82), .B1(n_137), .B2(n_206), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_40), .B(n_145), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_41), .B(n_155), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_42), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_43), .B(n_149), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_44), .A2(n_137), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g230 ( .A(n_45), .B(n_158), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_46), .B(n_149), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_47), .B(n_158), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_48), .B(n_155), .Y(n_462) );
INVx1_ASAP7_75t_L g141 ( .A(n_49), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_49), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_50), .B(n_145), .Y(n_512) );
AND2x2_ASAP7_75t_L g478 ( .A(n_51), .B(n_158), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_52), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_53), .B(n_155), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_54), .B(n_149), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_55), .B(n_149), .Y(n_472) );
AND2x2_ASAP7_75t_L g162 ( .A(n_56), .B(n_158), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_57), .B(n_155), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_58), .B(n_145), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_59), .B(n_155), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_60), .A2(n_137), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_61), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_62), .B(n_159), .Y(n_195) );
AND2x2_ASAP7_75t_L g493 ( .A(n_63), .B(n_159), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_64), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_65), .A2(n_137), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_66), .B(n_145), .Y(n_172) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_67), .B(n_193), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_68), .B(n_149), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_69), .B(n_149), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_70), .A2(n_93), .B1(n_137), .B2(n_206), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_71), .B(n_145), .Y(n_490) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_73), .B(n_149), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_74), .A2(n_137), .B(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_75), .A2(n_137), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_76), .A2(n_137), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g475 ( .A(n_77), .B(n_159), .Y(n_475) );
INVx1_ASAP7_75t_L g780 ( .A(n_78), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_79), .B(n_158), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_80), .B(n_155), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_81), .A2(n_84), .B1(n_155), .B2(n_201), .Y(n_278) );
INVx1_ASAP7_75t_L g119 ( .A(n_83), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_85), .B(n_149), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_86), .B(n_149), .Y(n_183) );
AND2x2_ASAP7_75t_L g544 ( .A(n_87), .B(n_193), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_88), .A2(n_137), .B(n_143), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_91), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_92), .A2(n_137), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_94), .B(n_145), .Y(n_542) );
INVxp67_ASAP7_75t_L g215 ( .A(n_95), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_96), .B(n_155), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_97), .B(n_145), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_98), .A2(n_137), .B(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g492 ( .A(n_99), .Y(n_492) );
BUFx2_ASAP7_75t_L g106 ( .A(n_100), .Y(n_106) );
BUFx2_ASAP7_75t_SL g771 ( .A(n_100), .Y(n_771) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_782), .B(n_792), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_121), .B(n_769), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp33_ASAP7_75t_SL g772 ( .A1(n_108), .A2(n_773), .B(n_776), .Y(n_772) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_120), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g775 ( .A(n_113), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x6_ASAP7_75t_SL g453 ( .A(n_114), .B(n_116), .Y(n_453) );
OR2x6_ASAP7_75t_SL g754 ( .A(n_114), .B(n_115), .Y(n_754) );
OR2x2_ASAP7_75t_L g768 ( .A(n_114), .B(n_116), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g787 ( .A(n_117), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AO221x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_755), .B2(n_763), .C(n_764), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_122), .Y(n_763) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_452), .B1(n_454), .B2(n_754), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_126), .B(n_761), .Y(n_760) );
AOI22x1_ASAP7_75t_L g776 ( .A1(n_126), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
INVx4_ASAP7_75t_L g777 ( .A(n_126), .Y(n_777) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_391), .Y(n_126) );
NOR3xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_284), .C(n_335), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_174), .B(n_231), .C(n_262), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_133), .B(n_236), .Y(n_399) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g244 ( .A(n_134), .B(n_165), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_134), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g261 ( .A(n_134), .B(n_251), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_134), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g298 ( .A(n_134), .B(n_274), .Y(n_298) );
INVx2_ASAP7_75t_L g324 ( .A(n_134), .Y(n_324) );
AND2x4_ASAP7_75t_L g333 ( .A(n_134), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g438 ( .A(n_134), .B(n_305), .Y(n_438) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_157), .B(n_162), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_154), .Y(n_135) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
BUFx3_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
AND2x6_ASAP7_75t_L g149 ( .A(n_139), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
AND2x4_ASAP7_75t_L g206 ( .A(n_140), .B(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x4_ASAP7_75t_L g145 ( .A(n_141), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B(n_152), .Y(n_143) );
AND2x4_ASAP7_75t_L g156 ( .A(n_146), .B(n_150), .Y(n_156) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_149), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_152), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_152), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_152), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_152), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_152), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_152), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_152), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_152), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_152), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_152), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_152), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_152), .A2(n_542), .B(n_543), .Y(n_541) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g155 ( .A(n_153), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g220 ( .A(n_156), .Y(n_220) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_157), .A2(n_237), .B(n_243), .Y(n_236) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_157), .A2(n_237), .B(n_243), .Y(n_251) );
AOI21x1_ASAP7_75t_L g499 ( .A1(n_157), .A2(n_500), .B(n_506), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_158), .Y(n_157) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_158), .A2(n_180), .B(n_184), .Y(n_179) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_158), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_158), .A2(n_539), .B(n_540), .Y(n_538) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x4_ASAP7_75t_L g173 ( .A(n_160), .B(n_161), .Y(n_173) );
AND2x2_ASAP7_75t_L g322 ( .A(n_163), .B(n_323), .Y(n_322) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_163), .A2(n_327), .A3(n_331), .B1(n_338), .B2(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_163), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g259 ( .A(n_164), .B(n_260), .Y(n_259) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_164), .B(n_254), .C(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g358 ( .A(n_164), .B(n_261), .Y(n_358) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_165), .Y(n_248) );
INVx5_ASAP7_75t_L g283 ( .A(n_165), .Y(n_283) );
AND2x4_ASAP7_75t_L g339 ( .A(n_165), .B(n_251), .Y(n_339) );
OR2x2_ASAP7_75t_L g354 ( .A(n_165), .B(n_274), .Y(n_354) );
OR2x2_ASAP7_75t_L g380 ( .A(n_165), .B(n_236), .Y(n_380) );
AND2x2_ASAP7_75t_L g388 ( .A(n_165), .B(n_334), .Y(n_388) );
AND2x4_ASAP7_75t_SL g413 ( .A(n_165), .B(n_333), .Y(n_413) );
OR2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_173), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_173), .B(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_173), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_173), .B(n_215), .Y(n_214) );
NOR3xp33_ASAP7_75t_L g218 ( .A(n_173), .B(n_219), .C(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_173), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_173), .A2(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_175), .B(n_333), .Y(n_409) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_185), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_176), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR2x6_ASAP7_75t_SL g233 ( .A(n_177), .B(n_234), .Y(n_233) );
INVxp67_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g258 ( .A(n_178), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_178), .B(n_293), .Y(n_311) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_178), .Y(n_449) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
AND2x2_ASAP7_75t_L g291 ( .A(n_179), .B(n_222), .Y(n_291) );
INVx2_ASAP7_75t_L g319 ( .A(n_179), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_179), .B(n_186), .Y(n_360) );
BUFx3_ASAP7_75t_L g384 ( .A(n_179), .Y(n_384) );
OR2x2_ASAP7_75t_L g396 ( .A(n_179), .B(n_186), .Y(n_396) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_179), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_185), .A2(n_427), .B1(n_430), .B2(n_431), .Y(n_426) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_196), .Y(n_185) );
INVx1_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
OR2x2_ASAP7_75t_L g265 ( .A(n_186), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g272 ( .A(n_186), .Y(n_272) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_186), .B(n_197), .Y(n_289) );
AND2x4_ASAP7_75t_L g294 ( .A(n_186), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g303 ( .A(n_186), .Y(n_303) );
OR2x2_ASAP7_75t_L g309 ( .A(n_186), .B(n_197), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_186), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_186), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_186), .B(n_291), .Y(n_425) );
OR2x2_ASAP7_75t_L g441 ( .A(n_186), .B(n_344), .Y(n_441) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_195), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_193), .Y(n_187) );
INVx2_ASAP7_75t_SL g276 ( .A(n_193), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_193), .A2(n_487), .B(n_488), .Y(n_486) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g217 ( .A(n_194), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_196), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_196), .B(n_258), .Y(n_374) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_221), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_197), .B(n_222), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_197), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_197), .B(n_266), .Y(n_270) );
INVx3_ASAP7_75t_L g295 ( .A(n_197), .Y(n_295) );
INVx1_ASAP7_75t_L g328 ( .A(n_197), .Y(n_328) );
AND2x2_ASAP7_75t_L g408 ( .A(n_197), .B(n_272), .Y(n_408) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_213), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_201), .B1(n_206), .B2(n_211), .Y(n_198) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_205), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2x1p5_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g468 ( .A(n_216), .Y(n_468) );
INVx4_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AOI21x1_ASAP7_75t_L g223 ( .A1(n_217), .A2(n_224), .B(n_230), .Y(n_223) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_217), .A2(n_508), .B(n_514), .Y(n_507) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_222), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
AND2x2_ASAP7_75t_L g318 ( .A(n_222), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g344 ( .A(n_222), .B(n_266), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_222), .B(n_295), .Y(n_361) );
INVx1_ASAP7_75t_L g367 ( .A(n_222), .Y(n_367) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
AOI222xp33_ASAP7_75t_SL g231 ( .A1(n_232), .A2(n_235), .B1(n_245), .B2(n_252), .C1(n_255), .C2(n_259), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_244), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_236), .B(n_305), .Y(n_356) );
AND2x4_ASAP7_75t_L g372 ( .A(n_236), .B(n_283), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g297 ( .A(n_248), .B(n_298), .Y(n_297) );
AOI222xp33_ASAP7_75t_L g262 ( .A1(n_249), .A2(n_263), .B1(n_268), .B2(n_273), .C1(n_281), .C2(n_796), .Y(n_262) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g401 ( .A(n_250), .B(n_305), .Y(n_401) );
OR2x2_ASAP7_75t_L g444 ( .A(n_250), .B(n_350), .Y(n_444) );
AND2x2_ASAP7_75t_L g273 ( .A(n_251), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g334 ( .A(n_251), .Y(n_334) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_251), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g362 ( .A1(n_252), .A2(n_363), .B(n_368), .C(n_369), .Y(n_362) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g390 ( .A(n_254), .Y(n_390) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
AND2x2_ASAP7_75t_L g304 ( .A(n_260), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g313 ( .A(n_260), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI31xp33_ASAP7_75t_L g355 ( .A1(n_263), .A2(n_281), .A3(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_264), .A2(n_314), .B(n_358), .C(n_359), .Y(n_357) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
OR2x2_ASAP7_75t_L g346 ( .A(n_265), .B(n_295), .Y(n_346) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
BUFx2_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
AND2x2_ASAP7_75t_L g323 ( .A(n_274), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_275), .Y(n_305) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .B(n_280), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_283), .B(n_340), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_296), .B(n_299), .C(n_321), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_292), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_318), .Y(n_325) );
OR2x2_ASAP7_75t_L g301 ( .A(n_290), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g331 ( .A(n_290), .B(n_305), .Y(n_331) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g407 ( .A(n_291), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g430 ( .A(n_292), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_294), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_294), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g442 ( .A(n_294), .B(n_318), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_294), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g385 ( .A(n_295), .B(n_367), .Y(n_385) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AOI322xp5_ASAP7_75t_L g439 ( .A1(n_298), .A2(n_318), .A3(n_372), .B1(n_397), .B2(n_440), .C1(n_442), .C2(n_443), .Y(n_439) );
AOI211xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_304), .B(n_306), .C(n_315), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_302), .B(n_330), .Y(n_352) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g317 ( .A(n_303), .B(n_318), .Y(n_317) );
NOR2x1p5_ASAP7_75t_L g383 ( .A(n_303), .B(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_303), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_304), .A2(n_322), .B(n_325), .C(n_326), .Y(n_321) );
AND2x4_ASAP7_75t_L g340 ( .A(n_305), .B(n_324), .Y(n_340) );
INVx2_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_305), .B(n_339), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_305), .B(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_305), .B(n_429), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_305), .B(n_333), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B(n_312), .Y(n_306) );
AND2x2_ASAP7_75t_L g402 ( .A(n_308), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g330 ( .A(n_311), .Y(n_330) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_320), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_323), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g417 ( .A(n_323), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_329), .B(n_331), .C(n_332), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_330), .Y(n_414) );
INVx3_ASAP7_75t_SL g429 ( .A(n_333), .Y(n_429) );
NAND5xp2_ASAP7_75t_L g335 ( .A(n_336), .B(n_355), .C(n_362), .D(n_375), .E(n_386), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B1(n_345), .B2(n_347), .C1(n_351), .C2(n_353), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_338), .A2(n_419), .B1(n_423), .B2(n_424), .Y(n_418) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g368 ( .A(n_339), .B(n_340), .Y(n_368) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_349), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_350), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g387 ( .A(n_350), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g398 ( .A(n_350), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g428 ( .A(n_354), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g376 ( .A(n_361), .Y(n_376) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_373), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_372), .A2(n_376), .B1(n_377), .B2(n_381), .Y(n_375) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g389 ( .A(n_374), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g394 ( .A(n_376), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_SL g422 ( .A(n_385), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_410), .C(n_433), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_409), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B1(n_400), .B2(n_402), .C(n_405), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g434 ( .A(n_396), .B(n_422), .Y(n_434) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OAI321xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .A3(n_415), .B1(n_417), .B2(n_418), .C(n_426), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_424), .A2(n_446), .B1(n_450), .B2(n_451), .Y(n_445) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B(n_439), .C(n_445), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
CKINVDCx11_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_453), .Y(n_762) );
INVx4_ASAP7_75t_L g759 ( .A(n_454), .Y(n_759) );
AND3x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_632), .C(n_728), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_574), .C(n_601), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_494), .B(n_523), .C(n_547), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_476), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_458), .A2(n_525), .B(n_529), .C(n_535), .Y(n_524) );
OR2x2_ASAP7_75t_L g647 ( .A(n_458), .B(n_584), .Y(n_647) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g614 ( .A(n_459), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_459), .B(n_585), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_459), .B(n_730), .Y(n_745) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
AND2x2_ASAP7_75t_L g531 ( .A(n_460), .B(n_477), .Y(n_531) );
INVx1_ASAP7_75t_L g551 ( .A(n_460), .Y(n_551) );
OR2x2_ASAP7_75t_L g566 ( .A(n_460), .B(n_485), .Y(n_566) );
INVx2_ASAP7_75t_L g572 ( .A(n_460), .Y(n_572) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_460), .Y(n_627) );
INVx1_ASAP7_75t_L g704 ( .A(n_460), .Y(n_704) );
NOR2x1_ASAP7_75t_SL g553 ( .A(n_467), .B(n_485), .Y(n_553) );
AND2x2_ASAP7_75t_L g583 ( .A(n_467), .B(n_572), .Y(n_583) );
AO21x1_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_469), .B(n_475), .Y(n_467) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_468), .A2(n_469), .B(n_475), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
OR2x2_ASAP7_75t_L g577 ( .A(n_476), .B(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_476), .B(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g705 ( .A(n_476), .Y(n_705) );
NAND2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
OR2x2_ASAP7_75t_SL g565 ( .A(n_477), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g569 ( .A(n_477), .Y(n_569) );
INVx4_ASAP7_75t_L g585 ( .A(n_477), .Y(n_585) );
OR2x2_ASAP7_75t_L g600 ( .A(n_477), .B(n_533), .Y(n_600) );
AND2x2_ASAP7_75t_L g639 ( .A(n_477), .B(n_553), .Y(n_639) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_477), .Y(n_651) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g532 ( .A(n_485), .B(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g584 ( .A(n_485), .B(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g599 ( .A(n_485), .Y(n_599) );
AND2x2_ASAP7_75t_L g615 ( .A(n_485), .B(n_585), .Y(n_615) );
AND2x2_ASAP7_75t_L g628 ( .A(n_485), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g660 ( .A(n_485), .B(n_572), .Y(n_660) );
INVx2_ASAP7_75t_SL g730 ( .A(n_485), .Y(n_730) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NOR2xp67_ASAP7_75t_L g495 ( .A(n_496), .B(n_515), .Y(n_495) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_496), .A2(n_602), .B(n_606), .C(n_622), .Y(n_601) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g697 ( .A(n_497), .B(n_536), .Y(n_697) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx2_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
AND2x4_ASAP7_75t_SL g557 ( .A(n_498), .B(n_537), .Y(n_557) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_498), .Y(n_561) );
AND2x2_ASAP7_75t_L g619 ( .A(n_498), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g693 ( .A(n_498), .Y(n_693) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_499), .Y(n_595) );
AND2x2_ASAP7_75t_L g638 ( .A(n_499), .B(n_507), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
INVx2_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
AND2x2_ASAP7_75t_L g588 ( .A(n_507), .B(n_537), .Y(n_588) );
INVx2_ASAP7_75t_L g620 ( .A(n_507), .Y(n_620) );
OR2x2_ASAP7_75t_L g643 ( .A(n_507), .B(n_518), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_513), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_515), .B(n_560), .Y(n_667) );
AND2x2_ASAP7_75t_L g701 ( .A(n_515), .B(n_637), .Y(n_701) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI31xp33_ASAP7_75t_SL g622 ( .A1(n_516), .A2(n_603), .A3(n_623), .B(n_630), .Y(n_622) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_517), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx3_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
AND2x2_ASAP7_75t_L g573 ( .A(n_518), .B(n_536), .Y(n_573) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
AND2x4_ASAP7_75t_L g563 ( .A(n_519), .B(n_520), .Y(n_563) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g708 ( .A(n_526), .Y(n_708) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_528), .B(n_537), .Y(n_590) );
AND2x2_ASAP7_75t_L g631 ( .A(n_528), .B(n_546), .Y(n_631) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g611 ( .A(n_532), .B(n_569), .Y(n_611) );
AND2x2_ASAP7_75t_L g570 ( .A(n_533), .B(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_533), .Y(n_579) );
INVx2_ASAP7_75t_L g629 ( .A(n_533), .Y(n_629) );
AND2x2_ASAP7_75t_L g719 ( .A(n_533), .B(n_704), .Y(n_719) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g725 ( .A(n_535), .Y(n_725) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_536), .B(n_545), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_536), .B(n_595), .Y(n_664) );
AND2x2_ASAP7_75t_L g712 ( .A(n_536), .B(n_638), .Y(n_712) );
INVx4_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g621 ( .A(n_537), .B(n_593), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_537), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g642 ( .A(n_537), .Y(n_642) );
BUFx2_ASAP7_75t_L g658 ( .A(n_537), .Y(n_658) );
AND2x4_ASAP7_75t_L g692 ( .A(n_537), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g737 ( .A(n_537), .B(n_638), .Y(n_737) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_544), .Y(n_537) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AOI222xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_554), .B1(n_558), .B2(n_564), .C1(n_567), .C2(n_573), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_549), .A2(n_613), .B1(n_616), .B2(n_621), .Y(n_612) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g596 ( .A(n_550), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_550), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_550), .B(n_615), .Y(n_748) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g709 ( .A(n_551), .B(n_615), .Y(n_709) );
OR2x2_ASAP7_75t_L g686 ( .A(n_552), .B(n_568), .Y(n_686) );
OR2x2_ASAP7_75t_L g694 ( .A(n_552), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g678 ( .A(n_553), .B(n_571), .Y(n_678) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OR2x2_ASAP7_75t_L g586 ( .A(n_556), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g736 ( .A(n_556), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g687 ( .A(n_557), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_557), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g722 ( .A(n_557), .Y(n_722) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx2_ASAP7_75t_L g707 ( .A(n_560), .Y(n_707) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g609 ( .A(n_561), .B(n_588), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_562), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_562), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g711 ( .A(n_562), .B(n_583), .Y(n_711) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g645 ( .A(n_563), .B(n_631), .Y(n_645) );
AND2x2_ASAP7_75t_L g688 ( .A(n_563), .B(n_620), .Y(n_688) );
AND2x4_ASAP7_75t_L g603 ( .A(n_564), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g744 ( .A(n_566), .B(n_600), .Y(n_744) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_568), .B(n_583), .Y(n_727) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_569), .B(n_583), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_569), .A2(n_610), .B(n_711), .C(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g741 ( .A(n_569), .B(n_719), .Y(n_741) );
INVx1_ASAP7_75t_L g652 ( .A(n_570), .Y(n_652) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_573), .B(n_637), .Y(n_636) );
OAI21xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_586), .B(n_589), .Y(n_574) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_577), .A2(n_730), .B1(n_731), .B2(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g605 ( .A(n_579), .Y(n_605) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_585), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g677 ( .A(n_585), .Y(n_677) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_596), .Y(n_589) );
INVx1_ASAP7_75t_L g668 ( .A(n_590), .Y(n_668) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_610), .B(n_612), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g653 ( .A(n_608), .B(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g690 ( .A(n_608), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_608), .B(n_638), .Y(n_726) );
INVx1_ASAP7_75t_L g746 ( .A(n_609), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_611), .A2(n_714), .B1(n_717), .B2(n_720), .C(n_723), .Y(n_713) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI321xp33_ASAP7_75t_L g734 ( .A1(n_616), .A2(n_651), .A3(n_735), .B1(n_738), .B2(n_740), .C(n_742), .Y(n_734) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g675 ( .A(n_620), .Y(n_675) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g669 ( .A(n_625), .Y(n_669) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g695 ( .A(n_626), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_628), .A2(n_656), .B1(n_660), .B2(n_661), .C(n_666), .Y(n_655) );
INVxp67_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
INVx1_ASAP7_75t_L g654 ( .A(n_631), .Y(n_654) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_633), .B(n_679), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_655), .C(n_670), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_639), .B1(n_640), .B2(n_646), .C(n_648), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g753 ( .A(n_638), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_644), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_642), .B(n_688), .Y(n_733) );
INVx2_ASAP7_75t_SL g665 ( .A(n_643), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_644), .A2(n_649), .B1(n_650), .B2(n_653), .Y(n_648) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_652), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_653), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g659 ( .A(n_654), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_656), .A2(n_699), .B1(n_701), .B2(n_702), .C1(n_706), .C2(n_709), .Y(n_698) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_657), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g732 ( .A(n_657), .B(n_711), .Y(n_732) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_665), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_665), .B(n_725), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B(n_669), .Y(n_666) );
NAND2xp33_ASAP7_75t_SL g670 ( .A(n_671), .B(n_676), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_676), .B(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g679 ( .A(n_680), .B(n_698), .C(n_710), .D(n_713), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B(n_687), .C(n_689), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_686), .A2(n_690), .B1(n_694), .B2(n_696), .Y(n_689) );
INVx1_ASAP7_75t_L g716 ( .A(n_688), .Y(n_716) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_705), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_722), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_726), .B(n_727), .Y(n_723) );
NOR4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_734), .C(n_747), .D(n_749), .Y(n_728) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
CKINVDCx11_ASAP7_75t_R g758 ( .A(n_754), .Y(n_758) );
OAI21x1_ASAP7_75t_SL g755 ( .A1(n_756), .A2(n_759), .B(n_760), .Y(n_755) );
BUFx4f_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
INVxp33_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g794 ( .A(n_785), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_SL g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
endmodule