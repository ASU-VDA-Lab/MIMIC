module fake_jpeg_27265_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_46),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_31),
.B1(n_20),
.B2(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_35),
.B1(n_23),
.B2(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_17),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_30),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_65),
.A2(n_71),
.B(n_77),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_84),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_31),
.B1(n_20),
.B2(n_29),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_35),
.B1(n_42),
.B2(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_75),
.B1(n_81),
.B2(n_51),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_20),
.B1(n_29),
.B2(n_34),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_40),
.C(n_43),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_90),
.C(n_28),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_35),
.B1(n_42),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_86),
.B1(n_91),
.B2(n_51),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_40),
.B1(n_35),
.B2(n_42),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_28),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_21),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_32),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_36),
.B1(n_43),
.B2(n_24),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_92),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_98),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_30),
.B(n_54),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_113),
.B1(n_85),
.B2(n_66),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_105),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_112),
.B1(n_67),
.B2(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_50),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_36),
.B1(n_50),
.B2(n_43),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_50),
.B1(n_43),
.B2(n_28),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_93),
.B(n_80),
.C(n_90),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_32),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_83),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_65),
.B(n_87),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_120),
.A2(n_138),
.B(n_102),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_124),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_67),
.B1(n_76),
.B2(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_127),
.B1(n_143),
.B2(n_103),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_94),
.B(n_118),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_92),
.B1(n_66),
.B2(n_88),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_134),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_89),
.C(n_59),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_115),
.C(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_139),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_142),
.B1(n_113),
.B2(n_95),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_30),
.B1(n_32),
.B2(n_28),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_145),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_72),
.B1(n_59),
.B2(n_33),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_100),
.A2(n_33),
.B1(n_59),
.B2(n_4),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_2),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_107),
.B(n_98),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_151),
.B(n_153),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_170),
.C(n_171),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_123),
.B(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_169),
.B1(n_175),
.B2(n_2),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_168),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_114),
.B(n_117),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_133),
.B1(n_120),
.B2(n_124),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_126),
.C(n_129),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_106),
.C(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_119),
.C(n_94),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_135),
.C(n_33),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

AO22x2_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_102),
.B1(n_140),
.B2(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_179),
.B1(n_196),
.B2(n_153),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_135),
.B1(n_138),
.B2(n_33),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_197),
.C(n_198),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_185),
.B(n_190),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_188)
);

AO21x1_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_175),
.B(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_158),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_152),
.A2(n_163),
.B1(n_150),
.B2(n_154),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_3),
.C(n_5),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_3),
.C(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_204),
.Y(n_222)
);

OAI322xp33_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_172),
.A3(n_159),
.B1(n_166),
.B2(n_165),
.C1(n_162),
.C2(n_160),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_SL g220 ( 
.A(n_201),
.B(n_178),
.C(n_203),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_151),
.C(n_171),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_211),
.C(n_212),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_210),
.B1(n_217),
.B2(n_178),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_173),
.C(n_154),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_159),
.C(n_164),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_155),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_189),
.B1(n_180),
.B2(n_195),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_156),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_5),
.C(n_6),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_213),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_226),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_217),
.B1(n_206),
.B2(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_195),
.B1(n_179),
.B2(n_193),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_233),
.B1(n_216),
.B2(n_205),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_183),
.B1(n_188),
.B2(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_206),
.B1(n_199),
.B2(n_211),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_182),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_7),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_186),
.B(n_197),
.C(n_7),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_236),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_208),
.C(n_199),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_233),
.C(n_9),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_8),
.C(n_9),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_8),
.C(n_9),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_220),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_247),
.B(n_8),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_219),
.B(n_223),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_253),
.B(n_10),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_224),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_238),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_226),
.B(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_255),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_244),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_257),
.B(n_259),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_245),
.C(n_248),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_262),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_245),
.C(n_224),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_11),
.B(n_12),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_264),
.A2(n_11),
.B(n_13),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_13),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_260),
.B(n_15),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_13),
.B(n_16),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.Y(n_271)
);


endmodule