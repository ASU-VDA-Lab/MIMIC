module real_jpeg_17324_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_0),
.B(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_1),
.A2(n_55),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_1),
.A2(n_56),
.B1(n_423),
.B2(n_427),
.Y(n_422)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_2),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_74),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_4),
.A2(n_74),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_4),
.A2(n_74),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_26),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_5),
.A2(n_71),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_5),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_71),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_5),
.B(n_147),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_5),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_5),
.B(n_250),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_6),
.Y(n_172)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_15),
.B(n_17),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_8),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_8),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

BUFx4f_ASAP7_75t_L g329 ( 
.A(n_11),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_12),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_12),
.A2(n_29),
.B1(n_325),
.B2(n_330),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_12),
.A2(n_29),
.B1(n_218),
.B2(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_12),
.A2(n_29),
.B1(n_432),
.B2(n_434),
.Y(n_431)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_58),
.B(n_470),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_19),
.B(n_49),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_21),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_30),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_31),
.A2(n_41),
.B1(n_69),
.B2(n_72),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g333 ( 
.A1(n_31),
.A2(n_41),
.B1(n_69),
.B2(n_72),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_41),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_32),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_41),
.A2(n_51),
.B(n_458),
.Y(n_457)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_42),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_42),
.Y(n_194)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_42),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_43),
.Y(n_134)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_49),
.B(n_463),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_49),
.B(n_463),
.Y(n_469)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_50),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_54),
.A2(n_55),
.B1(n_339),
.B2(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_57),
.B(n_71),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_412),
.B(n_464),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

AO221x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_311),
.B1(n_405),
.B2(n_410),
.C(n_411),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_241),
.B(n_310),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_204),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_63),
.B(n_204),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_148),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_64),
.B(n_149),
.C(n_182),
.Y(n_401)
);

XOR2x1_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_65),
.A2(n_66),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_65),
.B(n_439),
.C(n_440),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_65),
.B(n_417),
.C(n_438),
.Y(n_453)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_66),
.B(n_351),
.C(n_356),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_66),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_67),
.A2(n_68),
.B1(n_357),
.B2(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_67),
.B(n_79),
.C(n_104),
.Y(n_399)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_69),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_71),
.B(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_104),
.B2(n_105),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_98),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_80),
.A2(n_89),
.B1(n_98),
.B2(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_80),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_80),
.B(n_89),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_87),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_84),
.Y(n_234)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_88),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_89),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_89),
.A2(n_337),
.B(n_346),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_92),
.Y(n_287)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_96),
.Y(n_269)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_98),
.Y(n_248)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_104),
.A2(n_105),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_104),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_104),
.A2(n_105),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_129),
.B1(n_141),
.B2(n_147),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_106),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_106),
.A2(n_129),
.B(n_147),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_106),
.A2(n_147),
.B1(n_422),
.B2(n_431),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_106),
.A2(n_129),
.B1(n_147),
.B2(n_422),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_122),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B1(n_117),
.B2(n_121),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_122),
.B(n_152),
.Y(n_456)
);

OA22x2_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g263 ( 
.A(n_124),
.Y(n_263)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_124),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_131),
.Y(n_435)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_135),
.A2(n_222),
.A3(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_221)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_140),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_140),
.Y(n_433)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_182),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.C(n_156),
.Y(n_149)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_150),
.B(n_364),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_150),
.A2(n_212),
.B1(n_333),
.B2(n_334),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_154),
.A2(n_156),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_156),
.B(n_278),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_161),
.B(n_169),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_170),
.B1(n_176),
.B2(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_165),
.Y(n_330)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_169),
.A2(n_317),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_170),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g355 ( 
.A(n_172),
.Y(n_355)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_178),
.Y(n_271)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_198),
.B2(n_199),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_184),
.B(n_198),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_195),
.B2(n_197),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_198),
.A2(n_199),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_199),
.B(n_289),
.Y(n_290)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_213),
.C(n_220),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_205),
.A2(n_206),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_210),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_210),
.B(n_259),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_211),
.B(n_333),
.C(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21x1_ASAP7_75t_L g362 ( 
.A1(n_212),
.A2(n_363),
.B(n_368),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_254),
.C(n_255),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_213),
.A2(n_255),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_213),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_213),
.A2(n_220),
.B1(n_297),
.B2(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_213),
.A2(n_297),
.B1(n_316),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_SL g348 ( 
.A(n_237),
.B(n_324),
.Y(n_348)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_240),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_301),
.B(n_309),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_256),
.B(n_300),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_253),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_247),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_246),
.A2(n_247),
.B1(n_353),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_R g293 ( 
.A(n_247),
.B(n_261),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_247),
.B(n_353),
.Y(n_352)
);

AO22x2_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_248),
.B(n_249),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_249),
.A2(n_250),
.B1(n_338),
.B2(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_303),
.C(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_292),
.B(n_299),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_276),
.B(n_291),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_264),
.A3(n_268),
.B1(n_270),
.B2(n_272),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_275),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_288),
.B(n_290),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_283),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_305),
.Y(n_309)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_375),
.C(n_388),
.Y(n_311)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_312),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_358),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_313),
.B(n_358),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_335),
.C(n_350),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_335),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_332),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_333),
.C(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_323),
.B1(n_324),
.B2(n_331),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_333),
.A2(n_334),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_333),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_348),
.B1(n_372),
.B2(n_374),
.Y(n_371)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_348),
.A2(n_370),
.B(n_372),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_387),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_369),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_362),
.B(n_369),
.C(n_451),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_365),
.B(n_437),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_368),
.B(n_442),
.C(n_444),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_368),
.B(n_442),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_373),
.B(n_459),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_406),
.B(n_407),
.C(n_409),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_386),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_386),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_382),
.C(n_384),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_379),
.B1(n_382),
.B2(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_391),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_400),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_393),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.C(n_398),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_396),
.A2(n_398),
.B1(n_399),
.B2(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_396),
.Y(n_404)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_402),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_452),
.C(n_462),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_446),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_414),
.A2(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_441),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_415),
.B(n_441),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_438),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_436),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_436),
.C(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_431),
.B(n_456),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_436),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_436),
.B(n_440),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_444),
.A2(n_445),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_450),
.Y(n_466)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_448),
.Y(n_449)
);

A2O1A1O1Ixp25_ASAP7_75t_L g464 ( 
.A1(n_452),
.A2(n_462),
.B(n_465),
.C(n_468),
.D(n_469),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_454),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_454),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_457),
.CI(n_460),
.CON(n_454),
.SN(n_454)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_457),
.C(n_460),
.Y(n_463)
);


endmodule