module real_jpeg_2037_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_2),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_33),
.B1(n_41),
.B2(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_3),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_41),
.C(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_52),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_28),
.C(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_3),
.B(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_21),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_22),
.C(n_25),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_36),
.Y(n_147)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_99)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_107),
.B1(n_165),
.B2(n_166),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_106),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_84),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_15),
.B(n_84),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_65),
.C(n_75),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_16),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_50),
.B2(n_64),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_34),
.B1(n_35),
.B2(n_49),
.Y(n_18)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_35),
.C(n_64),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_31),
.B(n_32),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_20),
.A2(n_31),
.B1(n_32),
.B2(n_99),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_20),
.A2(n_31),
.B1(n_32),
.B2(n_99),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_25),
.B(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22x1_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_28),
.B(n_140),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_34),
.A2(n_35),
.B1(n_97),
.B2(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_35),
.B(n_97),
.C(n_156),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B(n_45),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_40),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_44),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_41),
.B(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_53),
.B(n_56),
.C(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_61),
.B1(n_62),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_56),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_75),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_74),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_74),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_68),
.A2(n_69),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_117),
.C(n_147),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_80),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_92),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_80),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_132),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_83),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_93),
.B2(n_94),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_104),
.B2(n_105),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_98),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_126),
.B(n_164),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_111),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_118),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_138),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_117),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_118),
.B1(n_148),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_158),
.B(n_163),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_152),
.B(n_157),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_143),
.B(n_151),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_137),
.B(n_142),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B(n_136),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_150),
.Y(n_151)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_162),
.Y(n_163)
);


endmodule