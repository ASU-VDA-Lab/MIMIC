module fake_jpeg_1369_n_99 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_33),
.B1(n_35),
.B2(n_27),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_47),
.B1(n_6),
.B2(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_33),
.B1(n_28),
.B2(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_5),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_54),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_42),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_58),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_6),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_43),
.B1(n_46),
.B2(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_56),
.B1(n_15),
.B2(n_19),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_46),
.B1(n_16),
.B2(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_10),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_73),
.B1(n_67),
.B2(n_65),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_56),
.C(n_26),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_77),
.C(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_78),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_73),
.C2(n_23),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_11),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_81),
.C(n_61),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_59),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_71),
.B(n_62),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_81),
.C(n_83),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_92),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_88),
.C(n_85),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_90),
.B(n_80),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_12),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_13),
.Y(n_99)
);


endmodule