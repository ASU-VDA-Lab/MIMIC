module fake_jpeg_10244_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_41),
.Y(n_77)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_46),
.Y(n_59)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_60),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_26),
.B1(n_28),
.B2(n_19),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_23),
.B1(n_33),
.B2(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_47),
.B1(n_36),
.B2(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_65),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_29),
.B1(n_20),
.B2(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_89),
.Y(n_144)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_88),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_48),
.B1(n_29),
.B2(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_87),
.A2(n_27),
.B1(n_22),
.B2(n_44),
.Y(n_137)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_94),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_41),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_96),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_30),
.B1(n_27),
.B2(n_32),
.Y(n_120)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_37),
.C(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_100),
.Y(n_145)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_99),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_107),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_104),
.Y(n_125)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_68),
.Y(n_105)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_19),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_37),
.C(n_39),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_16),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_115),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_64),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_116),
.B1(n_39),
.B2(n_44),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_62),
.B(n_30),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_11),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_49),
.B(n_34),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_120),
.A2(n_121),
.B1(n_101),
.B2(n_78),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_44),
.B1(n_34),
.B2(n_32),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_141),
.B1(n_110),
.B2(n_116),
.Y(n_180)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_132),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_91),
.B(n_17),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_80),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_138),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_81),
.B1(n_94),
.B2(n_84),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_22),
.B1(n_24),
.B2(n_35),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_34),
.B1(n_35),
.B2(n_24),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_89),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_91),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_159),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_176),
.B1(n_180),
.B2(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_160),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_125),
.B(n_137),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_157),
.B(n_143),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_108),
.B(n_96),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_165),
.B(n_166),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_100),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_164),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_115),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_168),
.C(n_126),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_83),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_79),
.C(n_82),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_101),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_90),
.B1(n_88),
.B2(n_95),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_174),
.B1(n_118),
.B2(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_92),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_134),
.B(n_105),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_173),
.B(n_35),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_117),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_127),
.A2(n_106),
.B1(n_86),
.B2(n_111),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_17),
.B(n_34),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_124),
.B(n_17),
.Y(n_202)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_118),
.B1(n_139),
.B2(n_126),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_78),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_164),
.B1(n_150),
.B2(n_31),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_153),
.B1(n_174),
.B2(n_178),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_120),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_197),
.C(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_125),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_202),
.B(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_9),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_124),
.C(n_136),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_210),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_154),
.B1(n_177),
.B2(n_165),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_214),
.B1(n_15),
.B2(n_7),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_149),
.B(n_148),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_130),
.B(n_123),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_135),
.C(n_24),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_31),
.B(n_1),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_155),
.B1(n_152),
.B2(n_151),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_173),
.B(n_160),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_241),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_205),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_188),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_224),
.B1(n_233),
.B2(n_234),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_9),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_182),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_236),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_0),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_2),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_10),
.C(n_12),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_200),
.C(n_201),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_249),
.C(n_250),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_205),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_245),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_206),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_209),
.C(n_187),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_246),
.B(n_252),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_188),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_254),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_189),
.C(n_210),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_189),
.C(n_190),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_223),
.B(n_202),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_213),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_190),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_191),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_220),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_195),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_269),
.B1(n_278),
.B2(n_281),
.Y(n_286)
);

NAND2x1_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_239),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_271),
.B(n_215),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_192),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_203),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_243),
.A2(n_219),
.B1(n_215),
.B2(n_217),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_240),
.B1(n_252),
.B2(n_238),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_253),
.B(n_220),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_217),
.C(n_222),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_277),
.C(n_255),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_221),
.C(n_236),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_221),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_282),
.B1(n_199),
.B2(n_10),
.Y(n_295)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_208),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_292),
.C(n_3),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_246),
.B(n_254),
.C(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_245),
.B(n_233),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_5),
.B(n_11),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_296),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_260),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_280),
.B(n_265),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_276),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_275),
.B1(n_283),
.B2(n_274),
.Y(n_302)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

AOI221xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_10),
.B1(n_12),
.B2(n_5),
.C(n_8),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_302),
.A2(n_300),
.B1(n_289),
.B2(n_285),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_280),
.B(n_5),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_311),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_11),
.C(n_15),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_3),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_294),
.B1(n_286),
.B2(n_287),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_318),
.B1(n_299),
.B2(n_4),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_319),
.C(n_312),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_284),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_299),
.Y(n_326)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_284),
.B1(n_288),
.B2(n_291),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_317),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_324),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

AOI221xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_293),
.B1(n_306),
.B2(n_304),
.C(n_308),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_313),
.B(n_320),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_319),
.C(n_314),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_330),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_333),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_327),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_4),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_4),
.Y(n_337)
);


endmodule