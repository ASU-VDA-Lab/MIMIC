module fake_jpeg_17498_n_358 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_41),
.B(n_66),
.Y(n_114)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_SL g96 ( 
.A(n_43),
.Y(n_96)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_47),
.B(n_1),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_57),
.Y(n_69)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_63),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2x1_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_31),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_71),
.A2(n_87),
.B(n_68),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_31),
.B1(n_36),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_85),
.B1(n_97),
.B2(n_111),
.Y(n_125)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_22),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_101),
.Y(n_138)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_37),
.B1(n_18),
.B2(n_29),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_83),
.A2(n_103),
.B1(n_112),
.B2(n_117),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_36),
.B1(n_33),
.B2(n_30),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_18),
.B(n_35),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_44),
.B1(n_50),
.B2(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_27),
.B1(n_35),
.B2(n_25),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_100),
.A2(n_11),
.B1(n_12),
.B2(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_26),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_62),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_40),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_116),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_42),
.A2(n_24),
.B1(n_22),
.B2(n_30),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_24),
.B1(n_22),
.B2(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_1),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_140),
.B1(n_152),
.B2(n_128),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_144),
.B(n_159),
.Y(n_177)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_6),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_141),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_149),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_143),
.A2(n_142),
.B(n_126),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_76),
.A2(n_116),
.B(n_71),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_92),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_93),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_9),
.C(n_10),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_81),
.C(n_73),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_11),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_90),
.B1(n_106),
.B2(n_80),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_12),
.B1(n_93),
.B2(n_84),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_172)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_84),
.B1(n_95),
.B2(n_88),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_80),
.A2(n_77),
.B1(n_95),
.B2(n_106),
.Y(n_159)
);

BUFx2_ASAP7_75t_SL g160 ( 
.A(n_77),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_104),
.Y(n_161)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_163),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_161),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_204),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_86),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_168),
.A2(n_178),
.B(n_181),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_81),
.CI(n_73),
.CON(n_169),
.SN(n_169)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_169),
.B(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_132),
.B1(n_150),
.B2(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_89),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_202),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_153),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_125),
.A2(n_152),
.B(n_131),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_133),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_191),
.B1(n_193),
.B2(n_178),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_146),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_205),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_128),
.A2(n_158),
.B1(n_120),
.B2(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_121),
.B(n_137),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_123),
.B(n_147),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_201),
.B(n_206),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_163),
.Y(n_201)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_145),
.A2(n_151),
.A3(n_162),
.B1(n_130),
.B2(n_141),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_134),
.B(n_145),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_189),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_122),
.B(n_124),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_211),
.B1(n_217),
.B2(n_223),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_235),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_191),
.B1(n_171),
.B2(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_194),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_175),
.B1(n_168),
.B2(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_169),
.B1(n_201),
.B2(n_176),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_227),
.B1(n_229),
.B2(n_238),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_225),
.B(n_199),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_177),
.A2(n_169),
.B1(n_201),
.B2(n_202),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_169),
.B1(n_201),
.B2(n_206),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_206),
.B(n_187),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_228),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_241),
.Y(n_262)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_234),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_237),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_173),
.A2(n_179),
.B1(n_180),
.B2(n_188),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_179),
.B(n_180),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_188),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.C(n_226),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_252),
.C(n_264),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_246),
.A2(n_253),
.B(n_233),
.Y(n_282)
);

AOI22x1_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_227),
.B1(n_240),
.B2(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_253),
.B1(n_257),
.B2(n_261),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_251),
.B(n_236),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_230),
.B(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_196),
.C(n_207),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_226),
.A2(n_173),
.B(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_210),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_242),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_213),
.C(n_223),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_267),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_200),
.C(n_190),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_211),
.B(n_200),
.C(n_174),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_215),
.B(n_186),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_186),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

XOR2x2_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_277),
.Y(n_305)
);

OAI322xp33_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_209),
.A3(n_222),
.B1(n_220),
.B2(n_219),
.C1(n_239),
.C2(n_241),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_279),
.A2(n_280),
.B(n_281),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_225),
.B(n_237),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_239),
.C(n_238),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_283),
.B(n_285),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_248),
.A2(n_208),
.B(n_234),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_296),
.B1(n_249),
.B2(n_255),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_245),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_212),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_298),
.B1(n_299),
.B2(n_274),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_247),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_254),
.A2(n_266),
.B1(n_261),
.B2(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

OAI321xp33_ASAP7_75t_L g299 ( 
.A1(n_262),
.A2(n_242),
.A3(n_251),
.B1(n_250),
.B2(n_254),
.C(n_258),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_252),
.C(n_267),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_303),
.C(n_308),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_264),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_310),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_257),
.C(n_270),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_280),
.B1(n_275),
.B2(n_286),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_256),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_286),
.B1(n_293),
.B2(n_288),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_309),
.A2(n_287),
.B1(n_298),
.B2(n_272),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_274),
.C(n_265),
.Y(n_310)
);

NAND4xp25_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_263),
.C(n_255),
.D(n_268),
.Y(n_311)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_315),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_260),
.C(n_268),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_249),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_287),
.Y(n_325)
);

XOR2x2_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_276),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_318),
.A2(n_309),
.B(n_305),
.Y(n_338)
);

NAND4xp25_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_285),
.C(n_279),
.D(n_283),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_319),
.A2(n_306),
.B1(n_316),
.B2(n_259),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_289),
.B1(n_275),
.B2(n_272),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_308),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_282),
.B(n_290),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_324),
.B(n_330),
.C(n_315),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_320),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_326),
.B(n_328),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_259),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_318),
.A2(n_314),
.B(n_305),
.C(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_332),
.B(n_337),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_303),
.C(n_301),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_336),
.C(n_339),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_310),
.B1(n_330),
.B2(n_306),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_338),
.A2(n_325),
.B(n_328),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_342),
.C(n_327),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_327),
.A2(n_300),
.B1(n_324),
.B2(n_323),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_346),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_331),
.C(n_329),
.Y(n_347)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_342),
.B(n_336),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_SL g350 ( 
.A(n_343),
.B(n_337),
.C(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_350),
.B(n_351),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_348),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_352),
.B(n_344),
.CI(n_331),
.CON(n_353),
.SN(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_349),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_354),
.B(n_329),
.Y(n_356)
);

AOI321xp33_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_340),
.A3(n_335),
.B1(n_332),
.B2(n_353),
.C(n_334),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_353),
.Y(n_358)
);


endmodule