module fake_jpeg_28251_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_SL g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_20),
.B1(n_14),
.B2(n_9),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

AND2x6_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_1),
.B1(n_6),
.B2(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_26),
.B(n_12),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_9),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_8),
.C(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_24),
.B1(n_12),
.B2(n_22),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_23),
.B(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_10),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_10),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_1),
.C(n_10),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_42),
.B1(n_24),
.B2(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_40),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_50),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_49),
.Y(n_58)
);


endmodule