module fake_jpeg_2281_n_230 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_0),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_36),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_84),
.Y(n_86)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_1),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_80),
.B1(n_57),
.B2(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_96),
.B1(n_71),
.B2(n_56),
.Y(n_100)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_67),
.B1(n_82),
.B2(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_58),
.B1(n_73),
.B2(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_94),
.Y(n_107)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_64),
.B1(n_60),
.B2(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_71),
.B(n_69),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_116),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_65),
.Y(n_133)
);

OR2x6_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_70),
.B1(n_56),
.B2(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_31),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_138),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_66),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_74),
.A3(n_66),
.B1(n_85),
.B2(n_55),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_74),
.B(n_77),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_76),
.B(n_75),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_61),
.B(n_6),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_137),
.B(n_72),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_147),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_70),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_2),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_55),
.B1(n_85),
.B2(n_61),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_152),
.B1(n_119),
.B2(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_23),
.C(n_52),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_2),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_61),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_3),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_162),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_26),
.C(n_49),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_160),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_128),
.B1(n_135),
.B2(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_50),
.B1(n_45),
.B2(n_43),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_25),
.C(n_47),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_119),
.B(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_176),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_150),
.B1(n_148),
.B2(n_12),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_42),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_179),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_194),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_9),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_11),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_168),
.B(n_175),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_205),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_166),
.B1(n_176),
.B2(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_203),
.B1(n_208),
.B2(n_13),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_170),
.B1(n_174),
.B2(n_14),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_32),
.B(n_30),
.Y(n_216)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_27),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_191),
.C(n_190),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_185),
.B(n_189),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_213),
.B(n_28),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_214),
.Y(n_217)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_40),
.B(n_37),
.C(n_35),
.D(n_34),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_11),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.C(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_206),
.B1(n_200),
.B2(n_207),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_220),
.B(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_219),
.B1(n_221),
.B2(n_217),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.C(n_15),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_13),
.B(n_14),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_16),
.C(n_17),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_228),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_18),
.Y(n_230)
);


endmodule