module fake_jpeg_31539_n_126 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_22),
.C(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_18),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_27),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_20),
.B1(n_19),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_59),
.B1(n_32),
.B2(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_47),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_50),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_28),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_16),
.C(n_25),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_39),
.B(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_78)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_59),
.B1(n_51),
.B2(n_46),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_51),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_55),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_71),
.C(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_71),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_47),
.B1(n_50),
.B2(n_46),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_70),
.B(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_76),
.B1(n_60),
.B2(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_97),
.C(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_78),
.B1(n_96),
.B2(n_89),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_72),
.C(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_81),
.B(n_79),
.C(n_84),
.D(n_78),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_106),
.C(n_101),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_88),
.B(n_42),
.C(n_71),
.D(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_97),
.C(n_95),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_111),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_64),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_80),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_106),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_103),
.B(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_113),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_121),
.B(n_117),
.Y(n_122)
);

AOI31xp33_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_118),
.A3(n_48),
.B(n_12),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_123),
.B(n_10),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_11),
.B(n_12),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_48),
.Y(n_126)
);


endmodule