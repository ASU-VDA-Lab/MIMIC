module fake_aes_12322_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AOI22xp5_ASAP7_75t_L g11 ( .A1(n_2), .A2(n_5), .B1(n_9), .B2(n_1), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
A2O1A1Ixp33_ASAP7_75t_L g17 ( .A1(n_14), .A2(n_0), .B(n_1), .C(n_2), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
AO21x1_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_14), .B(n_11), .Y(n_19) );
NAND2xp33_ASAP7_75t_L g20 ( .A(n_18), .B(n_15), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_19), .B(n_16), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_17), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_0), .Y(n_25) );
INVx3_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_23), .B1(n_18), .B2(n_0), .Y(n_27) );
NAND5xp2_ASAP7_75t_L g28 ( .A(n_26), .B(n_1), .C(n_3), .D(n_4), .E(n_6), .Y(n_28) );
OAI22xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_18), .B1(n_4), .B2(n_7), .Y(n_29) );
NAND4xp75_ASAP7_75t_L g30 ( .A(n_28), .B(n_3), .C(n_8), .D(n_9), .Y(n_30) );
NOR2x1_ASAP7_75t_L g31 ( .A(n_28), .B(n_18), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_27), .B(n_18), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_29), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
OAI22x1_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_30), .B1(n_10), .B2(n_8), .Y(n_35) );
XNOR2xp5_ASAP7_75t_L g36 ( .A(n_35), .B(n_34), .Y(n_36) );
endmodule