module real_aes_5613_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_889;
wire n_696;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_892;
wire n_528;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_922;
wire n_633;
wire n_482;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_0), .A2(n_57), .B1(n_373), .B2(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_1), .A2(n_219), .B1(n_451), .B2(n_452), .Y(n_565) );
AO22x2_ASAP7_75t_L g547 ( .A1(n_2), .A2(n_548), .B1(n_567), .B2(n_568), .Y(n_547) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_2), .Y(n_567) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_3), .Y(n_654) );
AND2x4_ASAP7_75t_L g666 ( .A(n_3), .B(n_239), .Y(n_666) );
AND2x4_ASAP7_75t_L g671 ( .A(n_3), .B(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_4), .A2(n_47), .B1(n_694), .B2(n_695), .Y(n_701) );
INVx1_ASAP7_75t_L g893 ( .A(n_5), .Y(n_893) );
INVx1_ASAP7_75t_L g471 ( .A(n_6), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_7), .A2(n_90), .B1(n_885), .B2(n_887), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_8), .A2(n_183), .B1(n_373), .B2(n_411), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_9), .A2(n_98), .B1(n_663), .B2(n_667), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_10), .A2(n_81), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_11), .A2(n_210), .B1(n_410), .B2(n_518), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_12), .A2(n_15), .B1(n_445), .B2(n_446), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_13), .A2(n_23), .B1(n_415), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_14), .A2(n_193), .B1(n_383), .B2(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_16), .A2(n_107), .B1(n_937), .B2(n_938), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_17), .A2(n_29), .B1(n_459), .B2(n_460), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_18), .B(n_404), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_19), .A2(n_917), .B1(n_918), .B2(n_948), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_19), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_20), .A2(n_25), .B1(n_432), .B2(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_21), .A2(n_140), .B1(n_448), .B2(n_449), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_22), .A2(n_70), .B1(n_385), .B2(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_24), .A2(n_199), .B1(n_343), .B2(n_351), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_26), .A2(n_108), .B1(n_396), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_27), .A2(n_175), .B1(n_351), .B2(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_28), .Y(n_356) );
INVx1_ASAP7_75t_L g492 ( .A(n_30), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_31), .A2(n_189), .B1(n_294), .B2(n_460), .Y(n_585) );
INVx1_ASAP7_75t_L g365 ( .A(n_32), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_33), .A2(n_94), .B1(n_379), .B2(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g607 ( .A(n_34), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_35), .A2(n_319), .B(n_321), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_36), .A2(n_91), .B1(n_690), .B2(n_692), .Y(n_700) );
XNOR2x1_ASAP7_75t_L g484 ( .A(n_37), .B(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_38), .A2(n_157), .B1(n_940), .B2(n_941), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_39), .A2(n_467), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g402 ( .A(n_40), .Y(n_402) );
INVx1_ASAP7_75t_L g280 ( .A(n_41), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_41), .B(n_177), .Y(n_329) );
INVxp67_ASAP7_75t_L g350 ( .A(n_41), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_42), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_43), .A2(n_88), .B1(n_413), .B2(n_417), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_44), .A2(n_115), .B1(n_309), .B2(n_943), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_45), .A2(n_158), .B1(n_694), .B2(n_695), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_46), .A2(n_227), .B1(n_683), .B2(n_686), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g254 ( .A(n_47), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_48), .B(n_264), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_49), .A2(n_75), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI21xp33_ASAP7_75t_SL g550 ( .A1(n_50), .A2(n_474), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_51), .A2(n_228), .B1(n_432), .B2(n_433), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_52), .A2(n_151), .B1(n_336), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_53), .A2(n_202), .B1(n_303), .B2(n_305), .Y(n_302) );
BUFx2_ASAP7_75t_L g557 ( .A(n_54), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_55), .A2(n_87), .B1(n_445), .B2(n_446), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_56), .A2(n_102), .B1(n_663), .B2(n_667), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_58), .A2(n_178), .B1(n_445), .B2(n_446), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_59), .A2(n_237), .B1(n_303), .B2(n_305), .Y(n_593) );
INVx2_ASAP7_75t_L g652 ( .A(n_60), .Y(n_652) );
INVx1_ASAP7_75t_L g665 ( .A(n_61), .Y(n_665) );
AND2x4_ASAP7_75t_L g668 ( .A(n_61), .B(n_652), .Y(n_668) );
INVx1_ASAP7_75t_SL g691 ( .A(n_61), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_62), .A2(n_182), .B1(n_448), .B2(n_449), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_63), .A2(n_138), .B1(n_336), .B2(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_64), .A2(n_149), .B1(n_359), .B2(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_65), .B(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_66), .A2(n_205), .B1(n_430), .B2(n_433), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_67), .A2(n_223), .B1(n_373), .B2(n_411), .Y(n_628) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_68), .Y(n_264) );
XNOR2x2_ASAP7_75t_SL g590 ( .A(n_69), .B(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_69), .A2(n_139), .B1(n_694), .B2(n_695), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_71), .A2(n_179), .B1(n_448), .B2(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g509 ( .A(n_72), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_73), .A2(n_162), .B1(n_524), .B2(n_527), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_74), .A2(n_169), .B1(n_303), .B2(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_76), .A2(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g680 ( .A(n_77), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_78), .A2(n_245), .B1(n_690), .B2(n_692), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_79), .A2(n_197), .B1(n_380), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_80), .A2(n_133), .B1(n_351), .B2(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g265 ( .A(n_82), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_82), .B(n_176), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_83), .A2(n_229), .B1(n_305), .B2(n_372), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_84), .A2(n_89), .B1(n_690), .B2(n_692), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_85), .A2(n_209), .B1(n_410), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_86), .A2(n_153), .B1(n_258), .B2(n_283), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_92), .A2(n_194), .B1(n_319), .B2(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_93), .A2(n_135), .B1(n_336), .B2(n_578), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_95), .A2(n_215), .B1(n_611), .B2(n_612), .C(n_613), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_96), .A2(n_161), .B1(n_641), .B2(n_642), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_97), .A2(n_224), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_99), .A2(n_116), .B1(n_518), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_100), .A2(n_187), .B1(n_410), .B2(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g619 ( .A(n_101), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_101), .A2(n_181), .B1(n_686), .B2(n_694), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_103), .A2(n_244), .B1(n_442), .B2(n_443), .Y(n_563) );
INVxp33_ASAP7_75t_SL g687 ( .A(n_104), .Y(n_687) );
XNOR2x1_ASAP7_75t_L g455 ( .A(n_105), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_106), .A2(n_117), .B1(n_921), .B2(n_922), .Y(n_920) );
INVx1_ASAP7_75t_L g614 ( .A(n_109), .Y(n_614) );
INVx1_ASAP7_75t_L g931 ( .A(n_110), .Y(n_931) );
INVx1_ASAP7_75t_L g552 ( .A(n_111), .Y(n_552) );
INVx1_ASAP7_75t_L g464 ( .A(n_112), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_113), .A2(n_142), .B1(n_670), .B2(n_673), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_114), .A2(n_121), .B1(n_905), .B2(n_906), .Y(n_904) );
INVx1_ASAP7_75t_L g494 ( .A(n_118), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_119), .A2(n_166), .B1(n_283), .B2(n_370), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_120), .A2(n_238), .B1(n_442), .B2(n_443), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_122), .A2(n_143), .B1(n_294), .B2(n_299), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_123), .A2(n_206), .B1(n_334), .B2(n_433), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_124), .A2(n_126), .B1(n_351), .B2(n_376), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_125), .A2(n_359), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g602 ( .A(n_127), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_128), .A2(n_130), .B1(n_305), .B2(n_385), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_129), .A2(n_213), .B1(n_899), .B2(n_901), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_131), .A2(n_168), .B1(n_334), .B2(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g570 ( .A(n_132), .Y(n_570) );
INVx1_ASAP7_75t_L g322 ( .A(n_134), .Y(n_322) );
INVx1_ASAP7_75t_L g684 ( .A(n_136), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_137), .B(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_141), .A2(n_164), .B1(n_945), .B2(n_946), .Y(n_944) );
INVx1_ASAP7_75t_L g425 ( .A(n_144), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_145), .A2(n_226), .B1(n_309), .B2(n_313), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_146), .A2(n_195), .B1(n_303), .B2(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_147), .B(n_367), .Y(n_539) );
XOR2xp5_ASAP7_75t_L g389 ( .A(n_148), .B(n_390), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_150), .A2(n_216), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_152), .A2(n_170), .B1(n_885), .B2(n_924), .Y(n_923) );
OA22x2_ASAP7_75t_L g270 ( .A1(n_154), .A2(n_177), .B1(n_264), .B2(n_268), .Y(n_270) );
INVx1_ASAP7_75t_L g290 ( .A(n_154), .Y(n_290) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_155), .A2(n_927), .B(n_930), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_156), .A2(n_247), .B1(n_370), .B2(n_411), .Y(n_504) );
XOR2x2_ASAP7_75t_L g513 ( .A(n_159), .B(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_160), .A2(n_235), .B1(n_670), .B2(n_673), .Y(n_717) );
INVx1_ASAP7_75t_L g934 ( .A(n_163), .Y(n_934) );
INVx1_ASAP7_75t_L g609 ( .A(n_165), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_167), .A2(n_231), .B1(n_385), .B2(n_387), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_171), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_172), .B(n_400), .Y(n_428) );
BUFx2_ASAP7_75t_L g559 ( .A(n_173), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_174), .A2(n_204), .B1(n_448), .B2(n_449), .Y(n_566) );
INVx1_ASAP7_75t_L g282 ( .A(n_176), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_176), .B(n_288), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g291 ( .A1(n_177), .A2(n_198), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g777 ( .A(n_180), .Y(n_777) );
INVx1_ASAP7_75t_L g776 ( .A(n_184), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_184), .A2(n_914), .B1(n_916), .B2(n_949), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_185), .A2(n_203), .B1(n_690), .B2(n_692), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_186), .A2(n_207), .B1(n_595), .B2(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g490 ( .A(n_188), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_190), .A2(n_225), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI221x1_ASAP7_75t_SL g358 ( .A1(n_191), .A2(n_192), .B1(n_359), .B2(n_361), .C(n_364), .Y(n_358) );
INVx1_ASAP7_75t_L g634 ( .A(n_196), .Y(n_634) );
INVx1_ASAP7_75t_L g267 ( .A(n_198), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_198), .B(n_230), .Y(n_330) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_200), .A2(n_359), .B(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_201), .A2(n_234), .B1(n_506), .B2(n_507), .C(n_508), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_208), .A2(n_889), .B(n_892), .Y(n_888) );
INVx1_ASAP7_75t_L g581 ( .A(n_211), .Y(n_581) );
INVx1_ASAP7_75t_L g437 ( .A(n_212), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_214), .A2(n_233), .B1(n_309), .B2(n_383), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_217), .A2(n_435), .B(n_436), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_218), .A2(n_222), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_220), .A2(n_241), .B1(n_373), .B2(n_584), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_221), .A2(n_534), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_230), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_232), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_236), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g672 ( .A(n_239), .Y(n_672) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_239), .Y(n_951) );
INVxp33_ASAP7_75t_L g678 ( .A(n_240), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_242), .A2(n_243), .B1(n_309), .B2(n_383), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_246), .A2(n_248), .B1(n_383), .B2(n_415), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_540), .B(n_646), .C(n_655), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_250), .A2(n_540), .B(n_647), .Y(n_646) );
XNOR2xp5_ASAP7_75t_SL g250 ( .A(n_251), .B(n_420), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_353), .B1(n_418), .B2(n_419), .Y(n_251) );
INVx1_ASAP7_75t_L g418 ( .A(n_252), .Y(n_418) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
NOR2x1_ASAP7_75t_L g255 ( .A(n_256), .B(n_317), .Y(n_255) );
NAND4xp25_ASAP7_75t_L g256 ( .A(n_257), .B(n_293), .C(n_302), .D(n_308), .Y(n_256) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_259), .Y(n_373) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_259), .Y(n_500) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_259), .Y(n_595) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_271), .Y(n_259) );
AND2x4_ASAP7_75t_L g304 ( .A(n_260), .B(n_297), .Y(n_304) );
AND2x4_ASAP7_75t_L g310 ( .A(n_260), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g314 ( .A(n_260), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g442 ( .A(n_260), .B(n_301), .Y(n_442) );
AND2x4_ASAP7_75t_L g448 ( .A(n_260), .B(n_311), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_260), .B(n_315), .Y(n_449) );
AND2x4_ASAP7_75t_L g451 ( .A(n_260), .B(n_297), .Y(n_451) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_269), .Y(n_260) );
AND2x2_ASAP7_75t_L g320 ( .A(n_261), .B(n_270), .Y(n_320) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g296 ( .A(n_262), .B(n_270), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
NAND2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g268 ( .A(n_264), .Y(n_268) );
INVx3_ASAP7_75t_L g275 ( .A(n_264), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_264), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_264), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_265), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_267), .A2(n_292), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g348 ( .A(n_270), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g285 ( .A(n_271), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g443 ( .A(n_271), .B(n_286), .Y(n_443) );
AND2x4_ASAP7_75t_L g446 ( .A(n_271), .B(n_296), .Y(n_446) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
AND2x4_ASAP7_75t_L g297 ( .A(n_273), .B(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_L g311 ( .A(n_273), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g316 ( .A(n_273), .Y(n_316) );
AND2x2_ASAP7_75t_L g345 ( .A(n_273), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g288 ( .A(n_275), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_276), .B(n_287), .C(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g312 ( .A(n_278), .Y(n_312) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx5_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g584 ( .A(n_284), .Y(n_584) );
INVx3_ASAP7_75t_L g596 ( .A(n_284), .Y(n_596) );
INVx6_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx12f_ASAP7_75t_L g411 ( .A(n_285), .Y(n_411) );
AND2x4_ASAP7_75t_L g307 ( .A(n_286), .B(n_297), .Y(n_307) );
AND2x4_ASAP7_75t_L g337 ( .A(n_286), .B(n_315), .Y(n_337) );
AND2x4_ASAP7_75t_L g433 ( .A(n_286), .B(n_315), .Y(n_433) );
AND2x4_ASAP7_75t_L g452 ( .A(n_286), .B(n_297), .Y(n_452) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
BUFx4f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_295), .Y(n_459) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x4_ASAP7_75t_L g300 ( .A(n_296), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g341 ( .A(n_296), .B(n_315), .Y(n_341) );
AND2x2_ASAP7_75t_L g352 ( .A(n_296), .B(n_311), .Y(n_352) );
AND2x2_ASAP7_75t_L g386 ( .A(n_296), .B(n_297), .Y(n_386) );
AND2x4_ASAP7_75t_L g430 ( .A(n_296), .B(n_311), .Y(n_430) );
AND2x4_ASAP7_75t_L g445 ( .A(n_296), .B(n_297), .Y(n_445) );
AND2x2_ASAP7_75t_L g469 ( .A(n_296), .B(n_315), .Y(n_469) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx12f_ASAP7_75t_L g370 ( .A(n_300), .Y(n_370) );
BUFx3_ASAP7_75t_L g410 ( .A(n_300), .Y(n_410) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_300), .Y(n_460) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_300), .Y(n_519) );
BUFx12f_ASAP7_75t_L g521 ( .A(n_303), .Y(n_521) );
INVx1_ASAP7_75t_L g900 ( .A(n_303), .Y(n_900) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_304), .Y(n_372) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_304), .Y(n_413) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g387 ( .A(n_306), .Y(n_387) );
INVx4_ASAP7_75t_L g417 ( .A(n_306), .Y(n_417) );
INVx1_ASAP7_75t_L g462 ( .A(n_306), .Y(n_462) );
INVx1_ASAP7_75t_L g522 ( .A(n_306), .Y(n_522) );
INVx4_ASAP7_75t_L g908 ( .A(n_306), .Y(n_908) );
INVx1_ASAP7_75t_L g947 ( .A(n_306), .Y(n_947) );
INVx8_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_310), .Y(n_415) );
INVx3_ASAP7_75t_L g526 ( .A(n_310), .Y(n_526) );
AND2x4_ASAP7_75t_L g319 ( .A(n_311), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g360 ( .A(n_311), .B(n_320), .Y(n_360) );
AND2x4_ASAP7_75t_L g315 ( .A(n_312), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g906 ( .A(n_313), .Y(n_906) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_314), .Y(n_383) );
BUFx5_ASAP7_75t_L g527 ( .A(n_314), .Y(n_527) );
INVx1_ASAP7_75t_L g625 ( .A(n_314), .Y(n_625) );
AND2x4_ASAP7_75t_L g335 ( .A(n_315), .B(n_320), .Y(n_335) );
AND2x2_ASAP7_75t_L g435 ( .A(n_315), .B(n_320), .Y(n_435) );
NAND4xp25_ASAP7_75t_SL g317 ( .A(n_318), .B(n_333), .C(n_338), .D(n_342), .Y(n_317) );
INVx2_ASAP7_75t_L g603 ( .A(n_319), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_323), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_323), .B(n_614), .Y(n_613) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g367 ( .A(n_324), .Y(n_367) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_324), .Y(n_407) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g439 ( .A(n_325), .Y(n_439) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_327), .B(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_328), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g465 ( .A(n_334), .Y(n_465) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx8_ASAP7_75t_SL g379 ( .A(n_335), .Y(n_379) );
INVx2_ASAP7_75t_L g397 ( .A(n_335), .Y(n_397) );
BUFx3_ASAP7_75t_L g506 ( .A(n_335), .Y(n_506) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_335), .Y(n_578) );
INVx3_ASAP7_75t_L g491 ( .A(n_336), .Y(n_491) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
INVx3_ASAP7_75t_L g883 ( .A(n_337), .Y(n_883) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g576 ( .A(n_340), .Y(n_576) );
INVx2_ASAP7_75t_L g639 ( .A(n_340), .Y(n_639) );
INVx2_ASAP7_75t_L g891 ( .A(n_340), .Y(n_891) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g363 ( .A(n_341), .Y(n_363) );
BUFx3_ASAP7_75t_L g534 ( .A(n_341), .Y(n_534) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx5_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
BUFx4f_ASAP7_75t_L g497 ( .A(n_344), .Y(n_497) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_348), .Y(n_344) );
AND2x4_ASAP7_75t_L g404 ( .A(n_345), .B(n_348), .Y(n_404) );
AND2x2_ASAP7_75t_L g432 ( .A(n_345), .B(n_348), .Y(n_432) );
INVx2_ASAP7_75t_L g925 ( .A(n_351), .Y(n_925) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_352), .Y(n_489) );
INVx2_ASAP7_75t_L g538 ( .A(n_352), .Y(n_538) );
INVx1_ASAP7_75t_L g419 ( .A(n_353), .Y(n_419) );
XNOR2x1_ASAP7_75t_L g353 ( .A(n_354), .B(n_388), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
XOR2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND4xp75_ASAP7_75t_L g357 ( .A(n_358), .B(n_368), .C(n_374), .D(n_381), .Y(n_357) );
INVx4_ASAP7_75t_L g495 ( .A(n_359), .Y(n_495) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
BUFx3_ASAP7_75t_L g474 ( .A(n_360), .Y(n_474) );
BUFx3_ASAP7_75t_L g886 ( .A(n_360), .Y(n_886) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g507 ( .A(n_362), .Y(n_507) );
INVx2_ASAP7_75t_L g929 ( .A(n_362), .Y(n_929) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
BUFx2_ASAP7_75t_SL g940 ( .A(n_372), .Y(n_940) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g530 ( .A(n_377), .Y(n_530) );
INVx2_ASAP7_75t_L g574 ( .A(n_377), .Y(n_574) );
INVx2_ASAP7_75t_L g641 ( .A(n_377), .Y(n_641) );
HB1xp67_ASAP7_75t_L g921 ( .A(n_379), .Y(n_921) );
BUFx3_ASAP7_75t_L g922 ( .A(n_380), .Y(n_922) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
BUFx3_ASAP7_75t_L g945 ( .A(n_385), .Y(n_945) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx8_ASAP7_75t_L g518 ( .A(n_386), .Y(n_518) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2x1_ASAP7_75t_SL g390 ( .A(n_391), .B(n_408), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_395), .C(n_398), .Y(n_391) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g636 ( .A(n_397), .Y(n_636) );
BUFx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_405), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_403), .A2(n_556), .B1(n_558), .B2(n_560), .Y(n_555) );
INVx4_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_407), .B(n_581), .Y(n_580) );
NAND4xp25_ASAP7_75t_SL g408 ( .A(n_409), .B(n_412), .C(n_414), .D(n_416), .Y(n_408) );
BUFx3_ASAP7_75t_L g938 ( .A(n_411), .Y(n_938) );
XNOR2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_481), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_453), .B2(n_479), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
XNOR2x1_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_440), .Y(n_426) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .C(n_431), .D(n_434), .Y(n_427) );
INVx2_ASAP7_75t_L g560 ( .A(n_430), .Y(n_560) );
INVx1_ASAP7_75t_L g606 ( .A(n_430), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_433), .Y(n_608) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_435), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx4_ASAP7_75t_L g511 ( .A(n_438), .Y(n_511) );
INVx1_ASAP7_75t_L g896 ( .A(n_438), .Y(n_896) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g553 ( .A(n_439), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .C(n_447), .D(n_450), .Y(n_440) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g480 ( .A(n_455), .Y(n_480) );
NAND4xp75_ASAP7_75t_L g456 ( .A(n_457), .B(n_463), .C(n_472), .D(n_476), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .Y(n_457) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g881 ( .A(n_465), .Y(n_881) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_469), .Y(n_611) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_512), .B2(n_513), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND4xp75_ASAP7_75t_L g485 ( .A(n_486), .B(n_498), .C(n_502), .D(n_505), .Y(n_485) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g887 ( .A(n_489), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_496), .Y(n_493) );
INVx2_ASAP7_75t_SL g894 ( .A(n_497), .Y(n_894) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
BUFx3_ASAP7_75t_L g941 ( .A(n_500), .Y(n_941) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_528), .Y(n_514) );
NAND4xp25_ASAP7_75t_SL g515 ( .A(n_516), .B(n_517), .C(n_520), .D(n_523), .Y(n_515) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_519), .Y(n_937) );
BUFx4f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g905 ( .A(n_526), .Y(n_905) );
BUFx3_ASAP7_75t_L g943 ( .A(n_527), .Y(n_943) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .C(n_535), .D(n_539), .Y(n_528) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g642 ( .A(n_537), .Y(n_642) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_588), .B2(n_645), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
XOR2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_569), .Y(n_546) );
INVx1_ASAP7_75t_L g568 ( .A(n_548), .Y(n_568) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_549), .B(n_562), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .C(n_561), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_553), .B(n_634), .Y(n_633) );
INVx4_ASAP7_75t_L g933 ( .A(n_553), .Y(n_933) );
CKINVDCx16_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
CKINVDCx9p33_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .C(n_565), .D(n_566), .Y(n_562) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NOR2xp67_ASAP7_75t_L g571 ( .A(n_572), .B(n_582), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .C(n_577), .D(n_579), .Y(n_572) );
NAND4xp25_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .C(n_586), .D(n_587), .Y(n_582) );
BUFx2_ASAP7_75t_L g903 ( .A(n_584), .Y(n_903) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AO22x2_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_615), .B1(n_643), .B2(n_644), .Y(n_589) );
INVx2_ASAP7_75t_L g643 ( .A(n_590), .Y(n_643) );
NAND4xp75_ASAP7_75t_L g591 ( .A(n_592), .B(n_597), .C(n_600), .D(n_610), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
BUFx3_ASAP7_75t_L g901 ( .A(n_595), .Y(n_901) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_604), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_605) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g644 ( .A(n_617), .Y(n_644) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
XNOR2x1_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NOR2x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_629), .Y(n_620) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .C(n_627), .D(n_628), .Y(n_621) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_637), .C(n_640), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx10_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .C(n_654), .Y(n_649) );
AND2x2_ASAP7_75t_L g910 ( .A(n_650), .B(n_911), .Y(n_910) );
AND2x2_ASAP7_75t_L g915 ( .A(n_650), .B(n_912), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g952 ( .A1(n_650), .A2(n_654), .B(n_691), .Y(n_952) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AO21x1_ASAP7_75t_L g950 ( .A1(n_651), .A2(n_951), .B(n_952), .Y(n_950) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g664 ( .A(n_652), .B(n_665), .Y(n_664) );
AND3x4_ASAP7_75t_L g690 ( .A(n_652), .B(n_671), .C(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_653), .B(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_654), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_873), .B1(n_876), .B2(n_909), .C(n_913), .Y(n_655) );
AOI211x1_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_773), .B(n_779), .C(n_854), .Y(n_656) );
NAND5xp2_ASAP7_75t_L g657 ( .A(n_658), .B(n_731), .C(n_749), .D(n_759), .E(n_764), .Y(n_657) );
AOI332xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_696), .A3(n_706), .B1(n_707), .B2(n_711), .B3(n_720), .C1(n_721), .C2(n_725), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_674), .Y(n_659) );
INVx2_ASAP7_75t_L g719 ( .A(n_660), .Y(n_719) );
BUFx3_ASAP7_75t_L g792 ( .A(n_660), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_660), .B(n_715), .Y(n_799) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g729 ( .A(n_661), .Y(n_729) );
OR2x2_ASAP7_75t_L g826 ( .A(n_661), .B(n_688), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_669), .Y(n_661) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
AND2x4_ASAP7_75t_L g670 ( .A(n_664), .B(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g683 ( .A(n_664), .B(n_666), .Y(n_683) );
AND2x2_ASAP7_75t_L g694 ( .A(n_664), .B(n_666), .Y(n_694) );
AND2x2_ASAP7_75t_L g667 ( .A(n_666), .B(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g686 ( .A(n_666), .B(n_668), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_666), .B(n_668), .Y(n_695) );
AND2x4_ASAP7_75t_L g673 ( .A(n_668), .B(n_671), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_668), .B(n_671), .Y(n_679) );
AND2x4_ASAP7_75t_L g692 ( .A(n_668), .B(n_671), .Y(n_692) );
INVx3_ASAP7_75t_L g677 ( .A(n_670), .Y(n_677) );
INVx1_ASAP7_75t_L g789 ( .A(n_674), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_674), .B(n_839), .Y(n_838) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_688), .Y(n_674) );
INVx1_ASAP7_75t_L g714 ( .A(n_675), .Y(n_714) );
INVx2_ASAP7_75t_L g752 ( .A(n_675), .Y(n_752) );
AND2x2_ASAP7_75t_L g760 ( .A(n_675), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g768 ( .A(n_675), .B(n_688), .Y(n_768) );
AND2x2_ASAP7_75t_L g771 ( .A(n_675), .B(n_715), .Y(n_771) );
AND2x2_ASAP7_75t_L g821 ( .A(n_675), .B(n_716), .Y(n_821) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_681), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_677), .A2(n_679), .B1(n_776), .B2(n_777), .C(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g875 ( .A(n_677), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_685), .B2(n_687), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_688), .Y(n_720) );
INVx2_ASAP7_75t_L g739 ( .A(n_688), .Y(n_739) );
OR2x2_ASAP7_75t_L g748 ( .A(n_688), .B(n_729), .Y(n_748) );
AND2x2_ASAP7_75t_L g761 ( .A(n_688), .B(n_729), .Y(n_761) );
AND2x2_ASAP7_75t_L g781 ( .A(n_688), .B(n_728), .Y(n_781) );
OR2x2_ASAP7_75t_L g810 ( .A(n_688), .B(n_752), .Y(n_810) );
AND2x2_ASAP7_75t_L g844 ( .A(n_688), .B(n_752), .Y(n_844) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_693), .Y(n_688) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_705), .Y(n_697) );
INVx1_ASAP7_75t_L g724 ( .A(n_698), .Y(n_724) );
OR2x2_ASAP7_75t_L g758 ( .A(n_698), .B(n_708), .Y(n_758) );
OAI32xp33_ASAP7_75t_L g863 ( .A1(n_698), .A2(n_763), .A3(n_780), .B1(n_839), .B2(n_859), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_698), .B(n_756), .Y(n_872) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
AND2x2_ASAP7_75t_L g706 ( .A(n_699), .B(n_702), .Y(n_706) );
INVx1_ASAP7_75t_L g736 ( .A(n_699), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_699), .B(n_707), .Y(n_747) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
OR2x2_ASAP7_75t_L g735 ( .A(n_702), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g754 ( .A(n_702), .Y(n_754) );
AND2x2_ASAP7_75t_L g772 ( .A(n_702), .B(n_722), .Y(n_772) );
AND2x2_ASAP7_75t_L g787 ( .A(n_702), .B(n_736), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_702), .B(n_707), .Y(n_798) );
AOI211xp5_ASAP7_75t_SL g866 ( .A1(n_702), .A2(n_867), .B(n_868), .C(n_869), .Y(n_866) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g742 ( .A(n_706), .B(n_722), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_706), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g832 ( .A(n_706), .B(n_707), .Y(n_832) );
NOR2x1_ASAP7_75t_R g732 ( .A(n_707), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g753 ( .A(n_707), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g795 ( .A(n_707), .B(n_787), .Y(n_795) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g723 ( .A(n_708), .Y(n_723) );
OR2x2_ASAP7_75t_L g763 ( .A(n_708), .B(n_735), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_708), .B(n_734), .Y(n_804) );
AND2x2_ASAP7_75t_L g828 ( .A(n_708), .B(n_754), .Y(n_828) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_719), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_713), .A2(n_721), .B1(n_750), .B2(n_757), .C(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g730 ( .A(n_714), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_714), .B(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_715), .B(n_734), .Y(n_733) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_715), .Y(n_745) );
INVx2_ASAP7_75t_L g756 ( .A(n_715), .Y(n_756) );
INVx2_ASAP7_75t_L g767 ( .A(n_715), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_715), .B(n_753), .Y(n_816) );
AND2x2_ASAP7_75t_L g827 ( .A(n_715), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g839 ( .A(n_715), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g870 ( .A(n_715), .B(n_746), .Y(n_870) );
INVx4_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_716), .B(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g808 ( .A(n_716), .B(n_722), .Y(n_808) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_719), .A2(n_750), .B(n_753), .C(n_755), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_719), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g802 ( .A(n_719), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_719), .B(n_855), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g869 ( .A1(n_720), .A2(n_735), .B1(n_810), .B2(n_870), .C(n_871), .Y(n_869) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_721), .A2(n_797), .B(n_799), .Y(n_796) );
AND2x2_ASAP7_75t_L g853 ( .A(n_721), .B(n_756), .Y(n_853) );
A2O1A1O1Ixp25_ASAP7_75t_L g856 ( .A1(n_721), .A2(n_795), .B(n_844), .C(n_857), .D(n_858), .Y(n_856) );
INVx2_ASAP7_75t_SL g862 ( .A(n_721), .Y(n_862) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
AND2x2_ASAP7_75t_L g786 ( .A(n_722), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_725), .A2(n_768), .B1(n_815), .B2(n_817), .C(n_819), .Y(n_814) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .Y(n_726) );
INVx1_ASAP7_75t_SL g857 ( .A(n_727), .Y(n_857) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_730), .B(n_781), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_730), .B(n_848), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_737), .B(n_740), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_734), .B(n_807), .Y(n_818) );
INVx3_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_736), .B(n_821), .Y(n_820) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_736), .A2(n_757), .B1(n_771), .B2(n_784), .C(n_872), .Y(n_871) );
CKINVDCx14_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g836 ( .A(n_739), .B(n_821), .Y(n_836) );
AOI21xp33_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_743), .B(n_748), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_742), .B(n_757), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_742), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
AND2x2_ASAP7_75t_L g831 ( .A(n_744), .B(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_744), .B(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_745), .B(n_754), .Y(n_846) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_747), .A2(n_833), .B(n_859), .C(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g823 ( .A(n_748), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_748), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g784 ( .A(n_752), .Y(n_784) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_756), .B(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_756), .B(n_758), .Y(n_813) );
INVx1_ASAP7_75t_L g849 ( .A(n_756), .Y(n_849) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
OAI21xp5_ASAP7_75t_L g811 ( .A1(n_761), .A2(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g851 ( .A(n_761), .Y(n_851) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI21xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_769), .B(n_772), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
NAND2xp67_ASAP7_75t_L g785 ( .A(n_767), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g845 ( .A(n_768), .Y(n_845) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g859 ( .A(n_771), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_772), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g842 ( .A(n_772), .Y(n_842) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AOI211xp5_ASAP7_75t_SL g840 ( .A1(n_774), .A2(n_841), .B(n_847), .C(n_850), .Y(n_840) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_775), .B(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g855 ( .A(n_775), .Y(n_855) );
XNOR2x1_ASAP7_75t_L g877 ( .A(n_776), .B(n_878), .Y(n_877) );
OAI211xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_782), .B(n_788), .C(n_840), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR2xp67_ASAP7_75t_SL g783 ( .A(n_784), .B(n_785), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_784), .B(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g793 ( .A(n_786), .Y(n_793) );
AOI211xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B(n_800), .C(n_829), .Y(n_788) );
OAI211xp5_ASAP7_75t_SL g790 ( .A1(n_791), .A2(n_793), .B(n_794), .C(n_796), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g812 ( .A(n_794), .Y(n_812) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND3xp33_ASAP7_75t_SL g800 ( .A(n_801), .B(n_811), .C(n_814), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_SL g801 ( .A1(n_802), .A2(n_803), .B(n_805), .C(n_809), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI21xp33_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_822), .B(n_824), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_833), .B1(n_834), .B2(n_835), .C(n_837), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_845), .B2(n_846), .Y(n_841) );
INVx1_ASAP7_75t_L g867 ( .A(n_843), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B1(n_864), .B2(n_866), .Y(n_854) );
NOR2xp33_ASAP7_75t_SL g860 ( .A(n_861), .B(n_863), .Y(n_860) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
OR2x2_ASAP7_75t_L g878 ( .A(n_879), .B(n_897), .Y(n_878) );
NAND3xp33_ASAP7_75t_SL g879 ( .A(n_880), .B(n_884), .C(n_888), .Y(n_879) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
BUFx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
OAI21xp33_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B(n_895), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_894), .A2(n_931), .B1(n_932), .B2(n_934), .Y(n_930) );
NAND4xp25_ASAP7_75t_L g897 ( .A(n_898), .B(n_902), .C(n_904), .D(n_907), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
BUFx3_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g948 ( .A(n_918), .Y(n_948) );
OR2x2_ASAP7_75t_L g918 ( .A(n_919), .B(n_935), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_923), .C(n_926), .Y(n_919) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_SL g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
NAND4xp25_ASAP7_75t_SL g935 ( .A(n_936), .B(n_939), .C(n_942), .D(n_944), .Y(n_935) );
BUFx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
endmodule