module real_jpeg_30475_n_31 (n_17, n_8, n_0, n_21, n_212, n_2, n_29, n_209, n_201, n_10, n_9, n_12, n_24, n_6, n_28, n_208, n_207, n_202, n_203, n_213, n_23, n_11, n_14, n_211, n_25, n_205, n_7, n_22, n_18, n_3, n_206, n_210, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_30, n_204, n_16, n_15, n_13, n_31);

input n_17;
input n_8;
input n_0;
input n_21;
input n_212;
input n_2;
input n_29;
input n_209;
input n_201;
input n_10;
input n_9;
input n_12;
input n_24;
input n_6;
input n_28;
input n_208;
input n_207;
input n_202;
input n_203;
input n_213;
input n_23;
input n_11;
input n_14;
input n_211;
input n_25;
input n_205;
input n_7;
input n_22;
input n_18;
input n_3;
input n_206;
input n_210;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_30;
input n_204;
input n_16;
input n_15;
input n_13;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_179;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_75),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_43),
.C(n_182),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_3),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_45),
.B1(n_47),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_9),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_10),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_81),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_11),
.B(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_33),
.C(n_186),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_12),
.B(n_35),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_41),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

AOI221xp5_ASAP7_75t_L g126 ( 
.A1(n_13),
.A2(n_22),
.B1(n_127),
.B2(n_132),
.C(n_134),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_13),
.B(n_127),
.C(n_132),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_14),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_14),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_15),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_15),
.B(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_16),
.Y(n_198)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_17),
.B(n_88),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_19),
.B(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_20),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_21),
.A2(n_99),
.A3(n_101),
.B1(n_105),
.B2(n_161),
.C1(n_163),
.C2(n_211),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_22),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_28),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_194),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_41),
.B(n_42),
.C(n_185),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_38),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_92),
.B(n_166),
.Y(n_43)
);

NAND4xp25_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.C(n_79),
.D(n_86),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_53),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_50),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_64),
.C(n_68),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_56),
.B(n_176),
.C(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_57),
.B(n_63),
.Y(n_170)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_60),
.Y(n_102)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g174 ( 
.A1(n_64),
.A2(n_70),
.A3(n_175),
.B1(n_178),
.B2(n_179),
.C1(n_180),
.C2(n_213),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_67),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_69),
.A2(n_169),
.A3(n_170),
.B1(n_171),
.B2(n_174),
.C(n_212),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_80),
.A2(n_168),
.B(n_181),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_90),
.Y(n_192)
);

AOI31xp67_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_115),
.A3(n_149),
.B(n_156),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.C(n_112),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_94),
.A2(n_157),
.B(n_160),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_96),
.B(n_112),
.C(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_202),
.Y(n_101)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_144),
.C(n_145),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_138),
.B(n_143),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_126),
.B1(n_136),
.B2(n_137),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_207),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_142),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

BUFx4f_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_201),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_203),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_204),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_205),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_206),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_208),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_209),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_210),
.Y(n_152)
);


endmodule