module fake_jpeg_23206_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_22),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_19),
.B1(n_13),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_7),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_1),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_15),
.B(n_33),
.C(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_57),
.Y(n_69)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_36),
.B1(n_30),
.B2(n_18),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_60),
.B1(n_62),
.B2(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_63),
.Y(n_71)
);

OAI21x1_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_16),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_64),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_51),
.Y(n_80)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_66),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_59),
.B1(n_55),
.B2(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

AO221x1_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_86),
.B1(n_70),
.B2(n_47),
.C(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_55),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_69),
.B(n_75),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_80),
.C(n_81),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_91),
.B1(n_93),
.B2(n_57),
.C(n_71),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_75),
.C(n_78),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_76),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_59),
.B(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_86),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_98),
.C(n_67),
.Y(n_100)
);

INVxp33_ASAP7_75t_SL g99 ( 
.A(n_94),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_101),
.B(n_95),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_98),
.Y(n_105)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

AOI31xp67_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_86),
.A3(n_53),
.B(n_48),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_107),
.Y(n_109)
);

AOI222xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_9),
.B1(n_10),
.B2(n_41),
.C1(n_84),
.C2(n_99),
.Y(n_110)
);


endmodule