module fake_jpeg_2565_n_43 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_43);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_17),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_14),
.B1(n_13),
.B2(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_23),
.B(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_1),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_13),
.C(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_1),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_3),
.B(n_5),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_36),
.B(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B1(n_37),
.B2(n_8),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_37),
.B(n_9),
.Y(n_43)
);


endmodule