module fake_jpeg_13107_n_249 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_44),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_65),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_6),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_39),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_80),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_22),
.B(n_38),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_36),
.B(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_12),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_52),
.C(n_65),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_58),
.C(n_48),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_1),
.B(n_3),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_22),
.B1(n_24),
.B2(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_20),
.B1(n_31),
.B2(n_49),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_41),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_64),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_28),
.B1(n_26),
.B2(n_40),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_103),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_47),
.B(n_58),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_99),
.A2(n_111),
.B(n_77),
.C(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_123),
.B1(n_71),
.B2(n_7),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_84),
.C(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_108),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_69),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_112),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_57),
.B1(n_53),
.B2(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_31),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_25),
.B(n_15),
.C(n_12),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_R g119 ( 
.A(n_85),
.B(n_1),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_126),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_61),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_96),
.Y(n_136)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_87),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_110),
.C(n_8),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_118),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_137),
.B1(n_139),
.B2(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_115),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_74),
.B1(n_84),
.B2(n_66),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_77),
.B1(n_101),
.B2(n_9),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_71),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_152),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_125),
.B1(n_99),
.B2(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_167),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_102),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_163),
.B(n_164),
.C(n_175),
.D(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_99),
.B(n_122),
.C(n_116),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_162),
.B(n_165),
.Y(n_178)
);

CKINVDCx12_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_126),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_100),
.B1(n_84),
.B2(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_138),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_170),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_109),
.B1(n_106),
.B2(n_101),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_172),
.B(n_142),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_176),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_6),
.B(n_9),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_6),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_187),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_195),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_170),
.B(n_142),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_193),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_143),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_154),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_178),
.B(n_160),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_202),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_133),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_137),
.B1(n_155),
.B2(n_160),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_205),
.A2(n_194),
.B1(n_188),
.B2(n_179),
.Y(n_211)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_138),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_151),
.Y(n_209)
);

AO221x1_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_180),
.B1(n_185),
.B2(n_144),
.C(n_146),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_217),
.B1(n_198),
.B2(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_190),
.B1(n_186),
.B2(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_177),
.C(n_160),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_205),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_178),
.B1(n_193),
.B2(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_200),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_227),
.B1(n_211),
.B2(n_221),
.Y(n_230)
);

XOR2x2_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_196),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_223),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_217),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_210),
.B(n_203),
.Y(n_229)
);

AOI21x1_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_201),
.B(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_232),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_199),
.B1(n_216),
.B2(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_235),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_214),
.C(n_181),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_219),
.C(n_202),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_236),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_224),
.A3(n_185),
.B1(n_206),
.B2(n_144),
.C1(n_146),
.C2(n_151),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_233),
.C(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_239),
.C(n_237),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_SL g246 ( 
.A(n_244),
.B(n_239),
.C(n_234),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_10),
.C(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_10),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_10),
.Y(n_249)
);


endmodule