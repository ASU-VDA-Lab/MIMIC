module fake_jpeg_13734_n_86 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_86);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_1),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_21),
.Y(n_36)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_29),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_25),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_39),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_44),
.B1(n_35),
.B2(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_27),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_35),
.B1(n_12),
.B2(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_35),
.B1(n_37),
.B2(n_27),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_52),
.B(n_17),
.C(n_37),
.D(n_10),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_68),
.B(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_17),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_64),
.C(n_8),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_30),
.B(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_70),
.B1(n_27),
.B2(n_62),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_73),
.B(n_65),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_1),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_5),
.B(n_7),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_6),
.C(n_7),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_84),
.B1(n_81),
.B2(n_80),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_3),
.B(n_4),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_10),
.Y(n_86)
);


endmodule