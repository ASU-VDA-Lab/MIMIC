module fake_netlist_6_2827_n_2303 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2303);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2303;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_118),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_82),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_64),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_119),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_134),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_137),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_161),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_65),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_140),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_212),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_115),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_79),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_102),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_113),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_130),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_41),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_225),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_66),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_11),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_0),
.Y(n_256)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_111),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_168),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_13),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_93),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_65),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_23),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_110),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_148),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_122),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_80),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_81),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_6),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_146),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_97),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_133),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_29),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_178),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_126),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_75),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_105),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_151),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_27),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_132),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_63),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_46),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_206),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_173),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_125),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_7),
.Y(n_295)
);

INVx4_ASAP7_75t_R g296 ( 
.A(n_73),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_136),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_138),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_174),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_169),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_197),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_56),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_224),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_203),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_179),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_150),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_230),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_17),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_37),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_45),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_66),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_71),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_204),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_81),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_177),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_1),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_227),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_145),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_186),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_165),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_219),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_18),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_139),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_123),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_5),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_90),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_82),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_229),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_6),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_217),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_75),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_187),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_58),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_80),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_127),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_153),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_175),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_44),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_106),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_72),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_86),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_149),
.Y(n_345)
);

BUFx10_ASAP7_75t_L g346 ( 
.A(n_83),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_62),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_226),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_141),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_135),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_48),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_95),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_53),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_46),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_124),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_188),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_167),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_181),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_20),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_160),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_37),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_172),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_209),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_78),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_103),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_189),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_104),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_101),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_166),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_36),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_60),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_3),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_17),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_49),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_33),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_154),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_183),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_24),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_216),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_100),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_220),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_185),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_25),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_0),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_35),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_96),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_8),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_120),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_29),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_5),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_57),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_51),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_191),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_70),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_58),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_195),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_77),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_231),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_54),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_21),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_144),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_2),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_88),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_47),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_117),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_171),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_44),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_155),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_108),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_51),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_143),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_79),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_16),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_72),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_63),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_60),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_199),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_109),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_28),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_22),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_16),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_1),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_193),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_27),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_201),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_218),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_45),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_223),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_54),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_9),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_211),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_74),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_70),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_131),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_213),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_182),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_4),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_85),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_89),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_39),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_84),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_94),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_92),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_59),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_12),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_43),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_73),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_152),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_207),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_24),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_62),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_76),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_98),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_192),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_77),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_53),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_64),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_25),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_233),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_378),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_237),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_239),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_340),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_303),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_245),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_340),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_340),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_403),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_340),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_340),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_340),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_340),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_340),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_358),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_250),
.B(n_2),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_406),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_242),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_336),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_403),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_246),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_244),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_247),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_340),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_248),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_253),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_249),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_343),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_251),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_252),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_346),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_258),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_343),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_261),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_343),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_343),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_336),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_234),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_267),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_246),
.B(n_3),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_343),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_343),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_268),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_274),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_281),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_283),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_343),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_284),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_246),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_343),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_343),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_291),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_293),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_346),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_298),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_299),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g517 ( 
.A(n_241),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_300),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_265),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_346),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_428),
.B(n_7),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_250),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_304),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_307),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_308),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_315),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_447),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_319),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_320),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_321),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_236),
.B(n_8),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_271),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_271),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_309),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_309),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_265),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_347),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_235),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_452),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_322),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_236),
.B(n_9),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_452),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_455),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_323),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_347),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_325),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_292),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_360),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_347),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_458),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_326),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_334),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_256),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_238),
.B(n_10),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_337),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_348),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_R g562 ( 
.A(n_349),
.B(n_87),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_350),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_347),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_256),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_356),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_263),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_335),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_363),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_365),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_366),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_263),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_243),
.B(n_10),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_269),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_254),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_269),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_278),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_368),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_259),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_278),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_369),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_377),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_279),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_279),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_516),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_477),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_486),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_516),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_498),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_527),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_502),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_507),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_496),
.B(n_272),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_465),
.B(n_374),
.Y(n_595)
);

OA21x2_ASAP7_75t_L g596 ( 
.A1(n_559),
.A2(n_255),
.B(n_243),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_527),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_511),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_528),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_519),
.B(n_383),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_512),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_530),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_531),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_517),
.B(n_468),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_531),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_480),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_463),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_499),
.B(n_360),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_479),
.B(n_459),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_463),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_514),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_565),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_508),
.B(n_425),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_565),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_524),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_567),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_561),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_461),
.B(n_462),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_541),
.B(n_384),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_540),
.B(n_374),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_466),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_467),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_467),
.B(n_425),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_469),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_469),
.B(n_238),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_470),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_575),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_481),
.B(n_266),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_470),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_566),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_471),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_471),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_472),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_464),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_553),
.B(n_383),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_472),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_473),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_539),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_482),
.B(n_266),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_473),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_483),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_483),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_487),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_487),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_492),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_571),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_567),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_578),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_581),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_492),
.B(n_338),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_494),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_572),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_494),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_474),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_495),
.B(n_501),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_484),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_488),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_460),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_495),
.B(n_441),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_506),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_506),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_489),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_509),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_491),
.B(n_317),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_338),
.Y(n_671)
);

OA21x2_ASAP7_75t_L g672 ( 
.A1(n_509),
.A2(n_275),
.B(n_255),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_510),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_503),
.B(n_240),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_504),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_550),
.B(n_374),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_539),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_R g679 ( 
.A(n_505),
.B(n_380),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_476),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_515),
.B(n_342),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_628),
.B(n_633),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_594),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_624),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_609),
.Y(n_685)
);

INVx4_ASAP7_75t_SL g686 ( 
.A(n_664),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_613),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_611),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_675),
.B(n_518),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_611),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_664),
.B(n_441),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_660),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_628),
.B(n_342),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_678),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_613),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_660),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_644),
.B(n_523),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_664),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_628),
.B(n_441),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_671),
.B(n_525),
.Y(n_700)
);

BUFx4f_ASAP7_75t_L g701 ( 
.A(n_596),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_631),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_631),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_628),
.B(n_441),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_586),
.Y(n_705)
);

XNOR2xp5_ASAP7_75t_L g706 ( 
.A(n_624),
.B(n_552),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_681),
.B(n_441),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_616),
.B(n_526),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_616),
.B(n_529),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_678),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_588),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_611),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_660),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_612),
.B(n_532),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_660),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_623),
.B(n_475),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_664),
.B(n_275),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_616),
.B(n_533),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_616),
.B(n_611),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_605),
.B(n_564),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_594),
.B(n_579),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_631),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_622),
.B(n_543),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_600),
.B(n_548),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_631),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_630),
.B(n_655),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_626),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_631),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_673),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_630),
.B(n_551),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_607),
.A2(n_534),
.B1(n_573),
.B2(n_544),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_673),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_627),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_629),
.B(n_556),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_632),
.A2(n_395),
.B1(n_371),
.B2(n_485),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_634),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_632),
.A2(n_554),
.B1(n_521),
.B2(n_475),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_636),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_637),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_600),
.B(n_557),
.Y(n_743)
);

AND3x2_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_302),
.C(n_478),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_643),
.B(n_280),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_664),
.B(n_280),
.Y(n_746)
);

AND2x2_ASAP7_75t_SL g747 ( 
.A(n_596),
.B(n_286),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_664),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_640),
.B(n_560),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_643),
.B(n_286),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_640),
.B(n_563),
.Y(n_751)
);

XOR2xp5_ASAP7_75t_L g752 ( 
.A(n_639),
.B(n_568),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_630),
.B(n_569),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_592),
.B(n_570),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_586),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_659),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_625),
.A2(n_262),
.B1(n_264),
.B2(n_260),
.Y(n_758)
);

NOR2x1p5_ASAP7_75t_L g759 ( 
.A(n_662),
.B(n_385),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_670),
.B(n_582),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_604),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_673),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_673),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_673),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_641),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_638),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_642),
.B(n_510),
.Y(n_767)
);

INVx4_ASAP7_75t_SL g768 ( 
.A(n_664),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_662),
.B(n_490),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_595),
.B(n_513),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_647),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_641),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_643),
.B(n_297),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_649),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_650),
.B(n_277),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_658),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_668),
.B(n_520),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_668),
.B(n_522),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_667),
.B(n_287),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_676),
.B(n_677),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_643),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_679),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_669),
.B(n_294),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_643),
.B(n_297),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_648),
.B(n_306),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_619),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_676),
.B(n_584),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_619),
.Y(n_788)
);

BUFx8_ASAP7_75t_SL g789 ( 
.A(n_680),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_596),
.A2(n_272),
.B1(n_318),
.B2(n_385),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_648),
.B(n_339),
.Y(n_791)
);

INVxp33_ASAP7_75t_SL g792 ( 
.A(n_587),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_648),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_630),
.B(n_301),
.Y(n_794)
);

NAND3x1_ASAP7_75t_L g795 ( 
.A(n_608),
.B(n_289),
.C(n_285),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_587),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_645),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_645),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_608),
.B(n_574),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_666),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_655),
.B(n_301),
.Y(n_801)
);

XNOR2xp5_ASAP7_75t_L g802 ( 
.A(n_589),
.B(n_451),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_655),
.B(n_257),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_646),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_643),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_666),
.Y(n_806)
);

AND2x6_ASAP7_75t_L g807 ( 
.A(n_655),
.B(n_305),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_596),
.A2(n_273),
.B1(n_276),
.B2(n_270),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_589),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_656),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_666),
.B(n_305),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_656),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_610),
.B(n_574),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_665),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_610),
.Y(n_816)
);

NOR2x1p5_ASAP7_75t_L g817 ( 
.A(n_591),
.B(n_389),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_665),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_615),
.B(n_314),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_615),
.B(n_314),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_617),
.B(n_328),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_617),
.B(n_328),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_597),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_599),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_L g825 ( 
.A(n_620),
.B(n_330),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_620),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_652),
.B(n_657),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_674),
.B(n_576),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_652),
.B(n_330),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_585),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_585),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_657),
.B(n_332),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_SL g833 ( 
.A1(n_674),
.A2(n_318),
.B(n_332),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_585),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_602),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_603),
.B(n_344),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_606),
.B(n_396),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_590),
.B(n_341),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_590),
.B(n_576),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_585),
.B(n_398),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_585),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_672),
.B(n_257),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_591),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_692),
.A2(n_345),
.B(n_352),
.C(n_341),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_696),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_815),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_713),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_815),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_807),
.B(n_381),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_787),
.B(n_435),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_719),
.B(n_672),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_688),
.B(n_672),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_715),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_689),
.B(n_282),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_740),
.B(n_598),
.C(n_593),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_688),
.B(n_672),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_683),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_690),
.B(n_345),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_690),
.B(n_712),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_712),
.B(n_701),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_684),
.B(n_721),
.Y(n_861)
);

NOR3xp33_ASAP7_75t_L g862 ( 
.A(n_738),
.B(n_598),
.C(n_593),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_701),
.B(n_747),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_725),
.B(n_601),
.Y(n_864)
);

INVx5_ASAP7_75t_L g865 ( 
.A(n_842),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_682),
.B(n_352),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_716),
.B(n_601),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_682),
.B(n_785),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_791),
.B(n_355),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_759),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_716),
.A2(n_409),
.B1(n_382),
.B2(n_453),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_714),
.B(n_288),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_728),
.B(n_355),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_816),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_828),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_685),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_778),
.B(n_618),
.C(n_614),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_736),
.B(n_357),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_701),
.B(n_386),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_694),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_743),
.B(n_614),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_739),
.B(n_357),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_SL g883 ( 
.A1(n_780),
.A2(n_654),
.B1(n_653),
.B2(n_651),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_741),
.B(n_362),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_749),
.B(n_751),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_821),
.A2(n_822),
.B(n_832),
.C(n_829),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_742),
.B(n_362),
.Y(n_887)
);

INVx8_ASAP7_75t_L g888 ( 
.A(n_803),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_726),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_777),
.B(n_618),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_747),
.B(n_393),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_799),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_758),
.B(n_635),
.C(n_621),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_814),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_769),
.B(n_621),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_716),
.B(n_635),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_766),
.B(n_367),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_817),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_716),
.B(n_697),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_708),
.A2(n_418),
.B1(n_438),
.B2(n_436),
.Y(n_900)
);

OAI22xp33_ASAP7_75t_L g901 ( 
.A1(n_700),
.A2(n_427),
.B1(n_421),
.B2(n_389),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_694),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_839),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_808),
.B(n_401),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_687),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_771),
.B(n_367),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_793),
.B(n_411),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_760),
.B(n_651),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_727),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

OAI22xp33_ASAP7_75t_L g911 ( 
.A1(n_803),
.A2(n_427),
.B1(n_421),
.B2(n_313),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_826),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_774),
.B(n_376),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_776),
.B(n_376),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_827),
.B(n_379),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_695),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_840),
.B(n_379),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_800),
.B(n_388),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_L g920 ( 
.A(n_708),
.B(n_654),
.C(n_653),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_709),
.A2(n_718),
.B1(n_753),
.B2(n_733),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_782),
.B(n_562),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_789),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_806),
.B(n_388),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_734),
.A2(n_405),
.B1(n_408),
.B2(n_439),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_710),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_733),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_720),
.B(n_417),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_695),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_765),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_770),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_752),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_724),
.B(n_295),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_711),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_765),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_823),
.B(n_824),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_790),
.A2(n_426),
.B(n_405),
.C(n_408),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_835),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_772),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_709),
.A2(n_423),
.B1(n_426),
.B2(n_431),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_431),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_698),
.B(n_434),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_753),
.B(n_577),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_754),
.B(n_374),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_779),
.B(n_434),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_718),
.B(n_311),
.C(n_310),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_698),
.B(n_439),
.Y(n_947)
);

AO221x1_ASAP7_75t_L g948 ( 
.A1(n_702),
.A2(n_290),
.B1(n_457),
.B2(n_285),
.C(n_289),
.Y(n_948)
);

NAND3xp33_ASAP7_75t_L g949 ( 
.A(n_783),
.B(n_324),
.C(n_316),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_737),
.B(n_327),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_807),
.B(n_442),
.Y(n_951)
);

OAI22xp33_ASAP7_75t_SL g952 ( 
.A1(n_707),
.A2(n_442),
.B1(n_443),
.B2(n_448),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_698),
.B(n_443),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_707),
.B(n_448),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_786),
.B(n_449),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_836),
.B(n_449),
.Y(n_956)
);

INVx8_ASAP7_75t_L g957 ( 
.A(n_803),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_788),
.B(n_454),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_711),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_837),
.B(n_329),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_803),
.B(n_333),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_706),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_767),
.B(n_351),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_693),
.B(n_354),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_SL g965 ( 
.A(n_722),
.B(n_359),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_744),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_794),
.Y(n_967)
);

INVx8_ASAP7_75t_L g968 ( 
.A(n_807),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_702),
.B(n_454),
.Y(n_969)
);

OAI22xp33_ASAP7_75t_L g970 ( 
.A1(n_842),
.A2(n_290),
.B1(n_312),
.B2(n_313),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_794),
.B(n_420),
.C(n_399),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_698),
.B(n_361),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_722),
.B(n_577),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_702),
.B(n_580),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_693),
.B(n_364),
.Y(n_975)
);

AND3x1_ASAP7_75t_L g976 ( 
.A(n_795),
.B(n_312),
.C(n_404),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_703),
.B(n_580),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_698),
.B(n_372),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_729),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_703),
.B(n_583),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_703),
.B(n_583),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_842),
.B(n_801),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_833),
.A2(n_353),
.B(n_404),
.C(n_424),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_763),
.B(n_584),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_726),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_726),
.Y(n_986)
);

O2A1O1Ixp5_ASAP7_75t_L g987 ( 
.A1(n_699),
.A2(n_704),
.B(n_801),
.C(n_829),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_748),
.B(n_373),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_763),
.B(n_390),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_802),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_748),
.B(n_394),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_797),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_748),
.B(n_797),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_789),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_798),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_842),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_763),
.B(n_764),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_732),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_748),
.B(n_397),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_798),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_756),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_748),
.B(n_400),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_821),
.B(n_822),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_832),
.B(n_402),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_812),
.A2(n_446),
.B1(n_331),
.B2(n_353),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_764),
.B(n_414),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_L g1007 ( 
.A(n_807),
.B(n_812),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_804),
.B(n_415),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_699),
.B(n_416),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_764),
.B(n_419),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_804),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_809),
.B(n_422),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_925),
.A2(n_820),
.B(n_825),
.C(n_819),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_973),
.B(n_722),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_885),
.A2(n_807),
.B1(n_812),
.B2(n_704),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_970),
.A2(n_820),
.B(n_825),
.C(n_819),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_889),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_845),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_859),
.A2(n_730),
.B(n_723),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_851),
.A2(n_730),
.B(n_723),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_868),
.A2(n_730),
.B(n_723),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_865),
.B(n_731),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_872),
.A2(n_391),
.B(n_331),
.C(n_440),
.Y(n_1023)
);

AOI33xp33_ASAP7_75t_L g1024 ( 
.A1(n_874),
.A2(n_446),
.A3(n_370),
.B1(n_375),
.B2(n_387),
.B3(n_391),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_921),
.A2(n_843),
.B1(n_810),
.B2(n_796),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_865),
.B(n_731),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_845),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_847),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_889),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_852),
.A2(n_813),
.B(n_811),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_1001),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_856),
.A2(n_762),
.B(n_735),
.Y(n_1032)
);

OAI321xp33_ASAP7_75t_L g1033 ( 
.A1(n_901),
.A2(n_440),
.A3(n_370),
.B1(n_375),
.B2(n_387),
.C(n_392),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_854),
.B(n_811),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_885),
.B(n_731),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_860),
.A2(n_735),
.B(n_762),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_853),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_865),
.B(n_732),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_959),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_854),
.B(n_813),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_889),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_879),
.A2(n_818),
.B(n_750),
.C(n_773),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_970),
.A2(n_838),
.B(n_717),
.C(n_746),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_979),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_987),
.A2(n_818),
.B(n_812),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_850),
.B(n_705),
.C(n_838),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_865),
.B(n_732),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_879),
.A2(n_841),
.B(n_729),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_850),
.B(n_792),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_863),
.B(n_732),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_863),
.A2(n_812),
.B(n_735),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_963),
.B(n_830),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_860),
.A2(n_762),
.B(n_757),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_861),
.B(n_899),
.Y(n_1054)
);

OAI321xp33_ASAP7_75t_L g1055 ( 
.A1(n_901),
.A2(n_940),
.A3(n_911),
.B1(n_1004),
.B2(n_904),
.C(n_996),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_891),
.A2(n_429),
.B1(n_392),
.B2(n_457),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_933),
.B(n_830),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_899),
.A2(n_773),
.B1(n_750),
.B2(n_745),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_876),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_938),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_982),
.A2(n_757),
.B(n_761),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_982),
.A2(n_761),
.B(n_746),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_933),
.B(n_745),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_950),
.B(n_745),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_950),
.B(n_750),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_888),
.B(n_795),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_997),
.A2(n_834),
.B(n_781),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_960),
.B(n_773),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_960),
.B(n_784),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_846),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_888),
.B(n_792),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_944),
.B(n_755),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_SL g1073 ( 
.A1(n_965),
.A2(n_705),
.B1(n_756),
.B2(n_407),
.Y(n_1073)
);

AND2x4_ASAP7_75t_SL g1074 ( 
.A(n_943),
.B(n_784),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1007),
.A2(n_834),
.B(n_781),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_917),
.A2(n_805),
.B(n_781),
.Y(n_1076)
);

AND2x2_ASAP7_75t_SL g1077 ( 
.A(n_1005),
.B(n_717),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_917),
.A2(n_805),
.B(n_831),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_927),
.B(n_430),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_848),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_857),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_998),
.A2(n_831),
.B(n_691),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_926),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_866),
.A2(n_831),
.B(n_691),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_930),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_909),
.A2(n_910),
.B(n_936),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_967),
.B(n_1003),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1003),
.A2(n_784),
.B(n_424),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_889),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_891),
.A2(n_456),
.B1(n_450),
.B2(n_445),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_886),
.A2(n_429),
.B(n_437),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_993),
.A2(n_831),
.B(n_768),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_985),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_935),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_876),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_993),
.A2(n_768),
.B(n_686),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1004),
.A2(n_407),
.B(n_437),
.C(n_432),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_943),
.B(n_686),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_985),
.A2(n_986),
.B(n_858),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_926),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_892),
.B(n_894),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_939),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_985),
.A2(n_768),
.B(n_686),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_903),
.B(n_985),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_986),
.A2(n_555),
.B(n_549),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_875),
.B(n_535),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_994),
.B(n_91),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_986),
.A2(n_555),
.B(n_549),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_912),
.B(n_433),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_986),
.A2(n_547),
.B(n_546),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_992),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_934),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_968),
.A2(n_547),
.B(n_546),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_962),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_904),
.A2(n_915),
.B(n_937),
.C(n_918),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_888),
.A2(n_444),
.B1(n_542),
.B2(n_538),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_968),
.A2(n_545),
.B(n_542),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_869),
.B(n_535),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_964),
.A2(n_545),
.B(n_538),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_871),
.B(n_536),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_880),
.B(n_536),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_968),
.A2(n_1006),
.B(n_989),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_908),
.B(n_11),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1010),
.A2(n_951),
.B(n_849),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_880),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_964),
.B(n_537),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_995),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1000),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_902),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_975),
.A2(n_1009),
.B(n_1011),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_975),
.B(n_537),
.Y(n_1131)
);

OAI321xp33_ASAP7_75t_L g1132 ( 
.A1(n_911),
.A2(n_296),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_18),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_941),
.B(n_12),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_L g1134 ( 
.A(n_922),
.B(n_99),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1009),
.A2(n_232),
.B(n_222),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_907),
.A2(n_221),
.B(n_214),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_934),
.B(n_208),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_945),
.B(n_974),
.Y(n_1138)
);

OR2x6_ASAP7_75t_SL g1139 ( 
.A(n_923),
.B(n_14),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_957),
.A2(n_202),
.B1(n_200),
.B2(n_198),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_977),
.B(n_15),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_895),
.B(n_19),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_957),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_946),
.B(n_196),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_907),
.A2(n_190),
.B(n_184),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_864),
.B(n_19),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_961),
.A2(n_20),
.B(n_21),
.C(n_26),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_898),
.Y(n_1148)
);

AOI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_961),
.A2(n_26),
.B(n_28),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_969),
.A2(n_164),
.B(n_163),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1012),
.A2(n_159),
.B(n_158),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_870),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_905),
.A2(n_157),
.B(n_156),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_966),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_980),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_981),
.B(n_31),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_984),
.B(n_32),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_873),
.B(n_32),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_881),
.B(n_867),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_916),
.A2(n_147),
.B(n_142),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_929),
.B(n_129),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_919),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_955),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_972),
.A2(n_128),
.B(n_121),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_972),
.A2(n_116),
.B(n_114),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1008),
.A2(n_112),
.B1(n_107),
.B2(n_35),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_978),
.A2(n_33),
.B(n_34),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_978),
.A2(n_34),
.B(n_36),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_988),
.A2(n_991),
.B(n_999),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_844),
.A2(n_956),
.B(n_1008),
.C(n_983),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_957),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_958),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_878),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_882),
.B(n_38),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_988),
.A2(n_40),
.B(n_42),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_942),
.B(n_42),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_884),
.B(n_43),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_924),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_991),
.A2(n_47),
.B(n_48),
.Y(n_1179)
);

NOR2x1_ASAP7_75t_L g1180 ( 
.A(n_890),
.B(n_49),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_887),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_883),
.B(n_50),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_897),
.B(n_50),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_999),
.A2(n_52),
.B(n_55),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1005),
.A2(n_83),
.B1(n_55),
.B2(n_57),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_954),
.A2(n_52),
.B(n_59),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1002),
.A2(n_61),
.B(n_67),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_932),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_952),
.B(n_949),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_906),
.B(n_61),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1002),
.A2(n_947),
.B(n_953),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_931),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_971),
.B(n_67),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_896),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_900),
.B(n_913),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_928),
.B(n_68),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_942),
.A2(n_68),
.B(n_69),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_947),
.A2(n_69),
.B(n_71),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_953),
.A2(n_74),
.B(n_76),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_914),
.A2(n_78),
.B(n_948),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_931),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_976),
.B(n_893),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1028),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1072),
.B(n_877),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1083),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1186),
.A2(n_920),
.B(n_855),
.C(n_862),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1031),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1041),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1124),
.A2(n_990),
.B(n_1063),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1041),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1050),
.A2(n_1048),
.B(n_1052),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_1020),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1036),
.A2(n_1053),
.B(n_1122),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1087),
.B(n_1181),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1030),
.A2(n_1050),
.B(n_1169),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1014),
.B(n_1054),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1068),
.A2(n_1069),
.B(n_1057),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1049),
.A2(n_1035),
.B1(n_1054),
.B2(n_1159),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1081),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1049),
.B(n_1178),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1041),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1163),
.B(n_1172),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1192),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1041),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1021),
.A2(n_1051),
.B(n_1032),
.Y(n_1225)
);

BUFx2_ASAP7_75t_SL g1226 ( 
.A(n_1100),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_L g1227 ( 
.A1(n_1195),
.A2(n_1189),
.B(n_1130),
.C(n_1144),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1035),
.B(n_1143),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1115),
.A2(n_1062),
.B(n_1086),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1075),
.A2(n_1099),
.B(n_1061),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1018),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1037),
.Y(n_1232)
);

NAND2x1_ASAP7_75t_L g1233 ( 
.A(n_1017),
.B(n_1029),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1125),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1018),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1015),
.A2(n_1040),
.B1(n_1034),
.B2(n_1056),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1017),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1055),
.B(n_1046),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1195),
.A2(n_1191),
.B(n_1088),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1104),
.A2(n_1019),
.B(n_1038),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1162),
.B(n_1138),
.Y(n_1241)
);

AOI21xp33_ASAP7_75t_L g1242 ( 
.A1(n_1159),
.A2(n_1196),
.B(n_1079),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1083),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1121),
.B(n_1109),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1098),
.A2(n_1047),
.B(n_1038),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1067),
.A2(n_1150),
.B(n_1084),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1196),
.B(n_1146),
.C(n_1123),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1081),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_1114),
.B(n_1188),
.Y(n_1249)
);

CKINVDCx8_ASAP7_75t_R g1250 ( 
.A(n_1201),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1091),
.A2(n_1082),
.B(n_1092),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1060),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1155),
.B(n_1126),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1027),
.Y(n_1254)
);

OAI21xp33_ASAP7_75t_L g1255 ( 
.A1(n_1109),
.A2(n_1146),
.B(n_1123),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1135),
.A2(n_1153),
.B(n_1016),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1059),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1095),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1106),
.B(n_1079),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1131),
.B(n_1101),
.Y(n_1260)
);

INVx5_ASAP7_75t_L g1261 ( 
.A(n_1029),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1161),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1039),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1149),
.A2(n_1097),
.B(n_1147),
.C(n_1023),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1044),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1266)
);

OAI21xp33_ASAP7_75t_L g1267 ( 
.A1(n_1073),
.A2(n_1097),
.B(n_1182),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1077),
.B(n_1133),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1013),
.A2(n_1132),
.B(n_1077),
.C(n_1043),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1197),
.A2(n_1199),
.B(n_1184),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1161),
.A2(n_1137),
.B(n_1165),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1202),
.A2(n_1194),
.B1(n_1025),
.B2(n_1142),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1070),
.B(n_1080),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1023),
.A2(n_1147),
.A3(n_1200),
.B(n_1141),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1085),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1129),
.B(n_1158),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1137),
.A2(n_1164),
.B(n_1170),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1033),
.A2(n_1024),
.B(n_1193),
.C(n_1185),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1171),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1134),
.B(n_1058),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1171),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1129),
.B(n_1177),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1148),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1160),
.A2(n_1103),
.B(n_1151),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1096),
.A2(n_1144),
.B(n_1189),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1024),
.A2(n_1193),
.B(n_1167),
.C(n_1187),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1125),
.B(n_1152),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1094),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1026),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1136),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1174),
.B(n_1190),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1180),
.B(n_1071),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1168),
.A2(n_1179),
.B(n_1175),
.C(n_1173),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1128),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1102),
.Y(n_1296)
);

NAND2x1_ASAP7_75t_L g1297 ( 
.A(n_1112),
.B(n_1127),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1022),
.A2(n_1026),
.B(n_1117),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1111),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1145),
.A2(n_1113),
.B(n_1022),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1090),
.A2(n_1120),
.B(n_1183),
.C(n_1116),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1120),
.A2(n_1119),
.B(n_1118),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1118),
.Y(n_1303)
);

NOR2x1_ASAP7_75t_SL g1304 ( 
.A(n_1071),
.B(n_1066),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1166),
.A2(n_1066),
.B1(n_1176),
.B2(n_1071),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1176),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1198),
.A2(n_1140),
.A3(n_1105),
.B(n_1108),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1110),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1107),
.B(n_1066),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1139),
.A2(n_1048),
.B(n_1045),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1143),
.B(n_1171),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1115),
.A2(n_863),
.B(n_701),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1049),
.A2(n_1073),
.B(n_872),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1071),
.B(n_888),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1072),
.B(n_1014),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1050),
.A2(n_860),
.B(n_879),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1048),
.A2(n_1045),
.B(n_1042),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1049),
.B(n_872),
.C(n_850),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1186),
.A2(n_1077),
.B1(n_1185),
.B2(n_1149),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1087),
.B(n_872),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1048),
.A2(n_1045),
.B(n_1042),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1115),
.A2(n_863),
.B(n_701),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1087),
.B(n_872),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1115),
.A2(n_863),
.B(n_701),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_SL g1325 ( 
.A(n_1049),
.B(n_872),
.C(n_705),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1048),
.A2(n_1045),
.B(n_1042),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1124),
.A2(n_863),
.B(n_860),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1087),
.B(n_872),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1072),
.B(n_1014),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1083),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1048),
.A2(n_1045),
.B(n_1042),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1115),
.A2(n_863),
.B(n_701),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1041),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1072),
.B(n_1014),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1087),
.B(n_872),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1087),
.B(n_872),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1087),
.B(n_872),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1041),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1124),
.A2(n_863),
.B(n_860),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1186),
.A2(n_1016),
.B(n_1013),
.C(n_1196),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1087),
.B(n_872),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1124),
.A2(n_863),
.B(n_860),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1049),
.A2(n_872),
.B(n_850),
.Y(n_1343)
);

AOI221x1_ASAP7_75t_L g1344 ( 
.A1(n_1200),
.A2(n_1186),
.B1(n_1097),
.B2(n_1202),
.C(n_925),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1048),
.A2(n_1045),
.B(n_1042),
.Y(n_1345)
);

AND2x2_ASAP7_75t_SL g1346 ( 
.A(n_1077),
.B(n_1056),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1041),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1087),
.B(n_872),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1087),
.B(n_872),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1041),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1048),
.A2(n_1045),
.B(n_1042),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1087),
.B(n_872),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1041),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1087),
.B(n_872),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1124),
.A2(n_863),
.B(n_860),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1125),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1091),
.A2(n_1061),
.B(n_1045),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1087),
.B(n_872),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1115),
.A2(n_863),
.B(n_701),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1083),
.Y(n_1360)
);

AOI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1202),
.A2(n_1142),
.B(n_1158),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1115),
.A2(n_863),
.B(n_701),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1087),
.B(n_872),
.Y(n_1363)
);

AOI21xp33_ASAP7_75t_L g1364 ( 
.A1(n_1049),
.A2(n_872),
.B(n_854),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1287),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1241),
.B(n_1320),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1203),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1232),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1216),
.B(n_1315),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1243),
.Y(n_1370)
);

INVx3_ASAP7_75t_SL g1371 ( 
.A(n_1207),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1343),
.A2(n_1313),
.B1(n_1318),
.B2(n_1255),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1329),
.B(n_1334),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1364),
.A2(n_1247),
.B(n_1242),
.C(n_1301),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1244),
.B(n_1259),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1234),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1234),
.B(n_1356),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1325),
.A2(n_1204),
.B1(n_1218),
.B2(n_1267),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1220),
.B(n_1323),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1346),
.A2(n_1319),
.B1(n_1238),
.B2(n_1256),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1279),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1330),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1328),
.B(n_1335),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_SL g1384 ( 
.A1(n_1239),
.A2(n_1229),
.B(n_1319),
.C(n_1209),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1346),
.A2(n_1305),
.B1(n_1349),
.B2(n_1348),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1248),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1356),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1226),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1252),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1248),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1341),
.B(n_1352),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1340),
.A2(n_1227),
.B(n_1269),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1207),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1249),
.A2(n_1363),
.B1(n_1354),
.B2(n_1358),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1360),
.B(n_1222),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1360),
.B(n_1293),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1260),
.B(n_1253),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_1219),
.Y(n_1399)
);

INVx5_ASAP7_75t_L g1400 ( 
.A(n_1350),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1214),
.B(n_1276),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1225),
.A2(n_1362),
.B(n_1359),
.Y(n_1402)
);

NOR2xp67_ASAP7_75t_L g1403 ( 
.A(n_1272),
.B(n_1205),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1263),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1291),
.B(n_1268),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1314),
.B(n_1292),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1269),
.B(n_1340),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1238),
.A2(n_1206),
.B(n_1264),
.C(n_1278),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1206),
.B(n_1275),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1279),
.Y(n_1411)
);

INVx5_ASAP7_75t_L g1412 ( 
.A(n_1350),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1279),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1223),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1350),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1344),
.B(n_1286),
.C(n_1294),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1273),
.B(n_1265),
.Y(n_1417)
);

INVx3_ASAP7_75t_SL g1418 ( 
.A(n_1223),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1236),
.B(n_1278),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1288),
.B(n_1296),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1279),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1254),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1314),
.B(n_1304),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1231),
.B(n_1254),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1281),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1231),
.B(n_1299),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1261),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1312),
.A2(n_1332),
.B(n_1322),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1299),
.B(n_1303),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1324),
.A2(n_1342),
.B(n_1355),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1314),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1250),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1266),
.A2(n_1306),
.B1(n_1280),
.B2(n_1309),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1327),
.A2(n_1339),
.B(n_1357),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1306),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1280),
.A2(n_1309),
.B1(n_1235),
.B2(n_1258),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1250),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1257),
.Y(n_1438)
);

AOI21xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1310),
.A2(n_1286),
.B(n_1311),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1357),
.A2(n_1285),
.B(n_1302),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1357),
.A2(n_1213),
.B(n_1230),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_SL g1443 ( 
.A(n_1228),
.B(n_1261),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1281),
.B(n_1261),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1213),
.A2(n_1230),
.B(n_1277),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1208),
.Y(n_1446)
);

NAND2x1p5_ASAP7_75t_L g1447 ( 
.A(n_1261),
.B(n_1353),
.Y(n_1447)
);

INVx5_ASAP7_75t_L g1448 ( 
.A(n_1350),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1353),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1208),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1235),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1281),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1277),
.A2(n_1295),
.B(n_1251),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1311),
.A2(n_1281),
.B1(n_1338),
.B2(n_1233),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1237),
.B(n_1353),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1310),
.A2(n_1308),
.B1(n_1270),
.B2(n_1297),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1210),
.Y(n_1457)
);

CKINVDCx8_ASAP7_75t_R g1458 ( 
.A(n_1353),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1274),
.B(n_1210),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1251),
.A2(n_1215),
.B(n_1308),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1221),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1237),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1221),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1338),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1224),
.Y(n_1465)
);

O2A1O1Ixp5_ASAP7_75t_L g1466 ( 
.A1(n_1294),
.A2(n_1316),
.B(n_1240),
.C(n_1211),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1274),
.B(n_1333),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1298),
.A2(n_1245),
.B(n_1289),
.C(n_1224),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1333),
.A2(n_1347),
.B1(n_1274),
.B2(n_1361),
.Y(n_1469)
);

INVx8_ASAP7_75t_L g1470 ( 
.A(n_1347),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1274),
.B(n_1215),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1290),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1307),
.A2(n_1271),
.B1(n_1300),
.B2(n_1351),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1290),
.B(n_1262),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1307),
.B(n_1271),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1307),
.B(n_1321),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1300),
.Y(n_1477)
);

BUFx2_ASAP7_75t_SL g1478 ( 
.A(n_1307),
.Y(n_1478)
);

NAND2xp33_ASAP7_75t_L g1479 ( 
.A(n_1262),
.B(n_1284),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1317),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1351),
.B(n_1326),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1246),
.B(n_1345),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1331),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1212),
.A2(n_1217),
.B(n_1229),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1241),
.B(n_1320),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1234),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1243),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1279),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1241),
.B(n_1320),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1248),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1207),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1241),
.B(n_1320),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1346),
.A2(n_1319),
.B1(n_1247),
.B2(n_1269),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1223),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1207),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1234),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1234),
.B(n_1143),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1279),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1243),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1207),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1287),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1261),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1279),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1287),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1243),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1212),
.A2(n_1217),
.B(n_1229),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1313),
.A2(n_706),
.B(n_1049),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1346),
.A2(n_1319),
.B1(n_1247),
.B2(n_1269),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1364),
.B(n_1343),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1216),
.B(n_1315),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_SL g1512 ( 
.A(n_1314),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1364),
.B(n_1318),
.C(n_1343),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1226),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1340),
.A2(n_1227),
.B(n_1269),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1346),
.A2(n_1319),
.B1(n_1247),
.B2(n_1269),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1203),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1216),
.B(n_1315),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_SL g1519 ( 
.A(n_1234),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1241),
.B(n_1320),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1203),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1279),
.Y(n_1522)
);

AO22x1_ASAP7_75t_L g1523 ( 
.A1(n_1220),
.A2(n_1049),
.B1(n_780),
.B2(n_1035),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1360),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1203),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1346),
.A2(n_1319),
.B1(n_1247),
.B2(n_1269),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1241),
.B(n_1320),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1234),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1287),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1203),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1207),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1314),
.B(n_1226),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1234),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1364),
.A2(n_1343),
.B1(n_1318),
.B2(n_1255),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1445),
.A2(n_1460),
.B(n_1466),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1398),
.A2(n_1395),
.B1(n_1508),
.B2(n_1378),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1494),
.A2(n_1516),
.B1(n_1526),
.B2(n_1509),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1466),
.A2(n_1402),
.B(n_1485),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1398),
.A2(n_1372),
.B1(n_1385),
.B2(n_1534),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1449),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1420),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1523),
.B(n_1510),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1367),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1441),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1368),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1386),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1432),
.A2(n_1388),
.B1(n_1514),
.B2(n_1495),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1449),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1494),
.A2(n_1516),
.B1(n_1509),
.B2(n_1526),
.Y(n_1549)
);

NAND2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1449),
.B(n_1427),
.Y(n_1550)
);

BUFx8_ASAP7_75t_L g1551 ( 
.A(n_1519),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_SL g1552 ( 
.A(n_1414),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1438),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1377),
.Y(n_1554)
);

BUFx2_ASAP7_75t_R g1555 ( 
.A(n_1418),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1369),
.B(n_1511),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1383),
.B(n_1379),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1390),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1404),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1377),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1449),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1517),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1383),
.B(n_1389),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1407),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1366),
.A2(n_1527),
.B1(n_1490),
.B2(n_1486),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1401),
.B(n_1518),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1525),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1513),
.A2(n_1380),
.B1(n_1515),
.B2(n_1393),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1366),
.A2(n_1490),
.B1(n_1527),
.B2(n_1486),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1370),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1393),
.A2(n_1515),
.B1(n_1419),
.B2(n_1408),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1402),
.A2(n_1485),
.B(n_1507),
.Y(n_1573)
);

AO22x1_ASAP7_75t_L g1574 ( 
.A1(n_1392),
.A2(n_1520),
.B1(n_1493),
.B2(n_1423),
.Y(n_1574)
);

BUFx12f_ASAP7_75t_L g1575 ( 
.A(n_1437),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1408),
.A2(n_1443),
.B1(n_1419),
.B2(n_1405),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1442),
.A2(n_1434),
.B(n_1468),
.Y(n_1577)
);

INVx6_ASAP7_75t_L g1578 ( 
.A(n_1399),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1530),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1493),
.B(n_1520),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1403),
.A2(n_1433),
.B1(n_1374),
.B2(n_1405),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1417),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1396),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1375),
.A2(n_1373),
.B1(n_1410),
.B2(n_1423),
.Y(n_1584)
);

CKINVDCx11_ASAP7_75t_R g1585 ( 
.A(n_1531),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1416),
.A2(n_1428),
.B1(n_1397),
.B2(n_1491),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1428),
.A2(n_1391),
.B1(n_1431),
.B2(n_1512),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1468),
.A2(n_1430),
.B(n_1440),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1451),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1382),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1488),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1427),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1529),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1500),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1376),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1365),
.B(n_1502),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1376),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1506),
.A2(n_1524),
.B1(n_1429),
.B2(n_1435),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1429),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1394),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1505),
.A2(n_1532),
.B1(n_1436),
.B2(n_1464),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1503),
.B(n_1400),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1424),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1465),
.B(n_1533),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1376),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1424),
.Y(n_1606)
);

AO21x1_ASAP7_75t_L g1607 ( 
.A1(n_1409),
.A2(n_1469),
.B(n_1439),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1487),
.B(n_1533),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1503),
.A2(n_1447),
.B(n_1409),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1440),
.A2(n_1453),
.B(n_1472),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1463),
.Y(n_1611)
);

NAND2x1p5_ASAP7_75t_L g1612 ( 
.A(n_1400),
.B(n_1412),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1532),
.A2(n_1406),
.B1(n_1478),
.B2(n_1459),
.Y(n_1613)
);

AO21x2_ASAP7_75t_L g1614 ( 
.A1(n_1473),
.A2(n_1479),
.B(n_1384),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1426),
.B(n_1387),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1475),
.A2(n_1476),
.B(n_1471),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1426),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1400),
.Y(n_1618)
);

INVx5_ASAP7_75t_SL g1619 ( 
.A(n_1487),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1475),
.A2(n_1482),
.B(n_1481),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1447),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1492),
.Y(n_1622)
);

BUFx4f_ASAP7_75t_SL g1623 ( 
.A(n_1487),
.Y(n_1623)
);

AO21x1_ASAP7_75t_SL g1624 ( 
.A1(n_1467),
.A2(n_1456),
.B(n_1476),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1467),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1497),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1497),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1446),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1450),
.Y(n_1629)
);

CKINVDCx11_ASAP7_75t_R g1630 ( 
.A(n_1371),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1457),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1532),
.A2(n_1406),
.B1(n_1484),
.B2(n_1469),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1406),
.A2(n_1519),
.B1(n_1471),
.B2(n_1480),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1497),
.B(n_1533),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1528),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1462),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1415),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1461),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1455),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1483),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1444),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1400),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1444),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1461),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1528),
.B(n_1498),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1461),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1458),
.A2(n_1498),
.B1(n_1454),
.B2(n_1528),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1455),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1381),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1477),
.A2(n_1483),
.B1(n_1522),
.B2(n_1411),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1474),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1381),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1411),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1496),
.A2(n_1501),
.B1(n_1399),
.B2(n_1452),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1412),
.B(n_1448),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1489),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1474),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1412),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1499),
.A2(n_1504),
.B1(n_1421),
.B2(n_1425),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1413),
.A2(n_1448),
.B(n_1470),
.Y(n_1660)
);

BUFx2_ASAP7_75t_R g1661 ( 
.A(n_1470),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1470),
.A2(n_1255),
.B1(n_1247),
.B2(n_1343),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1448),
.A2(n_1246),
.B(n_1445),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1448),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1376),
.Y(n_1665)
);

AO21x1_ASAP7_75t_L g1666 ( 
.A1(n_1494),
.A2(n_1364),
.B(n_1313),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1423),
.B(n_1406),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1398),
.A2(n_1218),
.B1(n_1318),
.B2(n_1049),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1389),
.B(n_1392),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1529),
.Y(n_1670)
);

OAI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1508),
.A2(n_1313),
.B1(n_1318),
.B2(n_1218),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1494),
.A2(n_1318),
.B1(n_1049),
.B2(n_780),
.Y(n_1672)
);

CKINVDCx16_ASAP7_75t_R g1673 ( 
.A(n_1495),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1420),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1369),
.B(n_1511),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1445),
.A2(n_1246),
.B(n_1262),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1420),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1369),
.B(n_1511),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1420),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1420),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1386),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1420),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1376),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1420),
.Y(n_1684)
);

AND2x6_ASAP7_75t_L g1685 ( 
.A(n_1459),
.B(n_1408),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1420),
.Y(n_1686)
);

BUFx10_ASAP7_75t_L g1687 ( 
.A(n_1519),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1376),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1510),
.A2(n_1255),
.B1(n_1247),
.B2(n_1343),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1445),
.A2(n_1246),
.B(n_1262),
.Y(n_1690)
);

CKINVDCx11_ASAP7_75t_R g1691 ( 
.A(n_1495),
.Y(n_1691)
);

INVx6_ASAP7_75t_L g1692 ( 
.A(n_1449),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1376),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1449),
.Y(n_1694)
);

BUFx8_ASAP7_75t_L g1695 ( 
.A(n_1519),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1386),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1423),
.B(n_1406),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1420),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1437),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1495),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1510),
.A2(n_1255),
.B1(n_1247),
.B2(n_1343),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1422),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1420),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1510),
.A2(n_1255),
.B1(n_1247),
.B2(n_1343),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1422),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1386),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1386),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1420),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1377),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1420),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1407),
.Y(n_1711)
);

OAI22x1_ASAP7_75t_L g1712 ( 
.A1(n_1378),
.A2(n_1247),
.B1(n_1372),
.B2(n_1218),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1407),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_SL g1714 ( 
.A(n_1377),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1581),
.A2(n_1655),
.B(n_1612),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1640),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1672),
.A2(n_1549),
.B1(n_1537),
.B2(n_1689),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1557),
.B(n_1564),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1676),
.A2(n_1690),
.B(n_1610),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1625),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1616),
.B(n_1549),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1569),
.B(n_1544),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1616),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1620),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1620),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1546),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1668),
.A2(n_1671),
.B(n_1689),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1569),
.B(n_1544),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1667),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1553),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1657),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1572),
.B(n_1586),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1557),
.B(n_1564),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1681),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1685),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1607),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1642),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1663),
.A2(n_1535),
.B(n_1577),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1617),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1696),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1573),
.Y(n_1742)
);

INVxp33_ASAP7_75t_L g1743 ( 
.A(n_1556),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1612),
.A2(n_1655),
.B(n_1576),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1667),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1586),
.B(n_1573),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1614),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1660),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1706),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1538),
.Y(n_1751)
);

AND2x4_ASAP7_75t_SL g1752 ( 
.A(n_1667),
.B(n_1697),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1614),
.Y(n_1753)
);

CKINVDCx6p67_ASAP7_75t_R g1754 ( 
.A(n_1575),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1701),
.A2(n_1704),
.B(n_1542),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1589),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1538),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1572),
.B(n_1624),
.Y(n_1758)
);

OA21x2_ASAP7_75t_L g1759 ( 
.A1(n_1588),
.A2(n_1666),
.B(n_1650),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1685),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1567),
.B(n_1675),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1650),
.A2(n_1632),
.B(n_1542),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1685),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1566),
.A2(n_1570),
.B(n_1539),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1707),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1613),
.A2(n_1609),
.B(n_1633),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1685),
.B(n_1599),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1685),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1697),
.B(n_1641),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1685),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1660),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1701),
.A2(n_1704),
.B1(n_1580),
.B2(n_1587),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1697),
.B(n_1641),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1558),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1536),
.A2(n_1662),
.B(n_1601),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1712),
.B(n_1583),
.Y(n_1776)
);

AO31x2_ASAP7_75t_L g1777 ( 
.A1(n_1603),
.A2(n_1606),
.A3(n_1562),
.B(n_1568),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1559),
.Y(n_1778)
);

AO21x2_ASAP7_75t_L g1779 ( 
.A1(n_1563),
.A2(n_1579),
.B(n_1611),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1613),
.A2(n_1633),
.B(n_1540),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1582),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1541),
.B(n_1674),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1565),
.B(n_1711),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1574),
.B(n_1713),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1598),
.B(n_1584),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1677),
.B(n_1679),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1660),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1680),
.B(n_1682),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1684),
.B(n_1686),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1698),
.B(n_1703),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1598),
.B(n_1632),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1678),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_L g1793 ( 
.A(n_1662),
.B(n_1587),
.C(n_1669),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1548),
.B(n_1561),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1708),
.B(n_1710),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1571),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1554),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1628),
.Y(n_1798)
);

BUFx12f_ASAP7_75t_L g1799 ( 
.A(n_1585),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1591),
.B(n_1615),
.Y(n_1800)
);

OAI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1540),
.A2(n_1550),
.B(n_1705),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1594),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1702),
.B(n_1543),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1545),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1636),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1629),
.B(n_1631),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1592),
.A2(n_1621),
.B(n_1602),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1652),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1590),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1653),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1656),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1658),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1578),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1554),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1649),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1658),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1621),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1664),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1621),
.Y(n_1819)
);

AO21x2_ASAP7_75t_L g1820 ( 
.A1(n_1637),
.A2(n_1647),
.B(n_1644),
.Y(n_1820)
);

OR2x6_ASAP7_75t_L g1821 ( 
.A(n_1548),
.B(n_1561),
.Y(n_1821)
);

AO21x2_ASAP7_75t_L g1822 ( 
.A1(n_1638),
.A2(n_1646),
.B(n_1639),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1659),
.A2(n_1596),
.B(n_1634),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1560),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1643),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1593),
.Y(n_1826)
);

AO21x2_ASAP7_75t_L g1827 ( 
.A1(n_1604),
.A2(n_1605),
.B(n_1626),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1560),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1648),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1709),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1670),
.B(n_1709),
.Y(n_1831)
);

AOI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1635),
.A2(n_1627),
.B(n_1645),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1694),
.B(n_1618),
.Y(n_1833)
);

OA21x2_ASAP7_75t_L g1834 ( 
.A1(n_1608),
.A2(n_1597),
.B(n_1665),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1673),
.B(n_1619),
.Y(n_1835)
);

NAND2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1618),
.B(n_1688),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1692),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1692),
.Y(n_1838)
);

INVxp33_ASAP7_75t_L g1839 ( 
.A(n_1547),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1595),
.B(n_1688),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1714),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1692),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1714),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1595),
.B(n_1665),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1602),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1597),
.B(n_1693),
.Y(n_1846)
);

AO21x2_ASAP7_75t_L g1847 ( 
.A1(n_1654),
.A2(n_1714),
.B(n_1619),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1827),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1736),
.B(n_1683),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1779),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1722),
.B(n_1746),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1736),
.B(n_1683),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1760),
.B(n_1763),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1774),
.Y(n_1854)
);

AO21x2_ASAP7_75t_L g1855 ( 
.A1(n_1739),
.A2(n_1687),
.B(n_1693),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1760),
.B(n_1622),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1774),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1778),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1761),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1728),
.A2(n_1551),
.B1(n_1695),
.B2(n_1700),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1720),
.A2(n_1687),
.B(n_1695),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1778),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1770),
.B(n_1555),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1722),
.B(n_1699),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1834),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1770),
.B(n_1578),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1756),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1834),
.Y(n_1868)
);

OAI31xp33_ASAP7_75t_SL g1869 ( 
.A1(n_1718),
.A2(n_1551),
.A3(n_1695),
.B(n_1691),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1813),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1746),
.B(n_1699),
.Y(n_1871)
);

AOI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1755),
.A2(n_1600),
.B1(n_1700),
.B2(n_1622),
.C(n_1551),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1767),
.B(n_1578),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1827),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1834),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1727),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1735),
.Y(n_1877)
);

AND2x4_ASAP7_75t_SL g1878 ( 
.A(n_1826),
.B(n_1661),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1719),
.B(n_1691),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1767),
.B(n_1630),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1758),
.B(n_1630),
.Y(n_1881)
);

AND2x6_ASAP7_75t_L g1882 ( 
.A(n_1763),
.B(n_1623),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1758),
.B(n_1575),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1741),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1839),
.B(n_1552),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1764),
.A2(n_1600),
.B(n_1585),
.Y(n_1886)
);

AOI222xp33_ASAP7_75t_L g1887 ( 
.A1(n_1775),
.A2(n_1772),
.B1(n_1733),
.B2(n_1793),
.C1(n_1734),
.C2(n_1783),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1800),
.B(n_1750),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1799),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1749),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1768),
.B(n_1752),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1784),
.B(n_1768),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1834),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1776),
.B(n_1723),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1721),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1752),
.B(n_1749),
.Y(n_1896)
);

NAND2xp33_ASAP7_75t_R g1897 ( 
.A(n_1802),
.B(n_1823),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1765),
.B(n_1781),
.Y(n_1898)
);

INVxp67_ASAP7_75t_SL g1899 ( 
.A(n_1784),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1752),
.B(n_1771),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1776),
.B(n_1723),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1721),
.Y(n_1902)
);

OAI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1791),
.A2(n_1785),
.B1(n_1743),
.B2(n_1762),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1777),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1798),
.B(n_1796),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1771),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1764),
.B(n_1729),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1777),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1777),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1777),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1787),
.B(n_1730),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1802),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1777),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1809),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1715),
.B(n_1717),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1724),
.B(n_1747),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1797),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1823),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1822),
.Y(n_1919)
);

AND2x4_ASAP7_75t_SL g1920 ( 
.A(n_1815),
.B(n_1769),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1806),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1742),
.B(n_1725),
.Y(n_1922)
);

AOI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1764),
.A2(n_1737),
.B1(n_1792),
.B2(n_1791),
.C(n_1785),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1777),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1831),
.A2(n_1835),
.B1(n_1841),
.B2(n_1843),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1888),
.B(n_1914),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1899),
.B(n_1740),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1876),
.B(n_1740),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1894),
.B(n_1759),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1877),
.B(n_1737),
.Y(n_1930)
);

NOR3xp33_ASAP7_75t_L g1931 ( 
.A(n_1872),
.B(n_1838),
.C(n_1837),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1894),
.B(n_1759),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1901),
.B(n_1759),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1923),
.B(n_1769),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1869),
.A2(n_1835),
.B1(n_1744),
.B2(n_1716),
.C(n_1831),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1901),
.B(n_1759),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1884),
.B(n_1823),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_L g1938 ( 
.A(n_1887),
.B(n_1762),
.C(n_1744),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1860),
.A2(n_1769),
.B(n_1773),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1886),
.B(n_1762),
.C(n_1819),
.Y(n_1940)
);

OAI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1886),
.A2(n_1716),
.B1(n_1762),
.B2(n_1745),
.C(n_1806),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1898),
.B(n_1804),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1859),
.A2(n_1754),
.B1(n_1745),
.B2(n_1799),
.Y(n_1943)
);

OAI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1871),
.A2(n_1838),
.B1(n_1837),
.B2(n_1842),
.C(n_1814),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1871),
.A2(n_1769),
.B1(n_1773),
.B2(n_1766),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_R g1946 ( 
.A(n_1889),
.B(n_1754),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1864),
.A2(n_1847),
.B(n_1821),
.Y(n_1947)
);

AOI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1903),
.A2(n_1786),
.B1(n_1795),
.B2(n_1782),
.C(n_1790),
.Y(n_1948)
);

NAND3xp33_ASAP7_75t_L g1949 ( 
.A(n_1864),
.B(n_1819),
.C(n_1829),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1907),
.B(n_1829),
.C(n_1842),
.Y(n_1950)
);

OAI221xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1851),
.A2(n_1795),
.B1(n_1790),
.B2(n_1789),
.C(n_1788),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1921),
.B(n_1804),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1896),
.B(n_1780),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1905),
.B(n_1805),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1912),
.B(n_1805),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1892),
.B(n_1726),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1897),
.B(n_1842),
.C(n_1818),
.Y(n_1957)
);

NOR3xp33_ASAP7_75t_SL g1958 ( 
.A(n_1889),
.B(n_1840),
.C(n_1818),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1922),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1892),
.B(n_1895),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1902),
.B(n_1731),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1854),
.B(n_1808),
.Y(n_1962)
);

OAI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1879),
.A2(n_1794),
.B1(n_1821),
.B2(n_1828),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1857),
.B(n_1808),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1878),
.A2(n_1885),
.B1(n_1856),
.B2(n_1863),
.Y(n_1965)
);

NOR3xp33_ASAP7_75t_SL g1966 ( 
.A(n_1925),
.B(n_1816),
.C(n_1812),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1915),
.B(n_1748),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1858),
.B(n_1862),
.Y(n_1968)
);

NAND4xp25_ASAP7_75t_L g1969 ( 
.A(n_1881),
.B(n_1782),
.C(n_1786),
.D(n_1788),
.Y(n_1969)
);

OAI21xp33_ASAP7_75t_SL g1970 ( 
.A1(n_1868),
.A2(n_1766),
.B(n_1807),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1915),
.B(n_1748),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1883),
.A2(n_1773),
.B1(n_1847),
.B2(n_1820),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1870),
.B(n_1773),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1851),
.B(n_1748),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1853),
.B(n_1748),
.Y(n_1975)
);

OAI21xp33_ASAP7_75t_SL g1976 ( 
.A1(n_1863),
.A2(n_1807),
.B(n_1801),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1883),
.A2(n_1856),
.B1(n_1881),
.B2(n_1880),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1853),
.B(n_1753),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1853),
.B(n_1753),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1856),
.A2(n_1847),
.B1(n_1820),
.B2(n_1828),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1867),
.B(n_1866),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1866),
.B(n_1822),
.Y(n_1982)
);

NAND3xp33_ASAP7_75t_L g1983 ( 
.A(n_1848),
.B(n_1816),
.C(n_1812),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1873),
.B(n_1822),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1873),
.B(n_1803),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1878),
.A2(n_1833),
.B(n_1836),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1911),
.B(n_1753),
.Y(n_1987)
);

NAND3xp33_ASAP7_75t_L g1988 ( 
.A(n_1874),
.B(n_1817),
.C(n_1845),
.Y(n_1988)
);

NOR3xp33_ASAP7_75t_L g1989 ( 
.A(n_1861),
.B(n_1845),
.C(n_1738),
.Y(n_1989)
);

NAND4xp25_ASAP7_75t_L g1990 ( 
.A(n_1919),
.B(n_1789),
.C(n_1811),
.D(n_1810),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1880),
.A2(n_1830),
.B1(n_1824),
.B2(n_1828),
.Y(n_1991)
);

OAI21xp5_ASAP7_75t_SL g1992 ( 
.A1(n_1896),
.A2(n_1833),
.B(n_1836),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1911),
.B(n_1753),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1849),
.B(n_1811),
.Y(n_1994)
);

OA21x2_ASAP7_75t_L g1995 ( 
.A1(n_1850),
.A2(n_1757),
.B(n_1751),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1852),
.B(n_1732),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_SL g1997 ( 
.A1(n_1917),
.A2(n_1794),
.B(n_1821),
.Y(n_1997)
);

NAND3xp33_ASAP7_75t_L g1998 ( 
.A(n_1918),
.B(n_1817),
.C(n_1825),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1937),
.B(n_1960),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1956),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1974),
.Y(n_2001)
);

NOR2x1_ASAP7_75t_L g2002 ( 
.A(n_1957),
.B(n_1865),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1929),
.B(n_1865),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1929),
.B(n_1875),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1959),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1995),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1959),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1932),
.B(n_1919),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1933),
.B(n_1893),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1995),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1968),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1936),
.B(n_1904),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1946),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1975),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1936),
.B(n_1908),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1976),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1953),
.B(n_1890),
.Y(n_2017)
);

AOI211x1_ASAP7_75t_L g2018 ( 
.A1(n_1938),
.A2(n_1832),
.B(n_1846),
.C(n_1844),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1984),
.B(n_1916),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1962),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1927),
.B(n_1909),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1930),
.B(n_1910),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1964),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1961),
.Y(n_2024)
);

NAND2x1p5_ASAP7_75t_L g2025 ( 
.A(n_1934),
.B(n_1861),
.Y(n_2025)
);

AND2x2_ASAP7_75t_SL g2026 ( 
.A(n_1972),
.B(n_1896),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1989),
.B(n_1906),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1982),
.B(n_1913),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1998),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1981),
.B(n_1916),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1978),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1942),
.B(n_1924),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1952),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_1950),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1987),
.B(n_1906),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1979),
.B(n_1900),
.Y(n_2036)
);

INVxp67_ASAP7_75t_SL g2037 ( 
.A(n_1983),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1967),
.B(n_1900),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1967),
.B(n_1900),
.Y(n_2039)
);

AND2x2_ASAP7_75t_SL g2040 ( 
.A(n_1980),
.B(n_1920),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_1940),
.B(n_1855),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_1994),
.B(n_1955),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1987),
.B(n_1993),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_2014),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2043),
.B(n_1993),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2043),
.B(n_1971),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2033),
.B(n_2034),
.Y(n_2047)
);

INVxp67_ASAP7_75t_L g2048 ( 
.A(n_2029),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2005),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2009),
.B(n_1926),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2005),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2033),
.B(n_1985),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2034),
.B(n_1954),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2007),
.Y(n_2054)
);

INVxp67_ASAP7_75t_L g2055 ( 
.A(n_2029),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2043),
.B(n_1947),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2043),
.B(n_1947),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2007),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2035),
.B(n_1992),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2011),
.B(n_1934),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2035),
.B(n_1997),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2000),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2035),
.B(n_1997),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2035),
.B(n_1973),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2009),
.B(n_1990),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_2006),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2008),
.B(n_1928),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2031),
.B(n_2017),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2008),
.B(n_1996),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2011),
.B(n_1948),
.Y(n_2070)
);

NOR2x1_ASAP7_75t_L g2071 ( 
.A(n_2002),
.B(n_1988),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_2013),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2006),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1999),
.B(n_1949),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2031),
.B(n_1973),
.Y(n_2075)
);

INVx2_ASAP7_75t_SL g2076 ( 
.A(n_2014),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2006),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2021),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2010),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2031),
.B(n_1891),
.Y(n_2080)
);

NAND4xp75_ASAP7_75t_L g2081 ( 
.A(n_2002),
.B(n_1958),
.C(n_1970),
.D(n_1966),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2010),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_2021),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_2014),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_2025),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2010),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_2024),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_2016),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2001),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2001),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2048),
.B(n_2037),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2088),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2081),
.A2(n_2040),
.B1(n_2026),
.B2(n_1963),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2055),
.B(n_2047),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2049),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2049),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2051),
.Y(n_2097)
);

OR2x6_ASAP7_75t_L g2098 ( 
.A(n_2081),
.B(n_1986),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2065),
.B(n_1999),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2087),
.B(n_2037),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2065),
.B(n_2042),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2074),
.B(n_2024),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2045),
.B(n_2036),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2059),
.B(n_2017),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_2059),
.B(n_2017),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2051),
.Y(n_2106)
);

NOR2xp67_ASAP7_75t_L g2107 ( 
.A(n_2056),
.B(n_2027),
.Y(n_2107)
);

OAI211xp5_ASAP7_75t_SL g2108 ( 
.A1(n_2071),
.A2(n_2041),
.B(n_1977),
.C(n_1941),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2050),
.B(n_2042),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2070),
.B(n_2078),
.Y(n_2110)
);

OR2x6_ASAP7_75t_L g2111 ( 
.A(n_2071),
.B(n_2025),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_2088),
.B(n_2041),
.Y(n_2112)
);

NAND2x1_ASAP7_75t_L g2113 ( 
.A(n_2056),
.B(n_2016),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2050),
.B(n_2019),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2054),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2054),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2045),
.B(n_2036),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2083),
.B(n_2020),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2046),
.B(n_2038),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2058),
.Y(n_2120)
);

NAND2x1_ASAP7_75t_L g2121 ( 
.A(n_2057),
.B(n_2075),
.Y(n_2121)
);

AOI21x1_ASAP7_75t_SL g2122 ( 
.A1(n_2060),
.A2(n_2027),
.B(n_2022),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2058),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2089),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2067),
.B(n_2030),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2053),
.B(n_2020),
.Y(n_2126)
);

NOR2x1_ASAP7_75t_L g2127 ( 
.A(n_2072),
.B(n_1943),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_2044),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2046),
.B(n_2064),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2089),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_2052),
.B(n_1965),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2068),
.Y(n_2132)
);

OAI21xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2057),
.A2(n_2026),
.B(n_2040),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2064),
.B(n_2038),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2044),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2090),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2068),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2061),
.B(n_2039),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2067),
.B(n_2023),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2080),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2090),
.B(n_2023),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2069),
.B(n_2030),
.Y(n_2142)
);

INVx1_ASAP7_75t_SL g2143 ( 
.A(n_2076),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2080),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2092),
.Y(n_2145)
);

INVx1_ASAP7_75t_SL g2146 ( 
.A(n_2128),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2095),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_2111),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2096),
.Y(n_2149)
);

INVx2_ASAP7_75t_SL g2150 ( 
.A(n_2111),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2097),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2098),
.A2(n_2026),
.B1(n_2040),
.B2(n_2063),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2111),
.B(n_2061),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2106),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2112),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2115),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2112),
.Y(n_2157)
);

BUFx3_ASAP7_75t_L g2158 ( 
.A(n_2098),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2093),
.A2(n_2018),
.B1(n_2025),
.B2(n_1951),
.Y(n_2159)
);

AOI222xp33_ASAP7_75t_L g2160 ( 
.A1(n_2108),
.A2(n_1935),
.B1(n_1970),
.B2(n_1939),
.C1(n_1945),
.C2(n_2085),
.Y(n_2160)
);

INVx5_ASAP7_75t_L g2161 ( 
.A(n_2098),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2116),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2120),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2123),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2124),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2129),
.B(n_2063),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2107),
.B(n_2085),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2110),
.B(n_2062),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2130),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2104),
.B(n_2075),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2128),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2135),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_2143),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2127),
.B(n_2069),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_2143),
.Y(n_2175)
);

OAI21xp33_ASAP7_75t_L g2176 ( 
.A1(n_2108),
.A2(n_2091),
.B(n_2110),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_2136),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2135),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2141),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2141),
.Y(n_2180)
);

INVx1_ASAP7_75t_SL g2181 ( 
.A(n_2091),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2101),
.B(n_2062),
.Y(n_2182)
);

INVxp33_ASAP7_75t_SL g2183 ( 
.A(n_2131),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2104),
.B(n_2105),
.Y(n_2184)
);

NOR2x1_ASAP7_75t_L g2185 ( 
.A(n_2113),
.B(n_2073),
.Y(n_2185)
);

INVx1_ASAP7_75t_SL g2186 ( 
.A(n_2145),
.Y(n_2186)
);

AOI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2176),
.A2(n_2100),
.B1(n_2094),
.B2(n_2133),
.C(n_2102),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2184),
.B(n_2138),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2171),
.Y(n_2189)
);

NOR2x1_ASAP7_75t_L g2190 ( 
.A(n_2158),
.B(n_2094),
.Y(n_2190)
);

NOR3xp33_ASAP7_75t_L g2191 ( 
.A(n_2176),
.B(n_2100),
.C(n_2121),
.Y(n_2191)
);

OAI21xp33_ASAP7_75t_L g2192 ( 
.A1(n_2158),
.A2(n_2099),
.B(n_2102),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2184),
.B(n_2170),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2171),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2183),
.B(n_2126),
.Y(n_2195)
);

OAI21xp5_ASAP7_75t_SL g2196 ( 
.A1(n_2160),
.A2(n_2025),
.B(n_2105),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2145),
.B(n_2126),
.Y(n_2197)
);

NOR2x1_ASAP7_75t_L g2198 ( 
.A(n_2158),
.B(n_2118),
.Y(n_2198)
);

AO22x1_ASAP7_75t_L g2199 ( 
.A1(n_2161),
.A2(n_2084),
.B1(n_2076),
.B2(n_2132),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2173),
.Y(n_2200)
);

NAND3xp33_ASAP7_75t_L g2201 ( 
.A(n_2161),
.B(n_2018),
.C(n_1931),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2174),
.B(n_2137),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2173),
.Y(n_2203)
);

O2A1O1Ixp33_ASAP7_75t_L g2204 ( 
.A1(n_2159),
.A2(n_2118),
.B(n_2139),
.C(n_2084),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2175),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2152),
.A2(n_2109),
.B1(n_2125),
.B2(n_2142),
.Y(n_2206)
);

OAI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_2161),
.A2(n_2139),
.B(n_2027),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2185),
.Y(n_2208)
);

OAI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_2161),
.A2(n_1969),
.B1(n_1944),
.B2(n_2114),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2184),
.B(n_2134),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2159),
.A2(n_2140),
.B1(n_2144),
.B2(n_2027),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2185),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2161),
.A2(n_1882),
.B1(n_1820),
.B2(n_2117),
.Y(n_2213)
);

OAI21xp33_ASAP7_75t_L g2214 ( 
.A1(n_2160),
.A2(n_2028),
.B(n_2022),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2175),
.Y(n_2215)
);

OAI221xp5_ASAP7_75t_L g2216 ( 
.A1(n_2161),
.A2(n_2028),
.B1(n_2122),
.B2(n_2032),
.C(n_1991),
.Y(n_2216)
);

AOI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_2191),
.A2(n_2161),
.B1(n_2166),
.B2(n_2170),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_2191),
.A2(n_2166),
.B1(n_2170),
.B2(n_2181),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2186),
.B(n_2146),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2189),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2194),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2200),
.B(n_2146),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2203),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2193),
.B(n_2166),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2190),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2205),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2215),
.B(n_2181),
.Y(n_2227)
);

INVx1_ASAP7_75t_SL g2228 ( 
.A(n_2198),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2208),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2195),
.B(n_2172),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2197),
.B(n_2168),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_2202),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2195),
.B(n_2172),
.Y(n_2233)
);

NAND3xp33_ASAP7_75t_L g2234 ( 
.A(n_2204),
.B(n_2177),
.C(n_2169),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_2209),
.B(n_2153),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2188),
.B(n_2172),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2192),
.B(n_2178),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2196),
.A2(n_2148),
.B1(n_2150),
.B2(n_2153),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2208),
.Y(n_2239)
);

NOR3xp33_ASAP7_75t_L g2240 ( 
.A(n_2219),
.B(n_2206),
.C(n_2187),
.Y(n_2240)
);

OAI221xp5_ASAP7_75t_L g2241 ( 
.A1(n_2217),
.A2(n_2211),
.B1(n_2201),
.B2(n_2214),
.C(n_2207),
.Y(n_2241)
);

NAND4xp25_ASAP7_75t_SL g2242 ( 
.A(n_2228),
.B(n_2216),
.C(n_2153),
.D(n_2213),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_2235),
.A2(n_2209),
.B(n_2199),
.Y(n_2243)
);

AOI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_2225),
.A2(n_2180),
.B1(n_2179),
.B2(n_2212),
.C(n_2150),
.Y(n_2244)
);

NAND2xp33_ASAP7_75t_SL g2245 ( 
.A(n_2224),
.B(n_2148),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2222),
.Y(n_2246)
);

OAI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_2234),
.A2(n_2212),
.B1(n_2148),
.B2(n_2150),
.Y(n_2247)
);

NAND3xp33_ASAP7_75t_L g2248 ( 
.A(n_2234),
.B(n_2213),
.C(n_2178),
.Y(n_2248)
);

AOI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_2218),
.A2(n_2238),
.B1(n_2232),
.B2(n_2237),
.C(n_2227),
.Y(n_2249)
);

AOI211xp5_ASAP7_75t_L g2250 ( 
.A1(n_2230),
.A2(n_2210),
.B(n_2155),
.C(n_2157),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2224),
.B(n_2178),
.Y(n_2251)
);

AOI211xp5_ASAP7_75t_SL g2252 ( 
.A1(n_2233),
.A2(n_2167),
.B(n_2177),
.C(n_2155),
.Y(n_2252)
);

AOI211xp5_ASAP7_75t_L g2253 ( 
.A1(n_2220),
.A2(n_2157),
.B(n_2155),
.C(n_2167),
.Y(n_2253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2254 ( 
.A1(n_2220),
.A2(n_2180),
.B(n_2179),
.C(n_2165),
.D(n_2169),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2243),
.A2(n_2231),
.B1(n_2236),
.B2(n_2223),
.Y(n_2255)
);

NAND3xp33_ASAP7_75t_L g2256 ( 
.A(n_2254),
.B(n_2223),
.C(n_2221),
.Y(n_2256)
);

NAND4xp75_ASAP7_75t_L g2257 ( 
.A(n_2249),
.B(n_2221),
.C(n_2226),
.D(n_2239),
.Y(n_2257)
);

OAI211xp5_ASAP7_75t_L g2258 ( 
.A1(n_2252),
.A2(n_2226),
.B(n_2231),
.C(n_2239),
.Y(n_2258)
);

NOR3x1_ASAP7_75t_L g2259 ( 
.A(n_2241),
.B(n_2165),
.C(n_2168),
.Y(n_2259)
);

NOR4xp75_ASAP7_75t_L g2260 ( 
.A(n_2251),
.B(n_2236),
.C(n_2167),
.D(n_2229),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2246),
.Y(n_2261)
);

NOR2x1_ASAP7_75t_L g2262 ( 
.A(n_2247),
.B(n_2229),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2240),
.A2(n_2157),
.B1(n_2156),
.B2(n_2162),
.Y(n_2263)
);

NAND4xp25_ASAP7_75t_L g2264 ( 
.A(n_2244),
.B(n_2149),
.C(n_2151),
.D(n_2154),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2250),
.B(n_2147),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2253),
.B(n_2103),
.Y(n_2266)
);

NOR3xp33_ASAP7_75t_L g2267 ( 
.A(n_2245),
.B(n_2149),
.C(n_2147),
.Y(n_2267)
);

OAI22xp33_ASAP7_75t_SL g2268 ( 
.A1(n_2262),
.A2(n_2151),
.B1(n_2156),
.B2(n_2162),
.Y(n_2268)
);

NOR2xp67_ASAP7_75t_L g2269 ( 
.A(n_2258),
.B(n_2248),
.Y(n_2269)
);

NOR2x1_ASAP7_75t_L g2270 ( 
.A(n_2257),
.B(n_2242),
.Y(n_2270)
);

NOR3xp33_ASAP7_75t_L g2271 ( 
.A(n_2255),
.B(n_2154),
.C(n_2163),
.Y(n_2271)
);

NAND4xp25_ASAP7_75t_L g2272 ( 
.A(n_2259),
.B(n_2164),
.C(n_2163),
.D(n_2182),
.Y(n_2272)
);

OAI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2256),
.A2(n_2164),
.B(n_2163),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2263),
.B(n_2164),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2269),
.A2(n_2266),
.B1(n_2267),
.B2(n_2265),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2274),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2268),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2270),
.A2(n_2261),
.B1(n_2264),
.B2(n_2182),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_2272),
.Y(n_2279)
);

NOR2x1_ASAP7_75t_L g2280 ( 
.A(n_2273),
.B(n_2260),
.Y(n_2280)
);

AOI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2271),
.A2(n_2073),
.B1(n_2077),
.B2(n_2079),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2272),
.B(n_2119),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2280),
.A2(n_2077),
.B(n_2073),
.Y(n_2283)
);

NOR4xp75_ASAP7_75t_SL g2284 ( 
.A(n_2275),
.B(n_2015),
.C(n_2012),
.D(n_2032),
.Y(n_2284)
);

NAND3xp33_ASAP7_75t_L g2285 ( 
.A(n_2278),
.B(n_2079),
.C(n_2077),
.Y(n_2285)
);

NAND3x1_ASAP7_75t_SL g2286 ( 
.A(n_2276),
.B(n_2004),
.C(n_2003),
.Y(n_2286)
);

INVxp67_ASAP7_75t_L g2287 ( 
.A(n_2277),
.Y(n_2287)
);

NOR2x1_ASAP7_75t_L g2288 ( 
.A(n_2279),
.B(n_2066),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2288),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2287),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2286),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2291),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2292),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2293),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2293),
.Y(n_2295)
);

AOI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2294),
.A2(n_2290),
.B(n_2295),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2295),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2297),
.B(n_2282),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2296),
.A2(n_2289),
.B(n_2283),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2299),
.B(n_2285),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_SL g2301 ( 
.A1(n_2300),
.A2(n_2298),
.B1(n_2284),
.B2(n_2066),
.Y(n_2301)
);

AOI221xp5_ASAP7_75t_L g2302 ( 
.A1(n_2301),
.A2(n_2281),
.B1(n_2079),
.B2(n_2086),
.C(n_2082),
.Y(n_2302)
);

AOI211xp5_ASAP7_75t_L g2303 ( 
.A1(n_2302),
.A2(n_2086),
.B(n_2082),
.C(n_2066),
.Y(n_2303)
);


endmodule