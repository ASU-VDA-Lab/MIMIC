module real_jpeg_26453_n_16 (n_5, n_4, n_8, n_0, n_12, n_360, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_360;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_1),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_1),
.A2(n_43),
.B1(n_80),
.B2(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_26),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_2),
.A2(n_70),
.B1(n_80),
.B2(n_81),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_3),
.A2(n_80),
.B1(n_81),
.B2(n_110),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_110),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_24),
.B1(n_71),
.B2(n_110),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_80),
.B1(n_81),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_127),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_127),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_4),
.A2(n_26),
.B1(n_39),
.B2(n_127),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_6),
.A2(n_80),
.B1(n_81),
.B2(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_119),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_6),
.A2(n_23),
.B1(n_119),
.B2(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_9),
.A2(n_25),
.B1(n_80),
.B2(n_81),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_9),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_68),
.B1(n_80),
.B2(n_81),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_68),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_11),
.A2(n_76),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_122),
.B1(n_146),
.B2(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_11),
.A2(n_34),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_11),
.B(n_45),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_15),
.Y(n_131)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_15),
.Y(n_139)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_93),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_46),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_20),
.B(n_46),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_21),
.A2(n_30),
.B(n_66),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_22),
.B(n_45),
.Y(n_87)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_23),
.Y(n_245)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_24),
.A2(n_31),
.A3(n_35),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_28),
.A2(n_45),
.B1(n_65),
.B2(n_69),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_28),
.A2(n_69),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_28),
.A2(n_45),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_28),
.A2(n_45),
.B1(n_232),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_29),
.A2(n_30),
.B1(n_244),
.B2(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_29),
.A2(n_40),
.B(n_262),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_29),
.A2(n_87),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_32),
.B(n_34),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_35),
.B1(n_54),
.B2(n_58),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_34),
.A2(n_54),
.A3(n_56),
.B1(n_162),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_35),
.B(n_106),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_39),
.A2(n_106),
.B(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_41),
.Y(n_311)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_42),
.B(n_106),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_85),
.C(n_88),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_47),
.A2(n_48),
.B1(n_353),
.B2(n_355),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_64),
.C(n_72),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_49),
.A2(n_50),
.B1(n_72),
.B2(n_73),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_52),
.A2(n_61),
.B(n_226),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_53),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_53),
.A2(n_60),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_56),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_55),
.B(n_58),
.Y(n_171)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_56),
.A2(n_78),
.B(n_106),
.C(n_112),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_59),
.A2(n_163),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_61),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_61),
.A2(n_90),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_61),
.A2(n_90),
.B1(n_189),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_61),
.A2(n_90),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_61),
.A2(n_302),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_63),
.B(n_90),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_64),
.B(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_72),
.A2(n_73),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_73),
.B(n_330),
.C(n_332),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_83),
.B(n_84),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_83),
.B1(n_109),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_74),
.A2(n_83),
.B1(n_118),
.B2(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_74),
.A2(n_84),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_74),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_79),
.B(n_106),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_79),
.B(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_79),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_79),
.A2(n_107),
.B1(n_251),
.B2(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_80),
.B(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_83),
.B(n_84),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_85),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_351),
.B(n_357),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_326),
.A3(n_344),
.B1(n_349),
.B2(n_350),
.C(n_360),
.Y(n_94)
);

AOI311xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_279),
.A3(n_316),
.B(n_320),
.C(n_321),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_234),
.C(n_274),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_206),
.B(n_233),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_182),
.B(n_205),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_155),
.B(n_181),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_132),
.B(n_154),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_102),
.B(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_104),
.B1(n_111),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_149),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_107),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_107),
.A2(n_269),
.B(n_294),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B(n_128),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_131),
.B1(n_136),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_122),
.A2(n_174),
.B(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_122),
.A2(n_149),
.B(n_173),
.Y(n_291)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_123),
.B(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_123),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_128),
.B(n_196),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_142),
.B(n_153),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_140),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_139),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_147),
.B(n_152),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_157),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_169),
.B1(n_179),
.B2(n_180),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_168),
.C(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_184),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_197),
.B2(n_198),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_200),
.C(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_192),
.C(n_193),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_202),
.B(n_252),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_208),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_223),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_222),
.C(n_223),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_214),
.B1(n_218),
.B2(n_219),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_218),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_214),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_227),
.C(n_230),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_235),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_254),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_236),
.B(n_254),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_246),
.C(n_247),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_238),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_246),
.B(n_247),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_250),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_266),
.B2(n_270),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_270),
.C(n_273),
.Y(n_318)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_265),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_268),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_280),
.A2(n_317),
.B(n_322),
.C(n_325),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_297),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_297),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.C(n_296),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_282),
.B(n_290),
.CI(n_296),
.CON(n_319),
.SN(n_319)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_289),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_286),
.C(n_287),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_295),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_291),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_295),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_306),
.B(n_310),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_315),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_305),
.B1(n_313),
.B2(n_314),
.Y(n_298)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_303),
.B(n_304),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_303),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_304),
.A2(n_328),
.B1(n_336),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_313),
.C(n_315),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_312),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_319),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_338),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_327),
.B(n_338),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_336),
.C(n_337),
.Y(n_327)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_335),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_330),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_342),
.C(n_343),
.Y(n_356)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_345),
.B(n_346),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_356),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_352),
.B(n_356),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_353),
.Y(n_355)
);


endmodule