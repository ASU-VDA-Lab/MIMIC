module fake_jpeg_10961_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_44),
.C(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_33),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_22),
.B1(n_41),
.B2(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_56),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_25),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_61),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_64),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_18),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_66),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_42),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_35),
.B1(n_33),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_30),
.B1(n_27),
.B2(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_44),
.B1(n_30),
.B2(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_81),
.B1(n_88),
.B2(n_26),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_47),
.B1(n_37),
.B2(n_40),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_89),
.B1(n_100),
.B2(n_26),
.Y(n_126)
);

AO22x2_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_47),
.B1(n_37),
.B2(n_40),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_63),
.B1(n_51),
.B2(n_60),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_32),
.B(n_24),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_84),
.C(n_85),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_36),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_36),
.C(n_19),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_40),
.B1(n_37),
.B2(n_41),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_31),
.B1(n_32),
.B2(n_19),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_101),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_29),
.B(n_24),
.C(n_23),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_51),
.B(n_34),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_116),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_54),
.B1(n_45),
.B2(n_57),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_41),
.B1(n_70),
.B2(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_114),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_70),
.B1(n_55),
.B2(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_70),
.B1(n_48),
.B2(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_118),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_54),
.B1(n_45),
.B2(n_46),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_12),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_0),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_0),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_122),
.C(n_107),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_46),
.B1(n_51),
.B2(n_60),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_87),
.B1(n_76),
.B2(n_78),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_1),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_60),
.B(n_46),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_77),
.B(n_90),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_129),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_128),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_99),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_140),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx2_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_143),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_155),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_95),
.B(n_82),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_81),
.B1(n_87),
.B2(n_80),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_154),
.Y(n_184)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_151),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_114),
.Y(n_162)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_78),
.B(n_76),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_110),
.B(n_104),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_142),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_165),
.B(n_173),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_119),
.C(n_123),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_169),
.C(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_122),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_136),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_13),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_130),
.B1(n_128),
.B2(n_117),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_161),
.B1(n_147),
.B2(n_154),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_121),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_117),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_189),
.C(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_117),
.B(n_127),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_141),
.B(n_188),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_155),
.B(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_117),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_11),
.C(n_16),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_127),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_135),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_10),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_193),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_202),
.B1(n_212),
.B2(n_183),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_149),
.B1(n_143),
.B2(n_131),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_163),
.B(n_171),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_205),
.B(n_206),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_184),
.B1(n_131),
.B2(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_155),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_211),
.C(n_163),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_149),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_148),
.B1(n_134),
.B2(n_135),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_152),
.B1(n_158),
.B2(n_144),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_157),
.B(n_11),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_182),
.B(n_164),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_222),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_153),
.B1(n_34),
.B2(n_28),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_220),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_248),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_179),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_204),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_238),
.B(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_198),
.C(n_196),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_197),
.C(n_26),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_164),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_202),
.A2(n_172),
.B1(n_178),
.B2(n_185),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_200),
.B1(n_197),
.B2(n_213),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_201),
.A2(n_168),
.B(n_153),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_168),
.B(n_189),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_8),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_215),
.B1(n_212),
.B2(n_209),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_251),
.A2(n_260),
.B1(n_245),
.B2(n_235),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_210),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_253),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_224),
.B(n_205),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_257),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_218),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_253),
.C(n_252),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_34),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_265),
.B(n_246),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_26),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_26),
.C(n_9),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_249),
.C(n_247),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_274),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_233),
.B1(n_225),
.B2(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_289),
.B1(n_248),
.B2(n_226),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_267),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_225),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_288),
.C(n_274),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_235),
.C(n_230),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_255),
.C(n_259),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_243),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_240),
.B1(n_250),
.B2(n_227),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_262),
.B(n_263),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_304),
.B(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

AO22x1_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_256),
.B1(n_262),
.B2(n_248),
.Y(n_295)
);

OAI211xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_285),
.B(n_279),
.C(n_277),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_268),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_239),
.C(n_9),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_299),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_239),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_7),
.C(n_15),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_6),
.C(n_15),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_10),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_278),
.B(n_7),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_279),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_275),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_311),
.A2(n_313),
.B(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_316),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_300),
.B(n_12),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_15),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_3),
.C(n_5),
.Y(n_316)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_318),
.B(n_320),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_295),
.B(n_297),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_323),
.B(n_13),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_301),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_5),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_13),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_16),
.C(n_1),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_312),
.B(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_321),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_307),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_331),
.C(n_327),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_330),
.C(n_322),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_1),
.B1(n_2),
.B2(n_327),
.Y(n_339)
);


endmodule