module fake_jpeg_17086_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_14),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_9),
.A2(n_4),
.B1(n_5),
.B2(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_5),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_6),
.B(n_10),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_10),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_20),
.B(n_21),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_6),
.B(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_17),
.B1(n_12),
.B2(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

XNOR2x1_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_7),
.B1(n_8),
.B2(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_23),
.B1(n_16),
.B2(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_3),
.B1(n_32),
.B2(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_20),
.B1(n_23),
.B2(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_16),
.C(n_0),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_31),
.C(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_35),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_33),
.A3(n_32),
.B1(n_41),
.B2(n_35),
.C1(n_37),
.C2(n_36),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_32),
.B(n_35),
.Y(n_44)
);


endmodule