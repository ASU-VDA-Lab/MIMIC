module fake_netlist_6_73_n_1697 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1697);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1697;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_165),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_56),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_57),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_133),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_0),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_48),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_78),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_8),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_15),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_81),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_64),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_15),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_97),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_38),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_134),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_51),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_31),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_17),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_28),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_114),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_59),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_9),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_48),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_129),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_49),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_40),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_63),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_80),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_118),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_18),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_161),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_74),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_38),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_96),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_126),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_93),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_154),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_163),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_123),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_115),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_39),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_146),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_66),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_89),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_157),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_29),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_5),
.Y(n_253)
);

CKINVDCx11_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_55),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_54),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_71),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_62),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_67),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_68),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_21),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_125),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_33),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_47),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_60),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_127),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_45),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_12),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_151),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_47),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_105),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_95),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_100),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_117),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_49),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_140),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_22),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_53),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_50),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_41),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_98),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_73),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_26),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_12),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_25),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_102),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_16),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_85),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_16),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_39),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_86),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_122),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_94),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_19),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_41),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_91),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_58),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_116),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_136),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_14),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_37),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_138),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_24),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_82),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_110),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_160),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_25),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_130),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_143),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_13),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_29),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_21),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_159),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_124),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_6),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_31),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_26),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_4),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_84),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_61),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_35),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_99),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_19),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_108),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_167),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_153),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_3),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_33),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_3),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_32),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_20),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_164),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_150),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_254),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_169),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

BUFx2_ASAP7_75t_SL g349 ( 
.A(n_193),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_172),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_197),
.B(n_1),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_200),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_206),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_241),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_207),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_205),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_250),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_175),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_172),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_210),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_1),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_211),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_295),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_175),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_213),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_193),
.B(n_6),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_175),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_191),
.B(n_7),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_183),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_216),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_220),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_181),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_257),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_229),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_191),
.B(n_8),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_196),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_257),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_175),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_221),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_232),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_196),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_233),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_239),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_240),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_175),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_257),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_208),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_208),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_257),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_288),
.B(n_9),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_219),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_208),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_208),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_261),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_261),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_244),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_294),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_223),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_262),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_245),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_178),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_294),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_246),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_309),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_288),
.B(n_17),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_182),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_248),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_260),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_272),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_333),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_274),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_332),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_225),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_276),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_186),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_194),
.B(n_18),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_278),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_281),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_195),
.B(n_20),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_353),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_345),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_376),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_R g439 ( 
.A(n_379),
.B(n_171),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_387),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_359),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_366),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_368),
.B(n_219),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_407),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_350),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_395),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_408),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_413),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_378),
.B(n_342),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_422),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_381),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_382),
.B(n_342),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_385),
.B(n_170),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_173),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_360),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_351),
.A2(n_247),
.B1(n_292),
.B2(n_290),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_400),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_349),
.B(n_171),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_365),
.B(n_338),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_402),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_385),
.B(n_257),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_390),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_391),
.Y(n_484)
);

INVx6_ASAP7_75t_L g485 ( 
.A(n_350),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_346),
.A2(n_348),
.B(n_347),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_426),
.B(n_275),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_369),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_346),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_385),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_384),
.B(n_202),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_347),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_348),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_392),
.B(n_179),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_369),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_415),
.B(n_202),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_405),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_352),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_352),
.Y(n_504)
);

BUFx8_ASAP7_75t_L g505 ( 
.A(n_350),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_409),
.B(n_184),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_453),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_434),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_489),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_445),
.B(n_412),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_453),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_488),
.A2(n_362),
.B1(n_357),
.B2(n_427),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_389),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_459),
.B(n_417),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_488),
.A2(n_374),
.B1(n_398),
.B2(n_383),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_497),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_465),
.B(n_418),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_468),
.B(n_419),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_421),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_431),
.B(n_344),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_498),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_469),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_504),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_503),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_L g529 ( 
.A(n_481),
.B(n_275),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_503),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_399),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_436),
.B(n_424),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_485),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_428),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_478),
.A2(n_414),
.B1(n_372),
.B2(n_349),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_495),
.B(n_358),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_432),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_485),
.B(n_354),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_442),
.B(n_429),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_495),
.B(n_403),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_476),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_450),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_433),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_485),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g549 ( 
.A(n_451),
.B(n_275),
.Y(n_549)
);

AND2x2_ASAP7_75t_SL g550 ( 
.A(n_474),
.B(n_275),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_442),
.B(n_202),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_441),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_487),
.A2(n_367),
.B1(n_192),
.B2(n_321),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_479),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_480),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_462),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_444),
.B(n_256),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_503),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_444),
.B(n_256),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_485),
.B(n_354),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_440),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_494),
.B(n_356),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_505),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_471),
.B(n_410),
.C(n_367),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_462),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_403),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_494),
.B(n_356),
.Y(n_573)
);

BUFx8_ASAP7_75t_SL g574 ( 
.A(n_474),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_463),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_463),
.Y(n_576)
);

AND2x2_ASAP7_75t_SL g577 ( 
.A(n_494),
.B(n_189),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_501),
.B(n_203),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_454),
.B(n_425),
.Y(n_581)
);

INVx4_ASAP7_75t_SL g582 ( 
.A(n_481),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_454),
.B(n_256),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_448),
.Y(n_584)
);

AND2x2_ASAP7_75t_SL g585 ( 
.A(n_493),
.B(n_199),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_466),
.B(n_234),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_441),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_505),
.B(n_252),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_441),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_448),
.B(n_404),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_439),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_461),
.A2(n_502),
.B1(n_484),
.B2(n_483),
.Y(n_594)
);

NOR3xp33_ASAP7_75t_L g595 ( 
.A(n_461),
.B(n_484),
.C(n_483),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_467),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g597 ( 
.A(n_441),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_473),
.B(n_361),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_496),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_481),
.A2(n_317),
.B1(n_280),
.B2(n_284),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_493),
.B(n_361),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_456),
.B(n_363),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_502),
.B(n_174),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_456),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_500),
.B(n_174),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_447),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_486),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_490),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_490),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_464),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_464),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_491),
.B(n_425),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_491),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_464),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_470),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_457),
.B(n_176),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_470),
.B(n_404),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_481),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_481),
.A2(n_277),
.B1(n_287),
.B2(n_341),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_470),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_470),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_470),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_482),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_482),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_482),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_458),
.B(n_209),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_460),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_453),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_475),
.B(n_283),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_434),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_487),
.Y(n_637)
);

OAI221xp5_ASAP7_75t_L g638 ( 
.A1(n_471),
.A2(n_339),
.B1(n_337),
.B2(n_297),
.C(n_406),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_488),
.A2(n_286),
.B1(n_285),
.B2(n_201),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

NOR2x1p5_ASAP7_75t_L g641 ( 
.A(n_431),
.B(n_187),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_481),
.B(n_212),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_503),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_577),
.B(n_224),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_637),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_510),
.B(n_226),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_540),
.B(n_187),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_513),
.B(n_406),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_549),
.B(n_176),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_572),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_514),
.B(n_227),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_599),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_520),
.B(n_235),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_549),
.B(n_177),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_577),
.A2(n_291),
.B1(n_305),
.B2(n_325),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_581),
.B(n_177),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_513),
.A2(n_296),
.B1(n_301),
.B2(n_302),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_637),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_518),
.A2(n_242),
.B1(n_238),
.B2(n_236),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_526),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_517),
.B(n_249),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_517),
.B(n_251),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_519),
.B(n_255),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_568),
.A2(n_258),
.B(n_259),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_637),
.B(n_265),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_593),
.B(n_526),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_581),
.B(n_180),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_637),
.B(n_303),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_266),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_572),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_553),
.A2(n_293),
.B1(n_343),
.B2(n_289),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_525),
.B(n_269),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_525),
.B(n_300),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_540),
.B(n_198),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_508),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_507),
.B(n_411),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_527),
.B(n_306),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_527),
.B(n_329),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_550),
.B(n_180),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_592),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_531),
.B(n_185),
.Y(n_682)
);

O2A1O1Ixp5_ASAP7_75t_L g683 ( 
.A1(n_560),
.A2(n_335),
.B(n_330),
.C(n_411),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_544),
.B(n_420),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_531),
.B(n_521),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_640),
.B(n_307),
.Y(n_686)
);

BUFx8_ASAP7_75t_L g687 ( 
.A(n_633),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_640),
.A2(n_308),
.B(n_336),
.C(n_334),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_523),
.B(n_185),
.Y(n_689)
);

NAND2x1_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_416),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_537),
.B(n_188),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_596),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_511),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_560),
.A2(n_318),
.B(n_336),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_512),
.B(n_188),
.Y(n_695)
);

OAI221xp5_ASAP7_75t_L g696 ( 
.A1(n_539),
.A2(n_638),
.B1(n_570),
.B2(n_639),
.C(n_614),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_550),
.B(n_190),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_511),
.B(n_635),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_634),
.B(n_312),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_544),
.B(n_215),
.C(n_217),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_543),
.B(n_312),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_596),
.B(n_314),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_604),
.B(n_632),
.C(n_595),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_535),
.B(n_314),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_535),
.B(n_315),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_524),
.B(n_522),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_580),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_579),
.A2(n_198),
.B1(n_340),
.B2(n_264),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_594),
.B(n_315),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_606),
.B(n_264),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_536),
.B(n_316),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_536),
.B(n_316),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_538),
.B(n_416),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_538),
.B(n_318),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_545),
.B(n_319),
.Y(n_715)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_632),
.A2(n_340),
.B1(n_310),
.B2(n_331),
.C(n_328),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_545),
.B(n_319),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_522),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_580),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_637),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_556),
.B(n_323),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_573),
.A2(n_566),
.B(n_542),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_551),
.B(n_323),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_585),
.B(n_324),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_556),
.B(n_324),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_585),
.A2(n_310),
.B1(n_331),
.B2(n_328),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_586),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_589),
.B(n_22),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_522),
.B(n_204),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_574),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_515),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_584),
.A2(n_311),
.B1(n_326),
.B2(n_322),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_533),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_532),
.B(n_334),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_557),
.B(n_214),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_516),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_584),
.A2(n_326),
.B1(n_322),
.B2(n_320),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_557),
.B(n_268),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_579),
.A2(n_270),
.B1(n_222),
.B2(n_304),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_558),
.B(n_267),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_562),
.B(n_271),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_579),
.A2(n_263),
.B1(n_230),
.B2(n_299),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_565),
.B(n_273),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_533),
.B(n_253),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_548),
.B(n_87),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_548),
.B(n_279),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_563),
.B(n_243),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_586),
.A2(n_298),
.B1(n_282),
.B2(n_237),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_614),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_563),
.B(n_231),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_597),
.A2(n_218),
.B(n_320),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_622),
.B(n_311),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_641),
.B(n_23),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_564),
.B(n_621),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_586),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_620),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_588),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_583),
.B(n_24),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_622),
.B(n_76),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_586),
.A2(n_65),
.B1(n_166),
.B2(n_162),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_621),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_554),
.B(n_52),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_541),
.B(n_27),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_608),
.B(n_77),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_547),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_567),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_618),
.B(n_168),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_618),
.B(n_149),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_609),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_569),
.B(n_578),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_574),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_534),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_633),
.B(n_30),
.C(n_32),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_600),
.B(n_30),
.C(n_34),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_528),
.A2(n_643),
.B1(n_530),
.B2(n_616),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_615),
.B(n_106),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_625),
.B(n_104),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_569),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_615),
.B(n_103),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_607),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_615),
.B(n_88),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_615),
.B(n_34),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_578),
.B(n_36),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_530),
.B(n_36),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_530),
.B(n_643),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_643),
.A2(n_626),
.B1(n_589),
.B2(n_624),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_703),
.B(n_589),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_692),
.B(n_589),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_718),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_685),
.B(n_626),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_772),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_666),
.B(n_509),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_685),
.B(n_624),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_769),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_698),
.B(n_617),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_658),
.A2(n_631),
.B(n_603),
.Y(n_796)
);

AOI21x1_ASAP7_75t_L g797 ( 
.A1(n_690),
.A2(n_628),
.B(n_598),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_612),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_656),
.B(n_612),
.Y(n_799)
);

AO21x1_ASAP7_75t_L g800 ( 
.A1(n_644),
.A2(n_628),
.B(n_602),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_675),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_720),
.A2(n_630),
.B(n_613),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_645),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_656),
.B(n_591),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_659),
.A2(n_623),
.B1(n_590),
.B2(n_587),
.Y(n_805)
);

BUFx4f_ASAP7_75t_L g806 ( 
.A(n_770),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_646),
.B(n_552),
.Y(n_807)
);

NOR3xp33_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_642),
.C(n_529),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_651),
.B(n_653),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_683),
.A2(n_576),
.B(n_636),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_667),
.B(n_590),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_707),
.B(n_719),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_SL g813 ( 
.A1(n_644),
.A2(n_576),
.B(n_636),
.C(n_575),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_761),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_706),
.B(n_615),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_765),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_587),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_645),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_720),
.A2(n_601),
.B(n_627),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_720),
.A2(n_627),
.B(n_588),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_645),
.A2(n_627),
.B(n_588),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_648),
.B(n_605),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_645),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_785),
.A2(n_627),
.B(n_588),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_694),
.A2(n_610),
.B(n_642),
.C(n_561),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_695),
.A2(n_561),
.B(n_555),
.C(n_546),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_687),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_689),
.B(n_582),
.Y(n_828)
);

AOI22x1_ASAP7_75t_SL g829 ( 
.A1(n_749),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_696),
.A2(n_610),
.B(n_575),
.C(n_591),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_733),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_659),
.A2(n_559),
.B(n_546),
.C(n_555),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_676),
.B(n_691),
.Y(n_833)
);

NOR2x1_ASAP7_75t_L g834 ( 
.A(n_693),
.B(n_611),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_733),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_785),
.A2(n_588),
.B(n_601),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_766),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_665),
.A2(n_601),
.B(n_619),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_665),
.A2(n_754),
.B(n_722),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_759),
.A2(n_559),
.B(n_571),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_668),
.A2(n_601),
.B(n_619),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_733),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_780),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_650),
.B(n_629),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_670),
.B(n_582),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_713),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_757),
.A2(n_582),
.B(n_44),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_741),
.A2(n_51),
.B(n_45),
.C(n_46),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_745),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_682),
.B(n_43),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_671),
.A2(n_50),
.B(n_680),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_756),
.B(n_681),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_684),
.B(n_682),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_763),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_671),
.B(n_745),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_655),
.A2(n_786),
.B1(n_649),
.B2(n_654),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_723),
.B(n_699),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_713),
.Y(n_858)
);

BUFx4f_ASAP7_75t_L g859 ( 
.A(n_728),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_655),
.A2(n_697),
.B1(n_679),
.B2(n_775),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_744),
.A2(n_746),
.B(n_747),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_758),
.A2(n_723),
.B(n_724),
.C(n_755),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_702),
.B(n_661),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_758),
.A2(n_737),
.B1(n_732),
.B2(n_726),
.Y(n_864)
);

INVx11_ASAP7_75t_L g865 ( 
.A(n_687),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_699),
.B(n_709),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_724),
.A2(n_752),
.B(n_782),
.C(n_688),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_776),
.B(n_779),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_729),
.B(n_647),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_750),
.A2(n_686),
.B(n_764),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_767),
.A2(n_768),
.B(n_777),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_752),
.A2(n_782),
.B(n_708),
.C(n_677),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_664),
.A2(n_700),
.B(n_784),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_662),
.B(n_672),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_663),
.B(n_678),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_731),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_784),
.A2(n_673),
.B(n_669),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_735),
.B(n_738),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_701),
.B(n_710),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_736),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_674),
.B(n_727),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_652),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_740),
.A2(n_762),
.B(n_751),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_704),
.B(n_715),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_657),
.B(n_734),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_753),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_781),
.A2(n_705),
.B(n_721),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_727),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_711),
.A2(n_725),
.B(n_712),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_714),
.A2(n_717),
.B1(n_743),
.B2(n_760),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_708),
.A2(n_783),
.B(n_748),
.C(n_774),
.Y(n_891)
);

AOI21xp33_ASAP7_75t_L g892 ( 
.A1(n_739),
.A2(n_742),
.B(n_716),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_732),
.A2(n_737),
.B(n_726),
.Y(n_893)
);

BUFx8_ASAP7_75t_SL g894 ( 
.A(n_730),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_773),
.A2(n_728),
.B(n_778),
.C(n_771),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_773),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_685),
.B(n_698),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_685),
.B(n_698),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_685),
.A2(n_646),
.B(n_653),
.C(n_651),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_644),
.A2(n_665),
.B(n_694),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_685),
.B(n_698),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_905)
);

NOR2x1p5_ASAP7_75t_SL g906 ( 
.A(n_675),
.B(n_560),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_769),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_666),
.B(n_685),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_685),
.B(n_593),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_660),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_769),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_685),
.B(n_593),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_659),
.A2(n_696),
.B1(n_518),
.B2(n_651),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_683),
.A2(n_560),
.B(n_487),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_685),
.A2(n_646),
.B(n_653),
.C(n_651),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_659),
.A2(n_696),
.B1(n_518),
.B2(n_651),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_666),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_659),
.A2(n_696),
.B1(n_518),
.B2(n_651),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_685),
.B(n_698),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_685),
.B(n_593),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_660),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_659),
.A2(n_696),
.B1(n_518),
.B2(n_651),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_685),
.B(n_698),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_683),
.A2(n_560),
.B(n_487),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_685),
.B(n_698),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_645),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_685),
.B(n_698),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_685),
.B(n_698),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_685),
.B(n_593),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_685),
.B(n_593),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_685),
.B(n_593),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_658),
.A2(n_720),
.B(n_637),
.Y(n_936)
);

OAI321xp33_ASAP7_75t_L g937 ( 
.A1(n_659),
.A2(n_518),
.A3(n_758),
.B1(n_708),
.B2(n_696),
.C(n_694),
.Y(n_937)
);

AND2x6_ASAP7_75t_L g938 ( 
.A(n_645),
.B(n_786),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_685),
.B(n_698),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_685),
.B(n_698),
.Y(n_940)
);

AO21x2_ASAP7_75t_L g941 ( 
.A1(n_839),
.A2(n_877),
.B(n_873),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_831),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_897),
.B(n_898),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_797),
.A2(n_838),
.B(n_841),
.Y(n_944)
);

AOI21xp33_ASAP7_75t_L g945 ( 
.A1(n_857),
.A2(n_919),
.B(n_914),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_900),
.A2(n_904),
.B(n_902),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_866),
.A2(n_893),
.B(n_937),
.C(n_892),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_921),
.A2(n_925),
.B(n_937),
.Y(n_948)
);

NAND3xp33_ASAP7_75t_L g949 ( 
.A(n_903),
.B(n_928),
.C(n_922),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_930),
.B(n_931),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_939),
.B(n_940),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_905),
.A2(n_917),
.B(n_907),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_821),
.A2(n_927),
.B(n_915),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_918),
.A2(n_936),
.B(n_934),
.Y(n_954)
);

OAI211xp5_ASAP7_75t_SL g955 ( 
.A1(n_920),
.A2(n_893),
.B(n_854),
.C(n_852),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_853),
.B(n_910),
.Y(n_956)
);

OAI22x1_ASAP7_75t_L g957 ( 
.A1(n_896),
.A2(n_879),
.B1(n_932),
.B2(n_923),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_913),
.B(n_933),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_935),
.B(n_926),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_909),
.B(n_869),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_833),
.B(n_806),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_810),
.A2(n_840),
.B(n_796),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_816),
.B(n_911),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_809),
.B(n_878),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_871),
.A2(n_875),
.B(n_874),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_864),
.A2(n_856),
.B1(n_860),
.B2(n_890),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_887),
.A2(n_861),
.B(n_870),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_864),
.A2(n_855),
.B1(n_851),
.B2(n_849),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_831),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_819),
.A2(n_820),
.B(n_802),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_806),
.B(n_816),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_851),
.B(n_815),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_867),
.A2(n_873),
.B(n_872),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_794),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_899),
.A2(n_916),
.B(n_830),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_884),
.B(n_804),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_850),
.A2(n_885),
.B1(n_886),
.B2(n_787),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_790),
.B(n_793),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_863),
.A2(n_807),
.B(n_822),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_832),
.A2(n_826),
.B(n_862),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_849),
.A2(n_812),
.B1(n_868),
.B2(n_912),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_924),
.B(n_843),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_831),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_848),
.A2(n_891),
.B(n_881),
.C(n_886),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_849),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_854),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_849),
.B(n_795),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_815),
.A2(n_883),
.B(n_811),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_792),
.A2(n_858),
.B1(n_846),
.B2(n_938),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_842),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_883),
.A2(n_817),
.B(n_828),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_789),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_803),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_825),
.A2(n_805),
.B(n_889),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_803),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_837),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_844),
.A2(n_845),
.B(n_929),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_908),
.B(n_814),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_888),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_818),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_823),
.A2(n_929),
.B(n_813),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_823),
.A2(n_842),
.B(n_835),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_798),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_938),
.B(n_858),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_827),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_788),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_938),
.B(n_882),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_808),
.A2(n_880),
.B(n_801),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_876),
.A2(n_834),
.B(n_847),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_788),
.A2(n_859),
.B(n_895),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_906),
.B(n_829),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_865),
.A2(n_839),
.B(n_914),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_894),
.A2(n_797),
.B(n_838),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_857),
.B(n_853),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_909),
.B(n_666),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_839),
.A2(n_836),
.B(n_824),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_897),
.B(n_898),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_791),
.Y(n_1019)
);

INVx3_ASAP7_75t_SL g1020 ( 
.A(n_837),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_831),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_853),
.B(n_703),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_897),
.B(n_898),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_909),
.B(n_666),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_849),
.B(n_842),
.Y(n_1028)
);

CKINVDCx16_ASAP7_75t_R g1029 ( 
.A(n_792),
.Y(n_1029)
);

AND2x6_ASAP7_75t_L g1030 ( 
.A(n_855),
.B(n_787),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_897),
.B(n_898),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_791),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_897),
.B(n_898),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_849),
.B(n_645),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_794),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_L g1036 ( 
.A1(n_857),
.A2(n_866),
.B1(n_896),
.B2(n_879),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_788),
.B(n_846),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_897),
.B(n_898),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_849),
.B(n_842),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_857),
.B(n_897),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_900),
.A2(n_720),
.B(n_658),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_797),
.A2(n_838),
.B(n_841),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_900),
.A2(n_720),
.B(n_658),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_897),
.B(n_898),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_788),
.B(n_846),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_909),
.B(n_666),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1047)
);

INVx6_ASAP7_75t_L g1048 ( 
.A(n_827),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_897),
.B(n_898),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_897),
.B(n_898),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_827),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_900),
.A2(n_720),
.B(n_658),
.Y(n_1052)
);

BUFx4_ASAP7_75t_SL g1053 ( 
.A(n_837),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_900),
.A2(n_720),
.B(n_658),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_897),
.B(n_898),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_794),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_797),
.A2(n_838),
.B(n_841),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_911),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_839),
.A2(n_919),
.B(n_914),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_791),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_900),
.A2(n_720),
.B(n_658),
.Y(n_1062)
);

AO31x2_ASAP7_75t_L g1063 ( 
.A1(n_901),
.A2(n_800),
.A3(n_919),
.B(n_914),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_909),
.B(n_666),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_797),
.A2(n_838),
.B(n_841),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_965),
.A2(n_967),
.B(n_988),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1040),
.B(n_964),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_960),
.B(n_1015),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_964),
.A2(n_991),
.B(n_979),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_943),
.B(n_1031),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_958),
.A2(n_966),
.B(n_947),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_1010),
.B(n_982),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1029),
.A2(n_972),
.B1(n_961),
.B2(n_1003),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_993),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_943),
.B(n_1031),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_963),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_993),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_972),
.B1(n_948),
.B2(n_1024),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_1028),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1033),
.B(n_1055),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1027),
.B(n_1046),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1035),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1058),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_1051),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1056),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_975),
.A2(n_1021),
.B(n_1018),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1064),
.B(n_1003),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1033),
.B(n_1055),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1018),
.A2(n_1023),
.B(n_1021),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_945),
.A2(n_948),
.B1(n_973),
.B2(n_1036),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1023),
.A2(n_1047),
.B(n_1060),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_982),
.B(n_971),
.Y(n_1092)
);

INVx3_ASAP7_75t_SL g1093 ( 
.A(n_992),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_994),
.A2(n_1034),
.B(n_952),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_994),
.A2(n_954),
.B(n_946),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_950),
.B(n_951),
.Y(n_1096)
);

INVx3_ASAP7_75t_SL g1097 ( 
.A(n_1020),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1014),
.B(n_1026),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_998),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_956),
.B(n_1017),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_976),
.B(n_986),
.Y(n_1101)
);

CKINVDCx8_ASAP7_75t_R g1102 ( 
.A(n_996),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1025),
.A2(n_1059),
.B(n_1047),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_993),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_1005),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_982),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1053),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1038),
.B(n_1044),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_995),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1005),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_999),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_942),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1025),
.A2(n_1060),
.B(n_1059),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_959),
.B(n_957),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_941),
.A2(n_980),
.B(n_978),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_984),
.A2(n_1012),
.B(n_1049),
.C(n_1050),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1012),
.A2(n_949),
.B(n_977),
.C(n_968),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_949),
.B(n_1006),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_968),
.B(n_1030),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_1004),
.B(n_1028),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_955),
.A2(n_1011),
.B(n_981),
.C(n_985),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1019),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_941),
.A2(n_981),
.B(n_987),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1032),
.B(n_1061),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1030),
.A2(n_1004),
.B1(n_989),
.B2(n_1007),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1030),
.B(n_1063),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1030),
.B(n_1063),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_942),
.Y(n_1130)
);

AND2x2_ASAP7_75t_SL g1131 ( 
.A(n_1022),
.B(n_942),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_969),
.B(n_983),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_995),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_1008),
.A2(n_1039),
.B(n_997),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_969),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_L g1136 ( 
.A(n_1048),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_983),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_995),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1039),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1022),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_1000),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1000),
.B(n_1063),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1013),
.B(n_1009),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1048),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_970),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_953),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1001),
.A2(n_962),
.B1(n_1065),
.B2(n_944),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_1016),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1042),
.A2(n_1057),
.B(n_1043),
.C(n_1052),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1041),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1054),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1062),
.A2(n_1040),
.B1(n_947),
.B2(n_964),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_963),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_960),
.B(n_1015),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1040),
.A2(n_857),
.B1(n_866),
.B2(n_376),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1040),
.B(n_964),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1040),
.B(n_857),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_942),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_964),
.B(n_963),
.Y(n_1161)
);

CKINVDCx11_ASAP7_75t_R g1162 ( 
.A(n_1051),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_963),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1040),
.B(n_964),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_960),
.B(n_1015),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_974),
.Y(n_1166)
);

BUFx4f_ASAP7_75t_L g1167 ( 
.A(n_1020),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1040),
.A2(n_706),
.B1(n_857),
.B2(n_864),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1040),
.A2(n_947),
.B1(n_964),
.B2(n_966),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1058),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1040),
.B(n_964),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_992),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_960),
.B(n_1015),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1040),
.B(n_964),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_964),
.B(n_963),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1040),
.A2(n_947),
.B1(n_964),
.B2(n_966),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_990),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_942),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1040),
.B(n_964),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_960),
.B(n_1015),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1058),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_958),
.A2(n_857),
.B(n_947),
.C(n_864),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1058),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1003),
.B(n_964),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1040),
.B(n_964),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_974),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_942),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_963),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1072),
.B(n_1111),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1158),
.A2(n_1156),
.B1(n_1168),
.B2(n_1108),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1181),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1166),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1072),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1067),
.A2(n_1171),
.B1(n_1179),
.B2(n_1174),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1186),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1083),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1072),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1082),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1070),
.B(n_1075),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1070),
.B(n_1075),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1080),
.B(n_1088),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1100),
.B(n_1067),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1085),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1143),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1113),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1071),
.A2(n_1169),
.B1(n_1176),
.B2(n_1116),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1083),
.Y(n_1208)
);

NAND2x1_ASAP7_75t_L g1209 ( 
.A(n_1079),
.B(n_1139),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_R g1210 ( 
.A(n_1157),
.B(n_1164),
.Y(n_1210)
);

CKINVDCx8_ASAP7_75t_R g1211 ( 
.A(n_1172),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1157),
.B(n_1164),
.Y(n_1212)
);

AO21x2_ASAP7_75t_L g1213 ( 
.A1(n_1095),
.A2(n_1066),
.B(n_1094),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1169),
.A2(n_1176),
.B1(n_1103),
.B2(n_1115),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1152),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1170),
.Y(n_1216)
);

BUFx12f_ASAP7_75t_L g1217 ( 
.A(n_1162),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1183),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1171),
.B(n_1174),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1133),
.Y(n_1220)
);

AO21x1_ASAP7_75t_SL g1221 ( 
.A1(n_1128),
.A2(n_1129),
.B(n_1121),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1179),
.A2(n_1185),
.B1(n_1096),
.B2(n_1088),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1163),
.Y(n_1223)
);

INVxp33_ASAP7_75t_L g1224 ( 
.A(n_1081),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1124),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1163),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1099),
.Y(n_1227)
);

CKINVDCx6p67_ASAP7_75t_R g1228 ( 
.A(n_1093),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1185),
.B(n_1096),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1080),
.B(n_1098),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1126),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1102),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1076),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1152),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1115),
.A2(n_1078),
.B1(n_1091),
.B2(n_1089),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1092),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1161),
.B(n_1175),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1120),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1125),
.A2(n_1119),
.B(n_1086),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1092),
.Y(n_1240)
);

BUFx8_ASAP7_75t_L g1241 ( 
.A(n_1084),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1122),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1089),
.A2(n_1091),
.B1(n_1086),
.B2(n_1087),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1135),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1068),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1137),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1184),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1105),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1149),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1149),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1138),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1090),
.B(n_1118),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1101),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1155),
.B(n_1165),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1073),
.A2(n_1092),
.B1(n_1127),
.B2(n_1182),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1173),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1154),
.A2(n_1189),
.B1(n_1167),
.B2(n_1097),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1180),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1132),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1130),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1167),
.A2(n_1121),
.B1(n_1153),
.B2(n_1136),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1153),
.B(n_1122),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1188),
.B(n_1160),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1112),
.Y(n_1264)
);

BUFx4_ASAP7_75t_R g1265 ( 
.A(n_1145),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1177),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1114),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1131),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1106),
.A2(n_1123),
.B1(n_1122),
.B2(n_1117),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1069),
.A2(n_1117),
.B(n_1128),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1111),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1074),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1187),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1074),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1147),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1146),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1110),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1150),
.A2(n_1148),
.B(n_1129),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1136),
.A2(n_1140),
.B1(n_1139),
.B2(n_1187),
.Y(n_1279)
);

BUFx4f_ASAP7_75t_L g1280 ( 
.A(n_1077),
.Y(n_1280)
);

NAND2x1_ASAP7_75t_L g1281 ( 
.A(n_1144),
.B(n_1141),
.Y(n_1281)
);

AO21x1_ASAP7_75t_L g1282 ( 
.A1(n_1151),
.A2(n_1142),
.B(n_1134),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1141),
.B(n_1159),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1077),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1104),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1159),
.B(n_1178),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1104),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1109),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1109),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1107),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1221),
.Y(n_1291)
);

CKINVDCx16_ASAP7_75t_R g1292 ( 
.A(n_1217),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1221),
.B(n_1243),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1213),
.A2(n_1282),
.B(n_1269),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1239),
.B(n_1235),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1239),
.B(n_1205),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1200),
.B(n_1201),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1213),
.A2(n_1282),
.B(n_1278),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1236),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1242),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1239),
.B(n_1262),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1275),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1191),
.A2(n_1214),
.B(n_1207),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1230),
.B(n_1262),
.Y(n_1304)
);

OR2x6_ASAP7_75t_L g1305 ( 
.A(n_1194),
.B(n_1198),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1270),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1194),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1230),
.B(n_1252),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1240),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1198),
.B(n_1281),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1252),
.A2(n_1255),
.B1(n_1261),
.B2(n_1240),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1238),
.Y(n_1312)
);

BUFx2_ASAP7_75t_R g1313 ( 
.A(n_1211),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1270),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1213),
.A2(n_1278),
.B(n_1249),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1200),
.B(n_1201),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1242),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1202),
.B(n_1278),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1250),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1242),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1227),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1199),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1204),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_1217),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1247),
.B(n_1276),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1222),
.A2(n_1203),
.B(n_1195),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1276),
.B(n_1244),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1246),
.A2(n_1225),
.B(n_1266),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1193),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1210),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1210),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1226),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1190),
.B(n_1215),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1234),
.B(n_1224),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1237),
.B(n_1226),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1224),
.B(n_1229),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1231),
.B(n_1212),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1223),
.B(n_1253),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1219),
.A2(n_1190),
.B(n_1279),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1190),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1197),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1268),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1259),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1260),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1251),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1268),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1305),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1304),
.B(n_1256),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1318),
.B(n_1245),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1304),
.B(n_1258),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1318),
.B(n_1254),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1318),
.B(n_1267),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1301),
.B(n_1287),
.Y(n_1354)
);

NOR2x1_ASAP7_75t_L g1355 ( 
.A(n_1326),
.B(n_1257),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1344),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1301),
.B(n_1208),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1303),
.A2(n_1192),
.B(n_1271),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1296),
.B(n_1288),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1291),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1292),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1296),
.B(n_1288),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_SL g1363 ( 
.A(n_1310),
.B(n_1273),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1296),
.B(n_1233),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1310),
.B(n_1291),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1310),
.B(n_1263),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1330),
.B(n_1216),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1330),
.B(n_1216),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1310),
.B(n_1263),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_R g1370 ( 
.A(n_1313),
.B(n_1277),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1328),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1331),
.B(n_1218),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_1339),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1328),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1328),
.Y(n_1375)
);

AND2x4_ASAP7_75t_SL g1376 ( 
.A(n_1317),
.B(n_1228),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1303),
.A2(n_1232),
.B1(n_1263),
.B2(n_1228),
.Y(n_1377)
);

NAND4xp25_ASAP7_75t_L g1378 ( 
.A(n_1326),
.B(n_1264),
.C(n_1232),
.D(n_1218),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1331),
.B(n_1300),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1328),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1316),
.B(n_1308),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1302),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1340),
.B(n_1211),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1344),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1322),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1305),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1305),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1308),
.B(n_1272),
.Y(n_1388)
);

OAI21xp33_ASAP7_75t_L g1389 ( 
.A1(n_1311),
.A2(n_1283),
.B(n_1286),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1308),
.B(n_1285),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_L g1391 ( 
.A(n_1340),
.B(n_1209),
.C(n_1289),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1293),
.B(n_1274),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1293),
.B(n_1335),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1293),
.B(n_1284),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1352),
.B(n_1333),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1393),
.B(n_1295),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1355),
.B(n_1307),
.C(n_1335),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_SL g1398 ( 
.A(n_1370),
.B(n_1313),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1393),
.B(n_1352),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1357),
.B(n_1333),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1358),
.A2(n_1347),
.B1(n_1343),
.B2(n_1295),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_L g1402 ( 
.A1(n_1355),
.A2(n_1337),
.B(n_1295),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1383),
.B(n_1334),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1378),
.A2(n_1334),
.B1(n_1341),
.B2(n_1305),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1391),
.B(n_1334),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1377),
.A2(n_1339),
.B1(n_1336),
.B2(n_1337),
.C(n_1342),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1357),
.B(n_1336),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1364),
.B(n_1342),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_L g1409 ( 
.A(n_1389),
.B(n_1307),
.C(n_1335),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1389),
.B(n_1345),
.C(n_1312),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1363),
.A2(n_1347),
.B1(n_1343),
.B2(n_1317),
.Y(n_1411)
);

NOR3xp33_ASAP7_75t_SL g1412 ( 
.A(n_1371),
.B(n_1324),
.C(n_1292),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1361),
.B(n_1334),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1373),
.A2(n_1343),
.B1(n_1347),
.B2(n_1324),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1363),
.A2(n_1320),
.B(n_1317),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1354),
.B(n_1315),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1364),
.B(n_1312),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1371),
.A2(n_1314),
.B(n_1306),
.Y(n_1418)
);

OAI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1367),
.A2(n_1299),
.B1(n_1309),
.B2(n_1341),
.C(n_1345),
.Y(n_1419)
);

NAND2xp33_ASAP7_75t_SL g1420 ( 
.A(n_1367),
.B(n_1317),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1350),
.B(n_1297),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1359),
.B(n_1294),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1368),
.B(n_1329),
.C(n_1332),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1368),
.B(n_1325),
.C(n_1327),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1350),
.B(n_1297),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1359),
.B(n_1294),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1381),
.B(n_1356),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1381),
.B(n_1325),
.Y(n_1428)
);

NAND3xp33_ASAP7_75t_L g1429 ( 
.A(n_1372),
.B(n_1325),
.C(n_1327),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1384),
.B(n_1319),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1373),
.A2(n_1265),
.B1(n_1290),
.B2(n_1277),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1372),
.B(n_1319),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1353),
.B(n_1319),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1392),
.A2(n_1341),
.B1(n_1309),
.B2(n_1299),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1353),
.B(n_1346),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1385),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1392),
.A2(n_1341),
.B1(n_1309),
.B2(n_1299),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1351),
.B(n_1346),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1348),
.A2(n_1320),
.B1(n_1317),
.B2(n_1294),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1362),
.B(n_1294),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1351),
.B(n_1338),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1349),
.B(n_1338),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1349),
.B(n_1302),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.B(n_1298),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1394),
.B(n_1323),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1382),
.B(n_1321),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1397),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1399),
.B(n_1365),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1399),
.B(n_1365),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1422),
.B(n_1374),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1436),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1396),
.B(n_1365),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1396),
.B(n_1365),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1436),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1446),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1444),
.B(n_1348),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1423),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1423),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1410),
.A2(n_1379),
.B1(n_1390),
.B2(n_1388),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1430),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1418),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1422),
.B(n_1374),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1432),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1400),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1418),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1426),
.B(n_1375),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1426),
.B(n_1375),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1416),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1418),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1440),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1435),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1440),
.B(n_1386),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1433),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1427),
.B(n_1395),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1438),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1445),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1443),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1408),
.B(n_1380),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1407),
.B(n_1417),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1439),
.B(n_1387),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1420),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1428),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1455),
.B(n_1402),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1457),
.B(n_1458),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1451),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1479),
.B(n_1421),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1451),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1454),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1490)
);

NOR2x1p5_ASAP7_75t_SL g1491 ( 
.A(n_1469),
.B(n_1380),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1454),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1457),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1458),
.B(n_1425),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1453),
.B(n_1387),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1481),
.B(n_1402),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1479),
.B(n_1442),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1482),
.B(n_1424),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1481),
.B(n_1360),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1460),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1482),
.B(n_1475),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1475),
.B(n_1429),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1460),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1448),
.B(n_1379),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1419),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1463),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1448),
.B(n_1360),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1463),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1464),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1476),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1449),
.B(n_1480),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1476),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1467),
.B(n_1410),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1474),
.Y(n_1515)
);

NOR2x1_ASAP7_75t_L g1516 ( 
.A(n_1459),
.B(n_1405),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1461),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1467),
.B(n_1409),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1478),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1465),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1449),
.B(n_1360),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1486),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1488),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1516),
.A2(n_1447),
.B(n_1403),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1493),
.B(n_1447),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1485),
.B(n_1478),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1485),
.B(n_1450),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1514),
.B(n_1450),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1514),
.B(n_1462),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1489),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1462),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1520),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1520),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1471),
.Y(n_1534)
);

AOI21xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1496),
.A2(n_1431),
.B(n_1459),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1518),
.B(n_1466),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1519),
.B(n_1466),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1471),
.Y(n_1538)
);

NOR3x1_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1414),
.C(n_1413),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1492),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1513),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1503),
.B(n_1468),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1494),
.B(n_1477),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1510),
.B(n_1477),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1496),
.B(n_1470),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1501),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1515),
.B(n_1474),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1473),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1502),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1484),
.A2(n_1480),
.B(n_1401),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1500),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1500),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1504),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1507),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1499),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1472),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1512),
.A2(n_1369),
.B1(n_1366),
.B2(n_1404),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1487),
.B(n_1473),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1509),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1562)
);

AND2x2_ASAP7_75t_SL g1563 ( 
.A(n_1512),
.B(n_1398),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1490),
.B(n_1456),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1540),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1540),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1525),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1563),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1563),
.B(n_1505),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1556),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1522),
.Y(n_1573)
);

AOI222xp33_ASAP7_75t_L g1574 ( 
.A1(n_1552),
.A2(n_1431),
.B1(n_1517),
.B2(n_1370),
.C1(n_1491),
.C2(n_1420),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1557),
.B(n_1490),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1524),
.B(n_1495),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1558),
.B(n_1505),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1554),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1517),
.C(n_1406),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1550),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1558),
.B(n_1550),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1561),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1553),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1546),
.B(n_1505),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1546),
.B(n_1508),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1538),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1561),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1415),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1539),
.B(n_1508),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1551),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1541),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1526),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1532),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1523),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1534),
.B(n_1495),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1241),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1551),
.B(n_1456),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1526),
.B(n_1241),
.C(n_1461),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1544),
.B(n_1549),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_R g1602 ( 
.A(n_1568),
.B(n_1248),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1531),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1579),
.A2(n_1559),
.B1(n_1536),
.B2(n_1531),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1574),
.A2(n_1567),
.B(n_1590),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1572),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1599),
.A2(n_1547),
.B(n_1542),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1597),
.B(n_1241),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1576),
.A2(n_1564),
.B1(n_1562),
.B2(n_1536),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1590),
.A2(n_1528),
.B1(n_1529),
.B2(n_1376),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1586),
.B(n_1578),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1569),
.A2(n_1555),
.B1(n_1530),
.B2(n_1545),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1581),
.B(n_1521),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1599),
.A2(n_1593),
.B(n_1595),
.C(n_1583),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1543),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1560),
.Y(n_1618)
);

OAI21xp33_ASAP7_75t_L g1619 ( 
.A1(n_1600),
.A2(n_1529),
.B(n_1528),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1573),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1588),
.Y(n_1621)
);

AOI211xp5_ASAP7_75t_L g1622 ( 
.A1(n_1569),
.A2(n_1543),
.B(n_1527),
.C(n_1415),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1583),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1591),
.A2(n_1527),
.B(n_1533),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1591),
.B(n_1537),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1626),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1623),
.B(n_1601),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1577),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1603),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1606),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1602),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1626),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1615),
.B(n_1581),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1624),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1604),
.A2(n_1611),
.B1(n_1610),
.B2(n_1619),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1585),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1613),
.B(n_1584),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1618),
.B(n_1584),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_SL g1642 ( 
.A(n_1618),
.B(n_1248),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1617),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1622),
.B(n_1577),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1592),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1637),
.A2(n_1621),
.B1(n_1620),
.B2(n_1614),
.C(n_1592),
.Y(n_1648)
);

AOI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1639),
.A2(n_1636),
.B(n_1643),
.C(n_1628),
.Y(n_1649)
);

NAND2x1_ASAP7_75t_L g1650 ( 
.A(n_1635),
.B(n_1589),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1638),
.A2(n_1598),
.B(n_1566),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1634),
.A2(n_1587),
.B1(n_1582),
.B2(n_1566),
.C(n_1565),
.Y(n_1652)
);

AND4x1_ASAP7_75t_L g1653 ( 
.A(n_1642),
.B(n_1265),
.C(n_1582),
.D(n_1587),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1632),
.A2(n_1589),
.B1(n_1565),
.B2(n_1594),
.C(n_1571),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1630),
.B(n_1571),
.Y(n_1655)
);

NOR3xp33_ASAP7_75t_L g1656 ( 
.A(n_1644),
.B(n_1594),
.C(n_1533),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_L g1657 ( 
.A1(n_1640),
.A2(n_1411),
.B(n_1537),
.C(n_1290),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1629),
.B(n_1589),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1655),
.Y(n_1659)
);

NOR3x1_ASAP7_75t_L g1660 ( 
.A(n_1651),
.B(n_1633),
.C(n_1627),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1650),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1653),
.B(n_1630),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1654),
.B(n_1627),
.Y(n_1663)
);

NAND4xp75_ASAP7_75t_L g1664 ( 
.A(n_1648),
.B(n_1645),
.C(n_1633),
.D(n_1631),
.Y(n_1664)
);

AND5x1_ASAP7_75t_L g1665 ( 
.A(n_1649),
.B(n_1646),
.C(n_1645),
.D(n_1641),
.E(n_1635),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1656),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1652),
.B(n_1647),
.Y(n_1667)
);

NOR2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1664),
.B(n_1658),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1663),
.B(n_1657),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1659),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1662),
.B(n_1589),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1667),
.B(n_1220),
.C(n_1206),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1669),
.A2(n_1661),
.B1(n_1668),
.B2(n_1671),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1670),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1672),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1669),
.B(n_1666),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1670),
.Y(n_1677)
);

NOR2x2_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1665),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1676),
.B(n_1660),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1674),
.B(n_1521),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1677),
.Y(n_1681)
);

INVx3_ASAP7_75t_SL g1682 ( 
.A(n_1678),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1673),
.B(n_1468),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1681),
.B(n_1675),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1679),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1680),
.Y(n_1686)
);

AO22x2_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1683),
.B1(n_1682),
.B2(n_1465),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1685),
.B(n_1684),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1688),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1688),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1689),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1690),
.A2(n_1684),
.B(n_1465),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1691),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1692),
.B(n_1280),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1694),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_R g1696 ( 
.A1(n_1695),
.A2(n_1692),
.B1(n_1437),
.B2(n_1434),
.C(n_1280),
.Y(n_1696)
);

AOI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1273),
.B(n_1220),
.C(n_1206),
.Y(n_1697)
);


endmodule