module fake_jpeg_27704_n_296 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx24_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_26),
.B1(n_18),
.B2(n_20),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_37),
.A2(n_28),
.B1(n_32),
.B2(n_17),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_21),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_14),
.B1(n_21),
.B2(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_58),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_66),
.Y(n_89)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

NAND5xp2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_30),
.C(n_29),
.D(n_31),
.E(n_20),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_15),
.B(n_20),
.C(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_32),
.B1(n_42),
.B2(n_39),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2x1_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_36),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_64),
.B(n_36),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_32),
.B1(n_42),
.B2(n_39),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_38),
.C(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_77),
.C(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_38),
.C(n_48),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_78),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_45),
.B1(n_50),
.B2(n_28),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_91),
.B1(n_56),
.B2(n_39),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_47),
.C(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_61),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_19),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_22),
.C(n_17),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_47),
.C(n_28),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_35),
.C(n_36),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_90),
.B1(n_70),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_42),
.B1(n_39),
.B2(n_47),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_16),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_97),
.B(n_99),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_105),
.B1(n_106),
.B2(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_63),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_107),
.B1(n_91),
.B2(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_70),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_72),
.B1(n_70),
.B2(n_65),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_53),
.B1(n_69),
.B2(n_67),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_57),
.B1(n_49),
.B2(n_59),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_71),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_23),
.B(n_22),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_117),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_75),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_36),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_133),
.B1(n_145),
.B2(n_23),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_78),
.B1(n_49),
.B2(n_94),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_128),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_140),
.B1(n_131),
.B2(n_146),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_131),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_73),
.B1(n_83),
.B2(n_93),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_73),
.B(n_22),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_152),
.B(n_119),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_141),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_95),
.B(n_75),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_138),
.B(n_142),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_49),
.B1(n_59),
.B2(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_88),
.B1(n_80),
.B2(n_79),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_88),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_36),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_49),
.B1(n_41),
.B2(n_71),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_99),
.B(n_120),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_110),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_157),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_110),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_104),
.C(n_115),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_168),
.C(n_177),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_164),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_163),
.A2(n_165),
.B(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_98),
.B(n_104),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_103),
.C(n_113),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_113),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_137),
.Y(n_186)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_124),
.B1(n_142),
.B2(n_25),
.Y(n_198)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_175),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_16),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_180),
.C(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_35),
.C(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_179),
.A2(n_182),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_16),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_24),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_25),
.B1(n_19),
.B2(n_14),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_150),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_155),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_132),
.C(n_130),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_203),
.C(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_133),
.B1(n_123),
.B2(n_135),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_209),
.B1(n_171),
.B2(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_19),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_24),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_35),
.C(n_24),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_174),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_176),
.B(n_185),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_24),
.C(n_2),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_170),
.B1(n_158),
.B2(n_182),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_167),
.B(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_219),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_216),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_191),
.B(n_194),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_222),
.B(n_198),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_181),
.B1(n_184),
.B2(n_168),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_225),
.B1(n_192),
.B2(n_190),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_195),
.B(n_206),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_1),
.C(n_3),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_220),
.C(n_215),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_4),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_210),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_206),
.B(n_202),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_231),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_189),
.C(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_243),
.C(n_210),
.Y(n_246)
);

BUFx12f_ASAP7_75t_SL g236 ( 
.A(n_223),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_225),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_204),
.C(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_244),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_200),
.C(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.C(n_252),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_200),
.C(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_212),
.C(n_226),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_219),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_232),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_233),
.B(n_239),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_4),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_268),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_240),
.B1(n_214),
.B2(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_243),
.C(n_245),
.Y(n_264)
);

OAI321xp33_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_231),
.A3(n_203),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_251),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_7),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_256),
.C(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_4),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_278),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_258),
.B1(n_5),
.B2(n_6),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_5),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_5),
.B(n_6),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_7),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_9),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_272),
.C(n_274),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_283),
.B(n_11),
.C(n_12),
.D(n_10),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_291),
.A2(n_288),
.B(n_287),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_292),
.B(n_11),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_10),
.B(n_12),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_295),
.A2(n_10),
.B(n_12),
.Y(n_296)
);


endmodule