module fake_jpeg_2392_n_223 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_223);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_SL g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_35),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_85),
.B1(n_57),
.B2(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_61),
.B1(n_84),
.B2(n_89),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_72),
.B1(n_60),
.B2(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_99),
.B1(n_80),
.B2(n_69),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_73),
.B1(n_63),
.B2(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_63),
.B1(n_73),
.B2(n_62),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_79),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_67),
.B1(n_65),
.B2(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_74),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_121),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_56),
.B1(n_61),
.B2(n_76),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_96),
.B1(n_89),
.B2(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_67),
.B1(n_56),
.B2(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_131),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_101),
.B1(n_98),
.B2(n_96),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_130),
.B1(n_133),
.B2(n_142),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_58),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_69),
.B1(n_76),
.B2(n_71),
.Y(n_133)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_96),
.C(n_118),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_20),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_21),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_24),
.B(n_51),
.C(n_49),
.D(n_48),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_68),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_152),
.Y(n_185)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_159),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_166),
.B(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_2),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_54),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_132),
.A3(n_144),
.B1(n_138),
.B2(n_10),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_3),
.B(n_6),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_7),
.B(n_8),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_6),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_7),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_178),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_171),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_26),
.B(n_41),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_186),
.B(n_36),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_28),
.B1(n_40),
.B2(n_39),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_47),
.B(n_38),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_151),
.C(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_197),
.C(n_161),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_29),
.B(n_13),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_162),
.Y(n_190)
);

AOI321xp33_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_173),
.A3(n_175),
.B1(n_179),
.B2(n_176),
.C(n_187),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_176),
.B1(n_182),
.B2(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_177),
.B(n_164),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_159),
.C(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_165),
.B1(n_171),
.B2(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_184),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_203),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_154),
.C(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_196),
.B(n_189),
.C(n_15),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_211),
.B(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_210),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_207),
.C(n_208),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_189),
.B(n_209),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_215),
.CI(n_208),
.CON(n_218),
.SN(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_12),
.B(n_14),
.Y(n_219)
);

OAI322xp33_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_16),
.A3(n_18),
.B1(n_19),
.B2(n_218),
.C1(n_188),
.C2(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_16),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_222),
.Y(n_223)
);


endmodule