module fake_netlist_6_652_n_4173 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_70, n_18, n_10, n_21, n_24, n_71, n_74, n_37, n_6, n_15, n_33, n_54, n_67, n_27, n_3, n_14, n_38, n_72, n_0, n_61, n_39, n_63, n_60, n_59, n_73, n_32, n_4, n_66, n_36, n_22, n_26, n_68, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_69, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_65, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_4173);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_70;
input n_18;
input n_10;
input n_21;
input n_24;
input n_71;
input n_74;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_67;
input n_27;
input n_3;
input n_14;
input n_38;
input n_72;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_73;
input n_32;
input n_4;
input n_66;
input n_36;
input n_22;
input n_26;
input n_68;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_69;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_65;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_4173;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_223;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_212;
wire n_3783;
wire n_700;
wire n_3773;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_3844;
wire n_168;
wire n_1237;
wire n_1061;
wire n_2534;
wire n_2353;
wire n_3089;
wire n_3301;
wire n_4099;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_77;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_3253;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_3222;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_350;
wire n_78;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_442;
wire n_480;
wire n_142;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_3706;
wire n_4050;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_3668;
wire n_1247;
wire n_2336;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_424;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_369;
wire n_287;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_3340;
wire n_461;
wire n_873;
wire n_383;
wire n_141;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_200;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_229;
wire n_3282;
wire n_2513;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_2645;
wire n_3757;
wire n_3904;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_3106;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_3031;
wire n_2019;
wire n_4029;
wire n_836;
wire n_3345;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_658;
wire n_616;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2739;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_3023;
wire n_3890;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_405;
wire n_213;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_155;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_112;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_126;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_224;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_407;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_163;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_4102;
wire n_757;
wire n_594;
wire n_1641;
wire n_3871;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2113;
wire n_2907;
wire n_577;
wire n_3438;
wire n_166;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_323;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_92;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_331;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4009;
wire n_2633;
wire n_483;
wire n_102;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_261;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_121;
wire n_3484;
wire n_433;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_219;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_264;
wire n_263;
wire n_3900;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_329;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_408;
wire n_932;
wire n_2998;
wire n_2831;
wire n_3446;
wire n_4158;
wire n_3317;
wire n_237;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_117;
wire n_175;
wire n_322;
wire n_993;
wire n_2692;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_3914;
wire n_2228;
wire n_3397;
wire n_134;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_136;
wire n_966;
wire n_3888;
wire n_3168;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_241;
wire n_3966;
wire n_2866;
wire n_1107;
wire n_2068;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_318;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_88;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_199;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_3581;
wire n_2428;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_3933;
wire n_702;
wire n_347;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_2510;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_195;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_286;
wire n_254;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_728;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_267;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2980;
wire n_2096;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_3510;
wire n_437;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_3289;
wire n_2824;
wire n_2733;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_388;
wire n_190;
wire n_2812;
wire n_484;
wire n_2644;
wire n_3326;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_170;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2921;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_3519;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_283;
wire n_2075;
wire n_4045;
wire n_2972;
wire n_2194;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_91;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_362;
wire n_148;
wire n_2279;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_304;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_125;
wire n_1634;
wire n_3252;
wire n_2078;
wire n_2932;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3431;
wire n_3337;
wire n_3450;
wire n_342;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_131;
wire n_1523;
wire n_2558;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_2750;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_382;
wire n_673;
wire n_2705;
wire n_2230;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_289;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_320;
wire n_108;
wire n_639;
wire n_963;
wire n_794;
wire n_2767;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_353;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_86;
wire n_3179;
wire n_104;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_305;
wire n_2554;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_413;
wire n_3171;
wire n_791;
wire n_1913;
wire n_3608;
wire n_510;
wire n_837;
wire n_2097;
wire n_79;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_147;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_153;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_3082;
wire n_3611;
wire n_2239;
wire n_1432;
wire n_156;
wire n_145;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2717;
wire n_1723;
wire n_2191;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_189;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_294;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2307;
wire n_2069;
wire n_3704;
wire n_2362;
wire n_425;
wire n_684;
wire n_2667;
wire n_2698;
wire n_2539;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_3020;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_290;
wire n_118;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_107;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_417;
wire n_2857;
wire n_446;
wire n_3693;
wire n_3788;
wire n_89;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2959;
wire n_2494;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_293;
wire n_4085;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_154;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_98;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_184;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_216;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_3056;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_3103;
wire n_3032;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_3393;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_312;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_100;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_150;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2788;
wire n_2218;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_124;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_211;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_319;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_3964;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_311;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_123;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_162;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_128;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_3481;
wire n_1092;
wire n_2329;
wire n_2237;
wire n_3026;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_444;
wire n_3033;
wire n_3724;
wire n_146;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_303;
wire n_511;
wire n_2990;
wire n_3847;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_113;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_4020;
wire n_266;
wire n_296;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_3407;
wire n_217;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_3425;
wire n_215;
wire n_2384;
wire n_3894;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_426;
wire n_317;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_90;
wire n_3986;
wire n_2601;
wire n_3454;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2502;
wire n_2131;
wire n_488;
wire n_3646;
wire n_2801;
wire n_2226;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_99;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_401;
wire n_4034;
wire n_324;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_335;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_120;
wire n_2732;
wire n_301;
wire n_2928;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_427;
wire n_2572;
wire n_2720;
wire n_1520;
wire n_496;
wire n_3126;
wire n_2204;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_3663;
wire n_2315;
wire n_4132;
wire n_351;
wire n_2955;
wire n_2995;
wire n_259;
wire n_1731;
wire n_177;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3360;
wire n_1437;
wire n_3051;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_379;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_410;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_171;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_169;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_341;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2875;
wire n_1103;
wire n_2448;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_144;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_106;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_186;
wire n_2984;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_392;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3276;
wire n_3113;
wire n_3250;
wire n_1934;
wire n_3194;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_349;
wire n_3448;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_140;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_421;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_280;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_198;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_179;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_3141;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_3839;
wire n_2823;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_466;
wire n_3041;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_235;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_101;
wire n_167;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_127;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_133;
wire n_1320;
wire n_2716;
wire n_96;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_137;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_397;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_122;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_218;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_172;
wire n_3536;
wire n_4109;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_3424;
wire n_2894;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_239;
wire n_2037;
wire n_97;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_220;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_80;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_402;
wire n_1870;
wire n_352;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_450;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2699;
wire n_3029;
wire n_2200;
wire n_2272;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_3329;
wire n_2704;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_260;
wire n_2670;
wire n_313;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_356;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_83;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_411;
wire n_2518;
wire n_2458;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_105;
wire n_2782;
wire n_3977;
wire n_227;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_1489;
wire n_164;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_4040;
wire n_804;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2562;
wire n_2141;
wire n_244;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_76;
wire n_2734;
wire n_548;
wire n_1782;
wire n_94;
wire n_282;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_345;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_139;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_273;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_3007;
wire n_2809;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_159;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_157;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_3517;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_346;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_138;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_4052;
wire n_2680;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_431;
wire n_3379;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_285;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_85;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_75;
wire n_743;
wire n_766;
wire n_3124;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_1804;
wire n_2923;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_251;
wire n_2508;
wire n_1019;
wire n_636;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_151;
wire n_110;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_262;
wire n_3602;
wire n_187;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_3391;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_332;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_194;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_278;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_384;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_310;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_84;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_143;
wire n_1536;
wire n_3846;
wire n_180;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_3874;
wire n_1379;
wire n_2814;
wire n_2528;
wire n_214;
wire n_246;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_181;
wire n_1810;
wire n_182;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_176;
wire n_114;
wire n_300;
wire n_222;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_372;
wire n_2076;
wire n_3583;
wire n_111;
wire n_2883;
wire n_2736;
wire n_314;
wire n_3860;
wire n_1408;
wire n_378;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_377;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_3774;
wire n_2182;
wire n_338;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_119;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_3739;
wire n_3898;
wire n_2485;
wire n_2284;
wire n_3520;
wire n_191;
wire n_2566;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_344;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_174;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_129;
wire n_3336;
wire n_647;
wire n_4160;
wire n_197;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_109;
wire n_445;
wire n_3553;
wire n_1561;
wire n_3114;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_82;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_270;
wire n_2265;
wire n_2615;
wire n_414;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_93;
wire n_839;
wire n_2437;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_3362;
wire n_3745;
wire n_2242;
wire n_4059;
wire n_1509;
wire n_103;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_185;
wire n_2222;
wire n_712;
wire n_3256;
wire n_348;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_376;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2466;
wire n_3982;
wire n_390;
wire n_2111;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_334;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_232;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_298;
wire n_1582;
wire n_492;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_265;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2950;
wire n_2483;
wire n_228;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_3123;
wire n_393;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_132;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_130;
wire n_3285;
wire n_519;
wire n_2523;
wire n_307;
wire n_469;
wire n_1218;
wire n_3769;
wire n_500;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_291;
wire n_4089;
wire n_1144;
wire n_3669;
wire n_3863;
wire n_2071;
wire n_357;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_436;
wire n_4075;
wire n_116;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_240;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_95;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_253;
wire n_3976;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_3876;
wire n_249;
wire n_201;
wire n_3198;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_115;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_467;
wire n_3187;
wire n_2540;
wire n_269;
wire n_359;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2461;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_158;
wire n_2107;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_3110;
wire n_87;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_207;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_205;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_412;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_640;
wire n_1322;
wire n_81;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_135;
wire n_3079;
wire n_165;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_364;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_361;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_192;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_27),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_15),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_11),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_7),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_40),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_15),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_13),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_6),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_14),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_12),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_32),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_48),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_1),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_43),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_24),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_32),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_4),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_31),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_5),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_23),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_21),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_20),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_30),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_23),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_13),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_51),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_49),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_4),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_3),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_9),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_9),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_10),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_45),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_17),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_0),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_38),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_21),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVxp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

BUFx2_ASAP7_75t_SL g164 ( 
.A(n_111),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_113),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_77),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_82),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_162),
.B(n_157),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_142),
.B1(n_83),
.B2(n_111),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_142),
.B1(n_83),
.B2(n_144),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

AOI22x1_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_86),
.B1(n_147),
.B2(n_144),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_147),
.B1(n_129),
.B2(n_86),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_117),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_150),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_82),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_89),
.B1(n_90),
.B2(n_129),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_202),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_163),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_152),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_166),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_163),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_117),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_99),
.B1(n_91),
.B2(n_90),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_169),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_81),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

AND3x1_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_98),
.C(n_91),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_177),
.B(n_169),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_175),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_187),
.A2(n_114),
.B(n_125),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_177),
.B(n_109),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_175),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_203),
.B(n_152),
.Y(n_266)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_201),
.B(n_109),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_182),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_114),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_191),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_195),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_201),
.B(n_119),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_182),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_119),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_191),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_182),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_191),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_192),
.B(n_120),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_182),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_205),
.A2(n_103),
.B1(n_99),
.B2(n_98),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_191),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_182),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_182),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_191),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_188),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_194),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_188),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_186),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_194),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_188),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_188),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_212),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_266),
.C(n_167),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_212),
.B(n_177),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_212),
.B(n_177),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g310 ( 
.A(n_210),
.B(n_213),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_231),
.B(n_164),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_212),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_224),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_241),
.A2(n_202),
.B1(n_196),
.B2(n_176),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_176),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_238),
.A2(n_201),
.B1(n_192),
.B2(n_186),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_211),
.B(n_176),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_233),
.B(n_252),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_192),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_232),
.B(n_196),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_233),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_192),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_232),
.B(n_196),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_252),
.B(n_201),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_211),
.B(n_202),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_224),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_211),
.B(n_166),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_238),
.A2(n_201),
.B1(n_192),
.B2(n_186),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_247),
.B(n_206),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_224),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_248),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_252),
.B(n_200),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_225),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_167),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_259),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_225),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_239),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_259),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_239),
.B(n_200),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g345 ( 
.A(n_271),
.B(n_186),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_239),
.B(n_200),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_201),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_250),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_243),
.A2(n_201),
.B1(n_208),
.B2(n_209),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_259),
.B(n_168),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_274),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_274),
.B(n_168),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_281),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_248),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_179),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_L g357 ( 
.A(n_210),
.B(n_116),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_250),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_248),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_250),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_248),
.B(n_153),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_248),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_210),
.B(n_120),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_256),
.B(n_165),
.Y(n_364)
);

AO22x2_ASAP7_75t_L g365 ( 
.A1(n_247),
.A2(n_183),
.B1(n_179),
.B2(n_181),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_241),
.B(n_116),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_256),
.B(n_165),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_256),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_257),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_257),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_257),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_217),
.Y(n_372)
);

BUFx8_ASAP7_75t_SL g373 ( 
.A(n_276),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_263),
.B(n_200),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_241),
.B(n_75),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_263),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_263),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_243),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_295),
.Y(n_379)
);

NOR2x1p5_ASAP7_75t_L g380 ( 
.A(n_278),
.B(n_126),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_264),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_217),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_264),
.B(n_179),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_217),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_264),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_276),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_265),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_217),
.Y(n_388)
);

AO22x2_ASAP7_75t_L g389 ( 
.A1(n_247),
.A2(n_183),
.B1(n_179),
.B2(n_181),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_217),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_265),
.B(n_187),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_265),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_272),
.B(n_183),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_272),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_272),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_275),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_267),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_275),
.A2(n_209),
.B1(n_208),
.B2(n_200),
.Y(n_398)
);

AND3x4_ASAP7_75t_L g399 ( 
.A(n_276),
.B(n_183),
.C(n_181),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_287),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_275),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_255),
.B(n_200),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_228),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_217),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_287),
.B(n_187),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_287),
.B(n_206),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_217),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_276),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_214),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_255),
.B(n_200),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_214),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_228),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_255),
.B(n_200),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_276),
.B(n_78),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_276),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_214),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_276),
.B(n_79),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_228),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_278),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_255),
.B(n_181),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_217),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_213),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_278),
.B(n_80),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_217),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_217),
.Y(n_425)
);

BUFx6f_ASAP7_75t_SL g426 ( 
.A(n_267),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_219),
.B(n_84),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_219),
.B(n_200),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_267),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_242),
.B(n_85),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_258),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_282),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_213),
.B(n_200),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_282),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_220),
.B(n_208),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_220),
.A2(n_125),
.B1(n_138),
.B2(n_146),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_242),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_267),
.A2(n_104),
.B1(n_97),
.B2(n_88),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_226),
.Y(n_439)
);

OR2x6_ASAP7_75t_L g440 ( 
.A(n_220),
.B(n_138),
.Y(n_440)
);

INVx8_ASAP7_75t_L g441 ( 
.A(n_267),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_221),
.B(n_89),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_214),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_221),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_221),
.B(n_87),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_222),
.B(n_126),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_282),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_222),
.A2(n_209),
.B1(n_208),
.B2(n_207),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_222),
.B(n_92),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_267),
.A2(n_209),
.B1(n_208),
.B2(n_207),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_226),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_258),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_289),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_223),
.B(n_93),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_215),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_223),
.B(n_121),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_226),
.Y(n_457)
);

NOR2x1p5_ASAP7_75t_L g458 ( 
.A(n_270),
.B(n_126),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_289),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_267),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_226),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_289),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_223),
.B(n_187),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_292),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_292),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_270),
.B(n_95),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_267),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_258),
.B(n_204),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_226),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_226),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_285),
.A2(n_136),
.B1(n_209),
.B2(n_208),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_292),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_L g473 ( 
.A(n_267),
.B(n_226),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_297),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_267),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_258),
.B(n_204),
.Y(n_476)
);

INVx4_ASAP7_75t_SL g477 ( 
.A(n_267),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_258),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_297),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_317),
.B(n_297),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_361),
.B(n_143),
.C(n_102),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_432),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_320),
.B(n_206),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_419),
.B(n_300),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_351),
.B(n_285),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_313),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_351),
.B(n_216),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_328),
.B(n_96),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_338),
.B(n_100),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_309),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_391),
.B(n_300),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_353),
.B(n_101),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_391),
.B(n_300),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_L g495 ( 
.A(n_315),
.B(n_145),
.C(n_107),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_305),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_405),
.B(n_301),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_308),
.B(n_216),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_313),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_405),
.B(n_301),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_308),
.B(n_216),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_437),
.B(n_301),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_329),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_329),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_333),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_330),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_333),
.Y(n_507)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_441),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_441),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_336),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_463),
.B(n_215),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_463),
.B(n_215),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_403),
.B(n_215),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_336),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_403),
.B(n_218),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_412),
.B(n_218),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_393),
.A2(n_267),
.B1(n_258),
.B2(n_246),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_412),
.B(n_218),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_418),
.B(n_339),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_418),
.B(n_218),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_364),
.A2(n_267),
.B1(n_258),
.B2(n_227),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_309),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_342),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g527 ( 
.A(n_330),
.B(n_52),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_305),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_308),
.A2(n_299),
.B1(n_298),
.B2(n_227),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_339),
.B(n_227),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_386),
.B(n_216),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_312),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_343),
.B(n_227),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_343),
.B(n_236),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_352),
.B(n_108),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_310),
.B(n_226),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_352),
.B(n_110),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_311),
.B(n_236),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_466),
.B(n_236),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_312),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_399),
.A2(n_106),
.B1(n_103),
.B2(n_123),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_386),
.B(n_216),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_427),
.B(n_236),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_342),
.B(n_237),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_354),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_408),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_348),
.B(n_237),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_348),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_360),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_382),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_383),
.A2(n_299),
.B1(n_298),
.B2(n_237),
.Y(n_552)
);

O2A1O1Ixp5_ASAP7_75t_L g553 ( 
.A1(n_456),
.A2(n_299),
.B(n_298),
.C(n_237),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_379),
.B(n_112),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_360),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_314),
.B(n_244),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_306),
.B(n_216),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_321),
.B(n_234),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_368),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_368),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_369),
.B(n_244),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_369),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_370),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_370),
.B(n_244),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_434),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_367),
.B(n_115),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_314),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_381),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_400),
.B(n_122),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_381),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_324),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_420),
.A2(n_299),
.B(n_298),
.C(n_294),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_337),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_385),
.B(n_244),
.Y(n_574)
);

AOI22x1_ASAP7_75t_L g575 ( 
.A1(n_458),
.A2(n_380),
.B1(n_341),
.B2(n_358),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_307),
.B(n_234),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_385),
.B(n_245),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_324),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_307),
.B(n_234),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_387),
.B(n_245),
.Y(n_580)
);

BUFx5_ASAP7_75t_L g581 ( 
.A(n_310),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_387),
.B(n_245),
.Y(n_582)
);

O2A1O1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_366),
.A2(n_357),
.B(n_436),
.C(n_335),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_447),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_395),
.B(n_245),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_L g586 ( 
.A(n_445),
.B(n_53),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_447),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_378),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_372),
.A2(n_277),
.B(n_294),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_395),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_382),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_310),
.B(n_226),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_453),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_340),
.A2(n_249),
.B1(n_253),
.B2(n_234),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_453),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_307),
.B(n_234),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_307),
.B(n_362),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_396),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_459),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_462),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_462),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_310),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_378),
.B(n_124),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_327),
.A2(n_261),
.B(n_294),
.C(n_290),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_396),
.B(n_246),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_337),
.B(n_127),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_323),
.B(n_141),
.C(n_132),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_349),
.B(n_130),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_327),
.B(n_246),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_307),
.B(n_234),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_349),
.B(n_131),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_408),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_362),
.B(n_249),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_318),
.B(n_249),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_340),
.B(n_246),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_341),
.B(n_251),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_406),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_464),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_464),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_465),
.Y(n_621)
);

BUFx5_ASAP7_75t_L g622 ( 
.A(n_310),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_415),
.A2(n_277),
.B1(n_294),
.B2(n_254),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_358),
.B(n_251),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_362),
.B(n_249),
.Y(n_625)
);

NAND3x1_ASAP7_75t_L g626 ( 
.A(n_399),
.B(n_123),
.C(n_106),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_356),
.B(n_133),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_458),
.B(n_380),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_465),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_302),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_362),
.B(n_249),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_472),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_302),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_371),
.B(n_251),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_371),
.B(n_251),
.Y(n_635)
);

INVx8_ASAP7_75t_L g636 ( 
.A(n_441),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_362),
.B(n_249),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_303),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_472),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_357),
.A2(n_260),
.B(n_290),
.C(n_254),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_303),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_376),
.A2(n_253),
.B1(n_288),
.B2(n_261),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_347),
.A2(n_277),
.B1(n_254),
.B2(n_260),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_356),
.B(n_134),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_326),
.B(n_135),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_376),
.B(n_254),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_SL g647 ( 
.A(n_426),
.B(n_226),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_345),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_304),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_377),
.B(n_260),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_415),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_365),
.A2(n_113),
.B1(n_140),
.B2(n_149),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_347),
.A2(n_261),
.B(n_290),
.C(n_262),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_440),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_345),
.B(n_137),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_382),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_304),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_382),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_316),
.B(n_253),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_377),
.B(n_262),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_440),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_440),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_316),
.B(n_253),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_316),
.B(n_253),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_440),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_409),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_334),
.B(n_253),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_334),
.B(n_288),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_474),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_392),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_334),
.B(n_288),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_409),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_322),
.A2(n_262),
.B(n_290),
.C(n_268),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_474),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_318),
.A2(n_269),
.B1(n_268),
.B2(n_277),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_382),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_355),
.B(n_288),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_411),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_411),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_355),
.B(n_288),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_406),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_416),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_319),
.B(n_268),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_392),
.B(n_268),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_331),
.B(n_269),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_394),
.B(n_269),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_394),
.B(n_269),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_482),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_491),
.B(n_449),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_573),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_547),
.B(n_359),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_487),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_482),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_537),
.A2(n_384),
.B(n_372),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_487),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_566),
.A2(n_399),
.B1(n_345),
.B2(n_375),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_491),
.B(n_454),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_490),
.B(n_345),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_524),
.B(n_401),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_588),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_583),
.A2(n_478),
.B(n_452),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_524),
.B(n_401),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_573),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_509),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_627),
.B(n_365),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_547),
.B(n_359),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_537),
.A2(n_388),
.B(n_384),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_551),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_551),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_499),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_603),
.B(n_581),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_588),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_483),
.B(n_332),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_603),
.B(n_421),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_489),
.B(n_325),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_551),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_499),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_521),
.B(n_310),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_613),
.B(n_429),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_481),
.A2(n_423),
.B1(n_430),
.B2(n_417),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_531),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_506),
.B(n_332),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_613),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_541),
.B(n_571),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_541),
.B(n_310),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_493),
.A2(n_414),
.B1(n_389),
.B2(n_365),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_485),
.B(n_460),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_571),
.B(n_428),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_509),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_628),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_503),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_681),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_503),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_508),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_591),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_504),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_648),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_508),
.B(n_446),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_546),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_485),
.B(n_429),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_604),
.B(n_373),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_504),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_516),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_535),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_516),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_495),
.A2(n_365),
.B1(n_389),
.B2(n_442),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_591),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_603),
.B(n_421),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_628),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_525),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_618),
.B(n_460),
.Y(n_753)
);

CKINVDCx11_ASAP7_75t_R g754 ( 
.A(n_618),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_508),
.B(n_446),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_644),
.B(n_389),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_538),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_505),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_505),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_683),
.B(n_442),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_683),
.B(n_442),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_685),
.B(n_442),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_525),
.Y(n_763)
);

BUFx6f_ASAP7_75t_SL g764 ( 
.A(n_654),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_536),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_592),
.A2(n_384),
.B(n_372),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_685),
.B(n_442),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_507),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_496),
.B(n_442),
.Y(n_769)
);

AND2x2_ASAP7_75t_SL g770 ( 
.A(n_655),
.B(n_473),
.Y(n_770)
);

AND2x6_ASAP7_75t_SL g771 ( 
.A(n_569),
.B(n_446),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_SL g772 ( 
.A(n_485),
.B(n_426),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_603),
.B(n_421),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_591),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_581),
.B(n_422),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_654),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_536),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_565),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_554),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_645),
.A2(n_389),
.B1(n_475),
.B2(n_438),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_528),
.B(n_442),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_532),
.B(n_431),
.Y(n_782)
);

NOR2x1p5_ASAP7_75t_L g783 ( 
.A(n_567),
.B(n_139),
.Y(n_783)
);

INVx5_ASAP7_75t_L g784 ( 
.A(n_591),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_578),
.B(n_344),
.Y(n_785)
);

CKINVDCx11_ASAP7_75t_R g786 ( 
.A(n_508),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_565),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_603),
.B(n_421),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_584),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_591),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_607),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_531),
.B(n_543),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_497),
.B(n_346),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_584),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_626),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_486),
.A2(n_475),
.B1(n_363),
.B2(n_426),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_500),
.B(n_374),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_507),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_484),
.B(n_468),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_581),
.B(n_421),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_531),
.B(n_477),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_510),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_510),
.B(n_636),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_609),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_581),
.B(n_425),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_608),
.A2(n_363),
.B1(n_446),
.B2(n_473),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_581),
.B(n_622),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_511),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_610),
.B(n_468),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_587),
.Y(n_810)
);

NOR2x2_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_416),
.Y(n_811)
);

NOR2x2_ASAP7_75t_L g812 ( 
.A(n_652),
.B(n_443),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_543),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_542),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_612),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_527),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_587),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_510),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_593),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_592),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_488),
.B(n_402),
.Y(n_821)
);

INVx5_ASAP7_75t_L g822 ( 
.A(n_510),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_615),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_593),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_511),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_610),
.B(n_476),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_595),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_498),
.B(n_501),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_R g829 ( 
.A(n_647),
.B(n_363),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_575),
.A2(n_363),
.B1(n_350),
.B2(n_476),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_670),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_661),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_595),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_661),
.B(n_410),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_543),
.B(n_477),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_662),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_SL g837 ( 
.A(n_519),
.B(n_148),
.C(n_450),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_662),
.B(n_413),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_665),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_480),
.B(n_492),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_670),
.A2(n_444),
.B1(n_422),
.B2(n_455),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_665),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_575),
.A2(n_363),
.B1(n_467),
.B2(n_397),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_581),
.B(n_425),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_515),
.B(n_433),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_615),
.B(n_477),
.Y(n_846)
);

NOR2x2_ASAP7_75t_L g847 ( 
.A(n_542),
.B(n_443),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_596),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_636),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_596),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_542),
.B(n_113),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_542),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_515),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_494),
.B(n_398),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_586),
.A2(n_444),
.B(n_450),
.C(n_435),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_581),
.B(n_425),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_556),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_523),
.A2(n_363),
.B(n_448),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_615),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_502),
.B(n_363),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_630),
.B(n_390),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_622),
.B(n_425),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_L g863 ( 
.A(n_622),
.B(n_425),
.Y(n_863)
);

AND2x6_ASAP7_75t_L g864 ( 
.A(n_630),
.B(n_439),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_633),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_636),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_526),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_556),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_526),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_557),
.A2(n_471),
.B(n_286),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_633),
.B(n_390),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_638),
.A2(n_451),
.B1(n_424),
.B2(n_469),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_636),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_638),
.B(n_390),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_600),
.Y(n_875)
);

NAND2x1p5_ASAP7_75t_L g876 ( 
.A(n_598),
.B(n_397),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_641),
.A2(n_657),
.B1(n_649),
.B2(n_669),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_622),
.B(n_439),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_641),
.B(n_477),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_649),
.B(n_439),
.Y(n_880)
);

BUFx10_ASAP7_75t_L g881 ( 
.A(n_600),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_601),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_549),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_601),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_657),
.B(n_404),
.Y(n_885)
);

BUFx12f_ASAP7_75t_SL g886 ( 
.A(n_647),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_549),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_602),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_512),
.B(n_404),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_550),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_550),
.B(n_286),
.Y(n_891)
);

BUFx12f_ASAP7_75t_L g892 ( 
.A(n_576),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_602),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_622),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_622),
.B(n_439),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_558),
.A2(n_397),
.B1(n_467),
.B2(n_439),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_513),
.B(n_404),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_555),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_555),
.B(n_407),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_559),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_559),
.B(n_407),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_619),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_560),
.Y(n_903)
);

AND2x6_ASAP7_75t_SL g904 ( 
.A(n_530),
.B(n_190),
.Y(n_904)
);

BUFx4f_ASAP7_75t_L g905 ( 
.A(n_619),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_560),
.B(n_286),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_562),
.B(n_563),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_SL g908 ( 
.A(n_540),
.B(n_190),
.C(n_197),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_562),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_563),
.B(n_407),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_620),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_620),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_568),
.B(n_470),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_621),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_621),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_568),
.B(n_286),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_570),
.B(n_470),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_653),
.A2(n_190),
.B(n_197),
.C(n_470),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_622),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_629),
.A2(n_397),
.B1(n_467),
.B2(n_457),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_629),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_570),
.B(n_457),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_590),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_590),
.B(n_457),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_599),
.B(n_457),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_599),
.B(n_457),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_632),
.Y(n_927)
);

INVx5_ASAP7_75t_L g928 ( 
.A(n_666),
.Y(n_928)
);

OR2x6_ASAP7_75t_L g929 ( 
.A(n_632),
.B(n_388),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_514),
.B(n_388),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_639),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_639),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_674),
.A2(n_397),
.B1(n_467),
.B2(n_461),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_674),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_666),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_672),
.B(n_208),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_679),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_672),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_678),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_517),
.B(n_424),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_SL g941 ( 
.A1(n_656),
.A2(n_397),
.B1(n_467),
.B2(n_5),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_677),
.B(n_467),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_716),
.B(n_518),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_815),
.B(n_520),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_710),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_701),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_779),
.B(n_522),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_840),
.B(n_544),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_699),
.B(n_714),
.C(n_746),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_857),
.B(n_539),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_791),
.B(n_533),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_757),
.B(n_534),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_804),
.B(n_679),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_804),
.B(n_678),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_706),
.B(n_682),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_693),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_710),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_756),
.B(n_682),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_697),
.A2(n_680),
.B1(n_663),
.B2(n_664),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_691),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_688),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_693),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_792),
.B(n_658),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_694),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_868),
.B(n_923),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_710),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_705),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_905),
.A2(n_553),
.B(n_572),
.C(n_676),
.Y(n_968)
);

AOI22x1_ASAP7_75t_L g969 ( 
.A1(n_820),
.A2(n_589),
.B1(n_451),
.B2(n_469),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_923),
.B(n_552),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_905),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_696),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_846),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_792),
.B(n_529),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_704),
.B(n_424),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_704),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_731),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_696),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_792),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_740),
.B(n_640),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_931),
.B(n_545),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_741),
.B(n_579),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_711),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_711),
.Y(n_984)
);

INVxp67_ASAP7_75t_SL g985 ( 
.A(n_863),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_865),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_739),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_739),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_690),
.B(n_548),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_745),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_747),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_770),
.B(n_597),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_723),
.B(n_611),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_728),
.A2(n_770),
.B1(n_795),
.B2(n_748),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_718),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_734),
.B(n_614),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_698),
.B(n_561),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_724),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_937),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_937),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_724),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_718),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_710),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_733),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_823),
.B(n_625),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_752),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_793),
.B(n_564),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_763),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_701),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_753),
.B(n_451),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_797),
.B(n_574),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_823),
.B(n_631),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_765),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_777),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_846),
.Y(n_1015)
);

AOI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_780),
.A2(n_673),
.B(n_659),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_720),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_733),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_751),
.Y(n_1019)
);

AND2x2_ASAP7_75t_SL g1020 ( 
.A(n_814),
.B(n_687),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_778),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_787),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_823),
.B(n_637),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_789),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_710),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_749),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_749),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_760),
.B(n_686),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_SL g1029 ( 
.A(n_806),
.B(n_623),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_859),
.B(n_643),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_863),
.A2(n_461),
.B(n_469),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_846),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_720),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_794),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_720),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_713),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_SL g1037 ( 
.A(n_743),
.B(n_713),
.Y(n_1037)
);

CKINVDCx11_ASAP7_75t_R g1038 ( 
.A(n_754),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_810),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_749),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_735),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_817),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_801),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_819),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_799),
.B(n_577),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_824),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_735),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_813),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_SL g1050 ( 
.A1(n_941),
.A2(n_684),
.B1(n_660),
.B2(n_650),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_827),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_754),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_749),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_833),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_859),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_738),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_801),
.B(n_605),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_749),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_785),
.B(n_580),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_738),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_744),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_774),
.Y(n_1062)
);

OR2x4_ASAP7_75t_L g1063 ( 
.A(n_873),
.B(n_616),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_809),
.B(n_826),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_744),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_852),
.A2(n_671),
.B1(n_668),
.B2(n_667),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_801),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_835),
.B(n_651),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_730),
.B(n_582),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_734),
.A2(n_675),
.B1(n_646),
.B2(n_617),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_732),
.B(n_585),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_758),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_758),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_864),
.Y(n_1074)
);

AO22x1_ASAP7_75t_L g1075 ( 
.A1(n_851),
.A2(n_635),
.B1(n_634),
.B2(n_624),
.Y(n_1075)
);

AOI22x1_ASAP7_75t_L g1076 ( 
.A1(n_858),
.A2(n_461),
.B1(n_190),
.B2(n_197),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_836),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_774),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_835),
.B(n_606),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_813),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_835),
.B(n_60),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_692),
.B(n_707),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_839),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_813),
.B(n_63),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_813),
.B(n_722),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_722),
.B(n_288),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_692),
.B(n_642),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_786),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_759),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_692),
.B(n_594),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_707),
.B(n_742),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_848),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_786),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_740),
.B(n_197),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_707),
.B(n_207),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_740),
.B(n_197),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_774),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_761),
.B(n_190),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_837),
.A2(n_204),
.B1(n_208),
.B2(n_209),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_SL g1100 ( 
.A1(n_721),
.A2(n_0),
.B1(n_2),
.B2(n_10),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_850),
.B(n_209),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_SL g1102 ( 
.A1(n_842),
.A2(n_2),
.B1(n_11),
.B2(n_12),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_875),
.B(n_209),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_811),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_882),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_811),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_894),
.A2(n_296),
.B1(n_293),
.B2(n_291),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_884),
.B(n_209),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_888),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_759),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_893),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_902),
.B(n_209),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_894),
.B(n_235),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_911),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_776),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_912),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_768),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_776),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_822),
.B(n_296),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_914),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_915),
.B(n_208),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_812),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_879),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_768),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_774),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_822),
.B(n_774),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_921),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_932),
.B(n_208),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_879),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_934),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_816),
.B(n_14),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_783),
.A2(n_204),
.B1(n_207),
.B2(n_198),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_700),
.B(n_207),
.Y(n_1133)
);

AND3x1_ASAP7_75t_SL g1134 ( 
.A(n_812),
.B(n_16),
.C(n_17),
.Y(n_1134)
);

BUFx8_ASAP7_75t_L g1135 ( 
.A(n_764),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_695),
.A2(n_193),
.B(n_199),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_771),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_798),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_927),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_725),
.B(n_16),
.Y(n_1140)
);

AO22x1_ASAP7_75t_L g1141 ( 
.A1(n_831),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_784),
.Y(n_1142)
);

INVxp33_ASAP7_75t_L g1143 ( 
.A(n_834),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_927),
.Y(n_1144)
);

CKINVDCx14_ASAP7_75t_R g1145 ( 
.A(n_849),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_879),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_703),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_907),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_762),
.A2(n_204),
.B1(n_207),
.B2(n_198),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_798),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_742),
.B(n_207),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_808),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_808),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_764),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_825),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_825),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_919),
.B(n_229),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_784),
.Y(n_1158)
);

BUFx8_ASAP7_75t_SL g1159 ( 
.A(n_764),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_832),
.B(n_18),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_742),
.B(n_193),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_767),
.A2(n_204),
.B1(n_199),
.B2(n_193),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_828),
.A2(n_204),
.B1(n_194),
.B2(n_198),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_821),
.B(n_193),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_919),
.B(n_296),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_860),
.A2(n_193),
.B(n_199),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_881),
.B(n_296),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_740),
.B(n_193),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_854),
.B(n_193),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_853),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_803),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_936),
.B(n_204),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_853),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_867),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_867),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_869),
.Y(n_1176)
);

AND3x1_ASAP7_75t_SL g1177 ( 
.A(n_847),
.B(n_19),
.C(n_22),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_881),
.B(n_296),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_869),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_784),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_845),
.B(n_877),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_883),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_883),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_838),
.B(n_199),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_782),
.B(n_199),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_890),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_719),
.B(n_204),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_890),
.B(n_204),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_717),
.Y(n_1189)
);

AOI22x1_ASAP7_75t_L g1190 ( 
.A1(n_708),
.A2(n_199),
.B1(n_293),
.B2(n_291),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_898),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_898),
.B(n_199),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_900),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_832),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_784),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_900),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_935),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_881),
.B(n_296),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_784),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_935),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_736),
.B(n_296),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_790),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_873),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_717),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_864),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_717),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_796),
.A2(n_296),
.B1(n_293),
.B2(n_291),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_849),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_930),
.B(n_194),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_891),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_938),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_889),
.B(n_194),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_938),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_892),
.A2(n_194),
.B1(n_198),
.B2(n_291),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_897),
.B(n_194),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_906),
.Y(n_1216)
);

INVx3_ASAP7_75t_SL g1217 ( 
.A(n_866),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_803),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_702),
.B(n_194),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_938),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_873),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_736),
.B(n_296),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_939),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_939),
.Y(n_1224)
);

OR2x6_ASAP7_75t_L g1225 ( 
.A(n_755),
.B(n_296),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_939),
.B(n_194),
.Y(n_1226)
);

NAND2xp33_ASAP7_75t_SL g1227 ( 
.A(n_829),
.B(n_293),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_717),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_892),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_903),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_830),
.B(n_194),
.Y(n_1231)
);

AND3x2_ASAP7_75t_SL g1232 ( 
.A(n_847),
.B(n_22),
.C(n_25),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_866),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_903),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_916),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_790),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_903),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_903),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_L g1239 ( 
.A1(n_1075),
.A2(n_807),
.B(n_855),
.C(n_856),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_944),
.B(n_909),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_949),
.A2(n_781),
.B1(n_769),
.B2(n_755),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1091),
.B(n_755),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1147),
.B(n_909),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1038),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1190),
.A2(n_870),
.B(n_766),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1038),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_948),
.A2(n_855),
.B(n_726),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1031),
.A2(n_775),
.B(n_872),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_943),
.A2(n_940),
.B(n_908),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1190),
.A2(n_918),
.B(n_925),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1136),
.A2(n_925),
.B(n_800),
.Y(n_1251)
);

AOI211x1_ASAP7_75t_L g1252 ( 
.A1(n_1141),
.A2(n_800),
.B(n_878),
.C(n_856),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_953),
.A2(n_887),
.B1(n_929),
.B2(n_755),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1074),
.B(n_790),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_985),
.A2(n_775),
.B(n_712),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1143),
.B(n_909),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1076),
.A2(n_805),
.B(n_862),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1076),
.A2(n_969),
.B(n_968),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_969),
.A2(n_805),
.B(n_862),
.Y(n_1259)
);

NAND2x1_ASAP7_75t_L g1260 ( 
.A(n_945),
.B(n_864),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1147),
.B(n_909),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1171),
.A2(n_844),
.B(n_878),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1227),
.A2(n_712),
.B(n_807),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_952),
.B(n_904),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1074),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1050),
.A2(n_772),
.B(n_843),
.C(n_887),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1171),
.A2(n_895),
.B(n_844),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1227),
.A2(n_772),
.B(n_788),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_950),
.B(n_689),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_947),
.B(n_689),
.Y(n_1270)
);

AOI21xp33_ASAP7_75t_L g1271 ( 
.A1(n_993),
.A2(n_929),
.B(n_926),
.Y(n_1271)
);

OAI21xp33_ASAP7_75t_SL g1272 ( 
.A1(n_994),
.A2(n_929),
.B(n_750),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_951),
.B(n_954),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1007),
.A2(n_788),
.B(n_773),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_961),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_961),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_956),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1064),
.A2(n_841),
.B(n_895),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_960),
.Y(n_1279)
);

AOI211x1_ASAP7_75t_L g1280 ( 
.A1(n_1141),
.A2(n_715),
.B(n_773),
.C(n_750),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1020),
.B(n_887),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1171),
.A2(n_1218),
.B(n_1029),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1052),
.Y(n_1283)
);

NAND2x1_ASAP7_75t_L g1284 ( 
.A(n_945),
.B(n_864),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_L g1285 ( 
.A1(n_1122),
.A2(n_1106),
.B1(n_1104),
.B2(n_1232),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_946),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1043),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1218),
.A2(n_901),
.B(n_899),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1011),
.A2(n_715),
.B(n_929),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_960),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_970),
.B(n_689),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1020),
.B(n_887),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1070),
.A2(n_896),
.B(n_885),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1045),
.A2(n_1181),
.B(n_1016),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_998),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_989),
.B(n_709),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_964),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_997),
.B(n_709),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_956),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1100),
.B(n_887),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1091),
.B(n_709),
.Y(n_1301)
);

O2A1O1Ixp5_ASAP7_75t_L g1302 ( 
.A1(n_1075),
.A2(n_922),
.B(n_924),
.C(n_874),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1225),
.A2(n_803),
.B(n_736),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_986),
.B(n_871),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1218),
.A2(n_913),
.B(n_910),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1029),
.A2(n_917),
.B(n_861),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1052),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_962),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1166),
.A2(n_876),
.B(n_729),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_998),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1119),
.A2(n_1126),
.B(n_1219),
.Y(n_1311)
);

AOI21x1_ASAP7_75t_SL g1312 ( 
.A1(n_1000),
.A2(n_886),
.B(n_829),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_965),
.B(n_727),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1119),
.A2(n_876),
.B(n_729),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1148),
.B(n_727),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1074),
.B(n_1205),
.Y(n_1316)
);

OR2x6_ASAP7_75t_L g1317 ( 
.A(n_980),
.B(n_803),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1148),
.B(n_727),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1140),
.A2(n_928),
.B(n_920),
.C(n_822),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_945),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1074),
.B(n_928),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1169),
.A2(n_933),
.B(n_942),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1017),
.B(n_727),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1059),
.A2(n_790),
.B(n_928),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_957),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_976),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_962),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_980),
.B(n_802),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1207),
.A2(n_1209),
.B(n_1144),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1017),
.B(n_737),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1043),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1033),
.B(n_737),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1164),
.A2(n_942),
.B(n_864),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1074),
.B(n_790),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1225),
.A2(n_802),
.B(n_818),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1033),
.B(n_737),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1035),
.B(n_737),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1184),
.A2(n_185),
.B(n_886),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1010),
.A2(n_928),
.B(n_822),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1119),
.A2(n_880),
.B(n_185),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1126),
.A2(n_880),
.B(n_185),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1028),
.A2(n_880),
.B(n_928),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1035),
.B(n_880),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1205),
.A2(n_822),
.B(n_818),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1107),
.A2(n_818),
.A3(n_802),
.B(n_880),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1001),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_955),
.B(n_873),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1205),
.A2(n_185),
.B(n_291),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1126),
.A2(n_185),
.B(n_291),
.Y(n_1349)
);

NOR2x1_ASAP7_75t_SL g1350 ( 
.A(n_1205),
.B(n_293),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_958),
.B(n_28),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_964),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1205),
.A2(n_293),
.B(n_291),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1069),
.A2(n_293),
.B(n_291),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_980),
.A2(n_1225),
.B(n_1157),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1212),
.A2(n_1215),
.B(n_1090),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_980),
.A2(n_293),
.B(n_291),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1192),
.A2(n_293),
.B(n_291),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1082),
.B(n_28),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1043),
.Y(n_1360)
);

INVx3_ASAP7_75t_SL g1361 ( 
.A(n_946),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1225),
.A2(n_293),
.B(n_284),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1113),
.A2(n_284),
.B(n_283),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1028),
.A2(n_29),
.B(n_30),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1185),
.A2(n_284),
.B(n_283),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1091),
.B(n_284),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_967),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1139),
.A2(n_284),
.B(n_283),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1139),
.A2(n_284),
.B(n_283),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_999),
.A2(n_284),
.B1(n_283),
.B2(n_279),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_975),
.A2(n_284),
.B(n_283),
.Y(n_1371)
);

NOR2x1_ASAP7_75t_L g1372 ( 
.A(n_1093),
.B(n_1115),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1226),
.A2(n_284),
.B(n_283),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1165),
.A2(n_284),
.B(n_283),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1144),
.A2(n_283),
.B(n_279),
.Y(n_1375)
);

AOI211x1_ASAP7_75t_L g1376 ( 
.A1(n_1042),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1077),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_981),
.B(n_33),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1167),
.A2(n_283),
.B(n_279),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1098),
.A2(n_279),
.B(n_273),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1098),
.A2(n_978),
.B(n_972),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_992),
.B(n_34),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1178),
.A2(n_279),
.B(n_273),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1003),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1187),
.A2(n_36),
.B(n_37),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_999),
.A2(n_279),
.B1(n_273),
.B2(n_240),
.Y(n_1386)
);

O2A1O1Ixp5_ASAP7_75t_L g1387 ( 
.A1(n_1198),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1019),
.B(n_39),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_972),
.A2(n_279),
.B(n_273),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_992),
.B(n_39),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1003),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_978),
.A2(n_279),
.B(n_273),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_R g1393 ( 
.A(n_1233),
.B(n_279),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_967),
.A2(n_41),
.B(n_42),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1104),
.B(n_41),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1106),
.B(n_42),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1131),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_983),
.A2(n_279),
.B(n_273),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_977),
.A2(n_273),
.B(n_240),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_957),
.A2(n_1027),
.B(n_966),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_996),
.B(n_44),
.Y(n_1401)
);

INVx8_ASAP7_75t_L g1402 ( 
.A(n_1168),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1187),
.A2(n_46),
.B(n_47),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_957),
.B(n_273),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_973),
.B(n_46),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_983),
.A2(n_229),
.B(n_240),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_966),
.B(n_229),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_L g1408 ( 
.A(n_1093),
.B(n_229),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_966),
.A2(n_229),
.B(n_240),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_984),
.A2(n_229),
.B(n_240),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1057),
.A2(n_229),
.B(n_240),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1009),
.B(n_229),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1210),
.B(n_194),
.Y(n_1413)
);

INVx5_ASAP7_75t_L g1414 ( 
.A(n_1003),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1003),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_984),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_959),
.A2(n_229),
.B(n_240),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1027),
.B(n_229),
.Y(n_1418)
);

O2A1O1Ixp5_ASAP7_75t_L g1419 ( 
.A1(n_1160),
.A2(n_273),
.B(n_240),
.C(n_235),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_995),
.A2(n_273),
.B(n_240),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_995),
.A2(n_240),
.B(n_235),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1027),
.A2(n_230),
.B(n_235),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1002),
.A2(n_230),
.B(n_235),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1210),
.B(n_194),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1002),
.A2(n_230),
.B(n_235),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_973),
.B(n_194),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1216),
.B(n_194),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_973),
.B(n_194),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1053),
.A2(n_230),
.B(n_235),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1063),
.A2(n_230),
.B1(n_235),
.B2(n_194),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1015),
.B(n_198),
.Y(n_1431)
);

AOI21x1_ASAP7_75t_L g1432 ( 
.A1(n_977),
.A2(n_230),
.B(n_235),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1063),
.A2(n_230),
.B1(n_235),
.B2(n_198),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1001),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1053),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1004),
.A2(n_230),
.B(n_189),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_982),
.A2(n_230),
.B(n_198),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1053),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1015),
.B(n_198),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1078),
.A2(n_1125),
.B(n_1097),
.Y(n_1440)
);

AND2x2_ASAP7_75t_SL g1441 ( 
.A(n_1232),
.B(n_230),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1078),
.A2(n_184),
.B(n_180),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_990),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_990),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1102),
.A2(n_198),
.B1(n_189),
.B2(n_180),
.C(n_184),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1078),
.A2(n_184),
.B(n_180),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1216),
.B(n_198),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1004),
.A2(n_1041),
.B(n_1018),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1003),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1015),
.B(n_198),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1083),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1032),
.B(n_198),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1071),
.A2(n_198),
.B(n_189),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1018),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1097),
.B(n_198),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1032),
.B(n_198),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1032),
.B(n_198),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1097),
.A2(n_184),
.B(n_189),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1049),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1235),
.B(n_180),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1125),
.B(n_1195),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1041),
.A2(n_180),
.B(n_189),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1047),
.A2(n_180),
.B(n_189),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1025),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1125),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1047),
.A2(n_180),
.B(n_189),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1235),
.B(n_180),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1081),
.A2(n_180),
.B(n_189),
.C(n_184),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1049),
.B(n_180),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1067),
.B(n_184),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_987),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1195),
.A2(n_184),
.B(n_189),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1056),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1025),
.Y(n_1474)
);

INVx8_ASAP7_75t_L g1475 ( 
.A(n_1168),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_SL g1476 ( 
.A1(n_991),
.A2(n_180),
.B(n_189),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_991),
.A2(n_189),
.B(n_180),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1094),
.B(n_180),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1123),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1025),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1056),
.Y(n_1481)
);

BUFx4_ASAP7_75t_SL g1482 ( 
.A(n_1036),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1067),
.B(n_184),
.Y(n_1483)
);

AOI21xp33_ASAP7_75t_L g1484 ( 
.A1(n_1057),
.A2(n_180),
.B(n_189),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1060),
.A2(n_180),
.B(n_189),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1006),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1067),
.B(n_184),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_L g1488 ( 
.A(n_1115),
.B(n_189),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_988),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_979),
.B(n_184),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1006),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1060),
.A2(n_189),
.B(n_184),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_979),
.B(n_184),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1061),
.A2(n_184),
.B(n_1065),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1061),
.A2(n_184),
.B(n_1065),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1195),
.Y(n_1496)
);

INVx3_ASAP7_75t_SL g1497 ( 
.A(n_1009),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1055),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1025),
.B(n_1026),
.Y(n_1499)
);

NOR4xp25_ASAP7_75t_L g1500 ( 
.A(n_1232),
.B(n_184),
.C(n_1134),
.D(n_1229),
.Y(n_1500)
);

NOR2x1_ASAP7_75t_SL g1501 ( 
.A(n_1025),
.B(n_184),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1066),
.A2(n_1231),
.B(n_1172),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1072),
.A2(n_1089),
.B(n_1073),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1037),
.B(n_1137),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_SL g1505 ( 
.A1(n_1008),
.A2(n_1014),
.B(n_1013),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_963),
.B(n_971),
.Y(n_1506)
);

AO31x2_ASAP7_75t_L g1507 ( 
.A1(n_1008),
.A2(n_1114),
.A3(n_1116),
.B(n_1111),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1137),
.B(n_971),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1072),
.A2(n_1197),
.B(n_1073),
.Y(n_1509)
);

INVx5_ASAP7_75t_L g1510 ( 
.A(n_1026),
.Y(n_1510)
);

CKINVDCx8_ASAP7_75t_R g1511 ( 
.A(n_1208),
.Y(n_1511)
);

AOI21x1_ASAP7_75t_SL g1512 ( 
.A1(n_1057),
.A2(n_1084),
.B(n_1087),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1089),
.A2(n_1197),
.B(n_1110),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_963),
.B(n_974),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1081),
.A2(n_1145),
.B(n_1084),
.Y(n_1515)
);

AOI221x1_ASAP7_75t_L g1516 ( 
.A1(n_1087),
.A2(n_1034),
.B1(n_1130),
.B2(n_1127),
.C(n_1120),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1055),
.B(n_1150),
.Y(n_1517)
);

O2A1O1Ixp5_ASAP7_75t_L g1518 ( 
.A1(n_1068),
.A2(n_1133),
.B(n_1234),
.C(n_1230),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1110),
.A2(n_1117),
.B(n_1124),
.Y(n_1519)
);

NAND2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1026),
.B(n_1040),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_963),
.B(n_974),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1013),
.A2(n_1127),
.B(n_1130),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1117),
.A2(n_1138),
.B(n_1124),
.Y(n_1523)
);

INVx5_ASAP7_75t_L g1524 ( 
.A(n_1026),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1138),
.A2(n_1179),
.B(n_1170),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1522),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1242),
.B(n_1168),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1317),
.B(n_1168),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1245),
.A2(n_1258),
.B(n_1432),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1266),
.A2(n_1081),
.B(n_1084),
.C(n_1030),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1390),
.B(n_1118),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1273),
.B(n_1044),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1522),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1244),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1514),
.B(n_1194),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1522),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1489),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1014),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1244),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1303),
.B(n_1094),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1390),
.B(n_1005),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1269),
.B(n_1046),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1507),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1287),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1240),
.B(n_1051),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1248),
.A2(n_1063),
.B(n_1096),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1504),
.A2(n_1154),
.B1(n_1208),
.B2(n_1088),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1507),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1255),
.A2(n_1096),
.B(n_1094),
.Y(n_1549)
);

NAND2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1265),
.B(n_1026),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1507),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1286),
.B(n_1233),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1317),
.B(n_1094),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1382),
.B(n_1395),
.Y(n_1554)
);

OR2x2_ASAP7_75t_SL g1555 ( 
.A(n_1401),
.B(n_1382),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1395),
.B(n_1005),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1266),
.A2(n_1030),
.B(n_1021),
.C(n_1022),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1361),
.A2(n_1217),
.B(n_1154),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1264),
.A2(n_1217),
.B1(n_1214),
.B2(n_1088),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1317),
.B(n_1096),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1417),
.A2(n_1096),
.B(n_1202),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1317),
.B(n_1237),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1316),
.A2(n_1319),
.B(n_1289),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1287),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1328),
.B(n_1237),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1287),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1507),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1359),
.B(n_1068),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1265),
.B(n_1316),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1507),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1505),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1319),
.A2(n_1058),
.B(n_1158),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1294),
.B(n_1054),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1441),
.A2(n_1036),
.B1(n_1068),
.B2(n_1123),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1328),
.B(n_1238),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1459),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1321),
.A2(n_1324),
.B(n_1303),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1482),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1321),
.A2(n_1058),
.B(n_1180),
.Y(n_1579)
);

AND2x2_ASAP7_75t_SL g1580 ( 
.A(n_1441),
.B(n_1040),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1287),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1275),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1397),
.A2(n_1129),
.B(n_1123),
.C(n_1146),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1295),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1276),
.Y(n_1585)
);

NOR2xp67_ASAP7_75t_L g1586 ( 
.A(n_1451),
.B(n_1238),
.Y(n_1586)
);

O2A1O1Ixp5_ASAP7_75t_L g1587 ( 
.A1(n_1329),
.A2(n_1120),
.B(n_1021),
.C(n_1022),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1331),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1331),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1290),
.B(n_1024),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1399),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1459),
.Y(n_1592)
);

BUFx4_ASAP7_75t_SL g1593 ( 
.A(n_1286),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1268),
.A2(n_1236),
.B(n_1142),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1364),
.A2(n_1105),
.B1(n_1109),
.B2(n_1092),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1297),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1352),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1385),
.A2(n_1039),
.B1(n_1111),
.B2(n_1024),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1357),
.A2(n_1236),
.B(n_1142),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1295),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1367),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1291),
.B(n_1034),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1304),
.B(n_1039),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1443),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1346),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1396),
.B(n_1012),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1328),
.B(n_1040),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1279),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1270),
.B(n_1351),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1396),
.B(n_1012),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1274),
.A2(n_1236),
.B(n_1040),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1444),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1256),
.B(n_1023),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1377),
.B(n_1114),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1397),
.A2(n_1132),
.B(n_1116),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1346),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1265),
.A2(n_1236),
.B(n_1040),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1486),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1331),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1434),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1290),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1265),
.A2(n_1236),
.B(n_1180),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1313),
.B(n_1150),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1331),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1310),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1310),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1265),
.A2(n_1180),
.B(n_1142),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1378),
.B(n_1152),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1335),
.A2(n_1180),
.B(n_1142),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1403),
.A2(n_1146),
.B(n_1129),
.C(n_1177),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1326),
.B(n_1152),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1511),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1300),
.A2(n_1471),
.B1(n_1515),
.B2(n_1511),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1360),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1301),
.B(n_1023),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1491),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1448),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1246),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1498),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1360),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1249),
.A2(n_1079),
.B(n_1172),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1498),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1360),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1506),
.B(n_1347),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1360),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1301),
.B(n_1095),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1335),
.A2(n_1142),
.B(n_1058),
.Y(n_1647)
);

INVx5_ASAP7_75t_L g1648 ( 
.A(n_1328),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1301),
.B(n_1095),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1419),
.A2(n_1199),
.B(n_1058),
.Y(n_1650)
);

BUFx12f_ASAP7_75t_L g1651 ( 
.A(n_1246),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1384),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1242),
.B(n_1048),
.Y(n_1653)
);

OR2x6_ASAP7_75t_SL g1654 ( 
.A(n_1388),
.B(n_1405),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1384),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1361),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1272),
.B(n_1146),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1285),
.B(n_1095),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1339),
.A2(n_1202),
.B(n_1058),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1372),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1241),
.A2(n_1079),
.B1(n_1085),
.B2(n_1135),
.Y(n_1661)
);

INVx3_ASAP7_75t_SL g1662 ( 
.A(n_1497),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1497),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1448),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1300),
.A2(n_1263),
.B(n_1342),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1384),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1517),
.Y(n_1667)
);

CKINVDCx11_ASAP7_75t_R g1668 ( 
.A(n_1283),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1508),
.A2(n_1079),
.B1(n_1085),
.B2(n_1135),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1517),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1277),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1307),
.A2(n_1085),
.B1(n_1135),
.B2(n_1129),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1277),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1391),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1243),
.B(n_1186),
.Y(n_1675)
);

INVx6_ASAP7_75t_L g1676 ( 
.A(n_1391),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1283),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1261),
.B(n_1186),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1468),
.A2(n_1199),
.B(n_1062),
.Y(n_1679)
);

INVx2_ASAP7_75t_SL g1680 ( 
.A(n_1307),
.Y(n_1680)
);

INVxp67_ASAP7_75t_SL g1681 ( 
.A(n_1399),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1502),
.A2(n_1048),
.B1(n_1080),
.B2(n_1221),
.Y(n_1682)
);

CKINVDCx16_ASAP7_75t_R g1683 ( 
.A(n_1412),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1271),
.B(n_1080),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1299),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1285),
.B(n_1228),
.Y(n_1686)
);

BUFx4f_ASAP7_75t_L g1687 ( 
.A(n_1384),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1468),
.A2(n_1062),
.B(n_1180),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1258),
.A2(n_1062),
.B(n_1199),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1242),
.B(n_1323),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1299),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1503),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1500),
.B(n_1228),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1387),
.B(n_1108),
.C(n_1128),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1330),
.B(n_1183),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1516),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1296),
.B(n_1183),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1503),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1308),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1332),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1469),
.B(n_1206),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1336),
.B(n_1156),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1280),
.A2(n_1203),
.B1(n_1221),
.B2(n_1151),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1474),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1247),
.B(n_1062),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1298),
.B(n_1156),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1308),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1344),
.A2(n_1062),
.B(n_1158),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1474),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1327),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1315),
.B(n_1191),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1327),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1253),
.A2(n_1112),
.B(n_1121),
.C(n_1101),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1469),
.B(n_1189),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1416),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1413),
.B(n_1189),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1278),
.A2(n_1199),
.B(n_1202),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1474),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1394),
.A2(n_1159),
.B1(n_1175),
.B2(n_1176),
.Y(n_1719)
);

INVxp67_ASAP7_75t_SL g1720 ( 
.A(n_1399),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1337),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1362),
.A2(n_1199),
.B(n_1202),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1282),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1416),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1318),
.B(n_1182),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1454),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1474),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1391),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1454),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1518),
.A2(n_1202),
.B(n_1158),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1302),
.A2(n_1151),
.B(n_1161),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_SL g1732 ( 
.A(n_1415),
.B(n_1159),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1473),
.Y(n_1733)
);

AO21x1_ASAP7_75t_L g1734 ( 
.A1(n_1281),
.A2(n_1182),
.B(n_1200),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1356),
.B(n_1191),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1293),
.A2(n_1158),
.B(n_1201),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1473),
.B(n_1200),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1509),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1415),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1415),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1355),
.B(n_1158),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1481),
.B(n_1155),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1481),
.B(n_1155),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1509),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1391),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1282),
.B(n_1203),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1343),
.B(n_1174),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1366),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1449),
.B(n_1464),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1329),
.A2(n_1201),
.B(n_1222),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1499),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1333),
.A2(n_1201),
.B(n_1222),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1513),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1513),
.Y(n_1754)
);

NOR2xp67_ASAP7_75t_L g1755 ( 
.A(n_1449),
.B(n_1151),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1356),
.B(n_1281),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1449),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1413),
.B(n_1424),
.Y(n_1758)
);

NAND2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1391),
.B(n_1204),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1464),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1353),
.A2(n_1222),
.B(n_1161),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1368),
.A2(n_1161),
.B(n_1223),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1322),
.B(n_1173),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_SL g1764 ( 
.A(n_1292),
.B(n_1193),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1464),
.Y(n_1765)
);

O2A1O1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1292),
.A2(n_1103),
.B(n_1193),
.C(n_1223),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1519),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1424),
.B(n_1196),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1320),
.B(n_1206),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1499),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1530),
.A2(n_1239),
.B(n_1350),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1576),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1600),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1593),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1537),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1576),
.B(n_1394),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1592),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1656),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1582),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1585),
.Y(n_1780)
);

A2O1A1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1530),
.A2(n_1402),
.B(n_1475),
.C(n_1257),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1592),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1644),
.B(n_1394),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1556),
.B(n_1408),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1644),
.B(n_1376),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1648),
.B(n_1414),
.Y(n_1786)
);

CKINVDCx14_ASAP7_75t_R g1787 ( 
.A(n_1668),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1633),
.A2(n_1402),
.B1(n_1475),
.B2(n_1478),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1541),
.B(n_1338),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1536),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1536),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1639),
.B(n_1381),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1626),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_SL g1794 ( 
.A(n_1662),
.B(n_1260),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1656),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1604),
.B(n_1338),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1555),
.A2(n_1252),
.B1(n_1478),
.B2(n_1402),
.Y(n_1797)
);

O2A1O1Ixp5_ASAP7_75t_L g1798 ( 
.A1(n_1705),
.A2(n_1763),
.B(n_1563),
.C(n_1577),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1604),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1557),
.A2(n_1354),
.B(n_1400),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1596),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1618),
.B(n_1338),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1654),
.A2(n_1478),
.B1(n_1475),
.B2(n_1402),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1618),
.B(n_1262),
.Y(n_1804)
);

A2O1A1Ixp33_ASAP7_75t_SL g1805 ( 
.A1(n_1719),
.A2(n_1320),
.B(n_1438),
.C(n_1465),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1636),
.B(n_1262),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1700),
.B(n_1721),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_SL g1808 ( 
.A(n_1534),
.B(n_1475),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1609),
.B(n_1479),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1636),
.B(n_1267),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1597),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1538),
.B(n_1381),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1667),
.B(n_1267),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1639),
.B(n_1288),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1648),
.B(n_1311),
.Y(n_1815)
);

OR2x6_ASAP7_75t_SL g1816 ( 
.A(n_1574),
.B(n_1512),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1557),
.A2(n_1440),
.B(n_1284),
.Y(n_1817)
);

NOR2xp67_ASAP7_75t_L g1818 ( 
.A(n_1558),
.B(n_1680),
.Y(n_1818)
);

AO31x2_ASAP7_75t_L g1819 ( 
.A1(n_1734),
.A2(n_1370),
.A3(n_1386),
.B(n_1501),
.Y(n_1819)
);

BUFx4f_ASAP7_75t_SL g1820 ( 
.A(n_1651),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1601),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1663),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1612),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1730),
.A2(n_1369),
.B(n_1368),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1621),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1670),
.B(n_1311),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1572),
.A2(n_1761),
.B(n_1705),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1580),
.B(n_1288),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1535),
.B(n_1447),
.Y(n_1829)
);

O2A1O1Ixp5_ASAP7_75t_L g1830 ( 
.A1(n_1763),
.A2(n_1437),
.B(n_1435),
.C(n_1496),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1736),
.A2(n_1647),
.B(n_1629),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1532),
.B(n_1447),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1580),
.B(n_1305),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1573),
.B(n_1460),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1602),
.B(n_1460),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1668),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1526),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1648),
.B(n_1305),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1630),
.A2(n_1559),
.B(n_1615),
.C(n_1583),
.Y(n_1839)
);

OA21x2_ASAP7_75t_L g1840 ( 
.A1(n_1529),
.A2(n_1245),
.B(n_1259),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1665),
.A2(n_1369),
.B(n_1368),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1593),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1642),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1648),
.B(n_1414),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1533),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1606),
.B(n_1366),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1595),
.B(n_1414),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1551),
.Y(n_1848)
);

OR2x6_ASAP7_75t_SL g1849 ( 
.A(n_1638),
.B(n_1427),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1613),
.B(n_1257),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1590),
.B(n_1519),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1630),
.A2(n_1478),
.B1(n_1510),
.B2(n_1414),
.Y(n_1852)
);

AOI21x1_ASAP7_75t_SL g1853 ( 
.A1(n_1746),
.A2(n_1366),
.B(n_1490),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1545),
.B(n_1467),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1747),
.B(n_1467),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1608),
.B(n_1493),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1610),
.B(n_1523),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1756),
.B(n_1523),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1661),
.A2(n_1435),
.B1(n_1325),
.B2(n_1320),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1534),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1746),
.B(n_1414),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1531),
.B(n_1204),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1747),
.B(n_1525),
.Y(n_1863)
);

CKINVDCx20_ASAP7_75t_R g1864 ( 
.A(n_1638),
.Y(n_1864)
);

AOI32xp33_ASAP7_75t_L g1865 ( 
.A1(n_1598),
.A2(n_1488),
.A3(n_1445),
.B1(n_1496),
.B2(n_1435),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1554),
.B(n_1520),
.Y(n_1866)
);

OAI21x1_ASAP7_75t_SL g1867 ( 
.A1(n_1764),
.A2(n_1476),
.B(n_1477),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1570),
.B(n_1525),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1542),
.B(n_1153),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1686),
.B(n_1543),
.Y(n_1870)
);

OR2x6_ASAP7_75t_SL g1871 ( 
.A(n_1677),
.B(n_1427),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1598),
.A2(n_1524),
.B1(n_1510),
.B2(n_1480),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1735),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1543),
.B(n_1259),
.Y(n_1874)
);

NOR2xp67_ASAP7_75t_L g1875 ( 
.A(n_1651),
.B(n_1325),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1548),
.B(n_1306),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1548),
.B(n_1306),
.Y(n_1877)
);

O2A1O1Ixp5_ASAP7_75t_L g1878 ( 
.A1(n_1546),
.A2(n_1325),
.B(n_1496),
.C(n_1438),
.Y(n_1878)
);

OR2x6_ASAP7_75t_SL g1879 ( 
.A(n_1677),
.B(n_1426),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1690),
.B(n_1153),
.Y(n_1880)
);

NAND2x1p5_ASAP7_75t_L g1881 ( 
.A(n_1674),
.B(n_1480),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1690),
.B(n_1170),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1600),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1567),
.B(n_1345),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1603),
.B(n_1179),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1567),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1662),
.B(n_1428),
.Y(n_1887)
);

NAND2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1674),
.B(n_1480),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1561),
.A2(n_1369),
.B(n_1334),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1595),
.A2(n_1250),
.B(n_1309),
.C(n_1480),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1671),
.Y(n_1891)
);

A2O1A1Ixp33_ASAP7_75t_SL g1892 ( 
.A1(n_1719),
.A2(n_1438),
.B(n_1465),
.C(n_1453),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1695),
.B(n_1196),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1625),
.Y(n_1894)
);

NAND2x1p5_ASAP7_75t_L g1895 ( 
.A(n_1728),
.B(n_1480),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1637),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1562),
.B(n_1345),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1702),
.B(n_1211),
.Y(n_1898)
);

OR2x6_ASAP7_75t_SL g1899 ( 
.A(n_1709),
.B(n_1431),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1599),
.A2(n_1334),
.B(n_1254),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1673),
.Y(n_1901)
);

A2O1A1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1549),
.A2(n_1250),
.B(n_1309),
.C(n_1510),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1660),
.B(n_1439),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1620),
.B(n_1345),
.Y(n_1904)
);

OA21x2_ASAP7_75t_L g1905 ( 
.A1(n_1587),
.A2(n_1365),
.B(n_1358),
.Y(n_1905)
);

NOR2xp67_ASAP7_75t_L g1906 ( 
.A(n_1663),
.B(n_1465),
.Y(n_1906)
);

NAND2x1p5_ASAP7_75t_L g1907 ( 
.A(n_1728),
.B(n_1510),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1562),
.B(n_1345),
.Y(n_1908)
);

O2A1O1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1628),
.A2(n_1450),
.B(n_1456),
.C(n_1457),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1722),
.A2(n_1254),
.B(n_1363),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1568),
.B(n_1211),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1746),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1562),
.B(n_1251),
.Y(n_1913)
);

O2A1O1Ixp5_ASAP7_75t_L g1914 ( 
.A1(n_1717),
.A2(n_1484),
.B(n_1452),
.C(n_1430),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1915)
);

INVxp67_ASAP7_75t_L g1916 ( 
.A(n_1584),
.Y(n_1916)
);

BUFx12f_ASAP7_75t_L g1917 ( 
.A(n_1539),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1616),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1723),
.B(n_1251),
.Y(n_1919)
);

AOI21x1_ASAP7_75t_SL g1920 ( 
.A1(n_1696),
.A2(n_1393),
.B(n_1487),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1682),
.A2(n_1520),
.B(n_1461),
.C(n_1483),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1568),
.B(n_1224),
.Y(n_1922)
);

A2O1A1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1750),
.A2(n_1524),
.B(n_1510),
.C(n_1314),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1723),
.B(n_1373),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1565),
.B(n_1373),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1626),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1614),
.B(n_1495),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1637),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1565),
.B(n_1365),
.Y(n_1929)
);

O2A1O1Ixp5_ASAP7_75t_L g1930 ( 
.A1(n_1641),
.A2(n_1433),
.B(n_1374),
.C(n_1470),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1616),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1623),
.B(n_1213),
.Y(n_1932)
);

OA21x2_ASAP7_75t_L g1933 ( 
.A1(n_1587),
.A2(n_1358),
.B(n_1371),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1575),
.B(n_1380),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1631),
.B(n_1494),
.Y(n_1935)
);

NOR2xp67_ASAP7_75t_L g1936 ( 
.A(n_1578),
.B(n_1524),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1675),
.B(n_1224),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1678),
.B(n_1220),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1575),
.B(n_1380),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1664),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1697),
.B(n_1220),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1575),
.B(n_1495),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1611),
.A2(n_1524),
.B(n_1409),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1605),
.Y(n_1944)
);

O2A1O1Ixp33_ASAP7_75t_L g1945 ( 
.A1(n_1713),
.A2(n_1731),
.B(n_1703),
.C(n_1696),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1607),
.B(n_1314),
.Y(n_1946)
);

O2A1O1Ixp5_ASAP7_75t_L g1947 ( 
.A1(n_1657),
.A2(n_1379),
.B(n_1383),
.C(n_1213),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1685),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1607),
.B(n_1371),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1607),
.B(n_1341),
.Y(n_1950)
);

A2O1A1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1657),
.A2(n_1429),
.B(n_1422),
.C(n_1340),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1635),
.B(n_1658),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1706),
.B(n_1461),
.Y(n_1953)
);

BUFx4_ASAP7_75t_R g1954 ( 
.A(n_1632),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1691),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1528),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1725),
.B(n_1188),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1699),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1553),
.B(n_1341),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1586),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1553),
.B(n_1494),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1664),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_SL g1963 ( 
.A(n_1539),
.B(n_1188),
.Y(n_1963)
);

O2A1O1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1694),
.A2(n_1766),
.B(n_1684),
.C(n_1732),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1692),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1692),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1528),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1679),
.A2(n_1340),
.B(n_1418),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1553),
.B(n_1398),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1560),
.B(n_1398),
.Y(n_1970)
);

BUFx12f_ASAP7_75t_L g1971 ( 
.A(n_1544),
.Y(n_1971)
);

AND2x2_ASAP7_75t_SL g1972 ( 
.A(n_1683),
.B(n_1312),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1560),
.B(n_1389),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1528),
.Y(n_1974)
);

CKINVDCx16_ASAP7_75t_R g1975 ( 
.A(n_1552),
.Y(n_1975)
);

NAND2x1p5_ASAP7_75t_L g1976 ( 
.A(n_1728),
.B(n_1375),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1646),
.B(n_1086),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1560),
.B(n_1389),
.Y(n_1978)
);

BUFx12f_ASAP7_75t_L g1979 ( 
.A(n_1544),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1739),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1698),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1711),
.B(n_1086),
.Y(n_1982)
);

A2O1A1Ixp33_ASAP7_75t_SL g1983 ( 
.A1(n_1684),
.A2(n_1149),
.B(n_1162),
.C(n_1442),
.Y(n_1983)
);

AND2x2_ASAP7_75t_SL g1984 ( 
.A(n_1527),
.B(n_1086),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1758),
.B(n_1421),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1707),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1698),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1594),
.A2(n_1446),
.B(n_1458),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1740),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1744),
.B(n_1420),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1710),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1741),
.Y(n_1992)
);

OA21x2_ASAP7_75t_L g1993 ( 
.A1(n_1591),
.A2(n_1681),
.B(n_1720),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1701),
.B(n_1420),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1753),
.B(n_1754),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1712),
.Y(n_1996)
);

INVxp67_ASAP7_75t_L g1997 ( 
.A(n_1714),
.Y(n_1997)
);

OA21x2_ASAP7_75t_L g1998 ( 
.A1(n_1591),
.A2(n_1375),
.B(n_1410),
.Y(n_1998)
);

OA21x2_ASAP7_75t_L g1999 ( 
.A1(n_1681),
.A2(n_1421),
.B(n_1425),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_SL g2000 ( 
.A1(n_1540),
.A2(n_1418),
.B(n_1407),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1571),
.B(n_1423),
.Y(n_2001)
);

NOR2x2_ASAP7_75t_L g2002 ( 
.A(n_1540),
.B(n_1411),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1716),
.B(n_1423),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1632),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1652),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1649),
.B(n_1455),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1715),
.B(n_1425),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1724),
.B(n_1410),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1694),
.A2(n_1455),
.B(n_1348),
.C(n_1407),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1748),
.B(n_1404),
.Y(n_2010)
);

BUFx4_ASAP7_75t_R g2011 ( 
.A(n_1751),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1653),
.B(n_1404),
.Y(n_2012)
);

BUFx3_ASAP7_75t_L g2013 ( 
.A(n_1652),
.Y(n_2013)
);

NOR2xp67_ASAP7_75t_L g2014 ( 
.A(n_1672),
.B(n_1472),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1837),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1837),
.Y(n_2016)
);

CKINVDCx6p67_ASAP7_75t_R g2017 ( 
.A(n_1836),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_R g2018 ( 
.A(n_1774),
.B(n_1709),
.Y(n_2018)
);

BUFx6f_ASAP7_75t_L g2019 ( 
.A(n_1773),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1845),
.Y(n_2020)
);

AO21x2_ASAP7_75t_L g2021 ( 
.A1(n_1902),
.A2(n_1689),
.B(n_1720),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1845),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1790),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1799),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1799),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1975),
.B(n_1669),
.Y(n_2026)
);

OAI21x1_ASAP7_75t_L g2027 ( 
.A1(n_1943),
.A2(n_1650),
.B(n_1738),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1807),
.B(n_1571),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1995),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1995),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1790),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1912),
.Y(n_2032)
);

NOR2xp67_ASAP7_75t_L g2033 ( 
.A(n_1912),
.B(n_1738),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1791),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1870),
.B(n_1767),
.Y(n_2035)
);

OAI21x1_ASAP7_75t_L g2036 ( 
.A1(n_1800),
.A2(n_1767),
.B(n_1569),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1791),
.Y(n_2037)
);

INVx3_ASAP7_75t_L g2038 ( 
.A(n_1912),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1815),
.B(n_1741),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1848),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1870),
.B(n_1741),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1775),
.B(n_1547),
.Y(n_2042)
);

OAI21x1_ASAP7_75t_L g2043 ( 
.A1(n_1824),
.A2(n_1831),
.B(n_1910),
.Y(n_2043)
);

OAI21x1_ASAP7_75t_L g2044 ( 
.A1(n_1841),
.A2(n_1569),
.B(n_1659),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1779),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1825),
.B(n_1693),
.Y(n_2046)
);

AO21x2_ASAP7_75t_L g2047 ( 
.A1(n_1902),
.A2(n_1708),
.B(n_1579),
.Y(n_2047)
);

INVxp67_ASAP7_75t_L g2048 ( 
.A(n_1894),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1780),
.Y(n_2049)
);

BUFx10_ASAP7_75t_L g2050 ( 
.A(n_1844),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1896),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1897),
.B(n_1540),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1801),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1811),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1821),
.Y(n_2055)
);

AND2x2_ASAP7_75t_SL g2056 ( 
.A(n_1984),
.B(n_1527),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1897),
.B(n_1769),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1823),
.Y(n_2058)
);

INVx4_ASAP7_75t_L g2059 ( 
.A(n_1954),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1896),
.Y(n_2060)
);

BUFx12f_ASAP7_75t_L g2061 ( 
.A(n_1860),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1873),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1772),
.B(n_1726),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1873),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1778),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1928),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_1778),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1891),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1901),
.Y(n_2069)
);

BUFx12f_ASAP7_75t_L g2070 ( 
.A(n_1860),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1948),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_1777),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1955),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1928),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1958),
.Y(n_2075)
);

AO21x2_ASAP7_75t_L g2076 ( 
.A1(n_1923),
.A2(n_1762),
.B(n_1688),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1940),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1986),
.Y(n_2078)
);

BUFx2_ASAP7_75t_R g2079 ( 
.A(n_1774),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1940),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1782),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1991),
.Y(n_2082)
);

BUFx2_ASAP7_75t_SL g2083 ( 
.A(n_1818),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1861),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1992),
.Y(n_2085)
);

OA21x2_ASAP7_75t_L g2086 ( 
.A1(n_1890),
.A2(n_1752),
.B(n_1406),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1861),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1962),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1908),
.B(n_1769),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1962),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1965),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_1980),
.Y(n_2092)
);

OAI21x1_ASAP7_75t_L g2093 ( 
.A1(n_1817),
.A2(n_1889),
.B(n_1968),
.Y(n_2093)
);

AO21x2_ASAP7_75t_L g2094 ( 
.A1(n_1923),
.A2(n_1890),
.B(n_1805),
.Y(n_2094)
);

AOI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_1839),
.A2(n_1653),
.B1(n_1768),
.B2(n_1733),
.C(n_1729),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1996),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1944),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1886),
.Y(n_2098)
);

OAI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_1964),
.A2(n_1640),
.B1(n_1645),
.B2(n_1588),
.C(n_1581),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_1803),
.A2(n_1640),
.B1(n_1588),
.B2(n_1581),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1965),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_1989),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1804),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_1926),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1861),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1966),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1773),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1966),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1804),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1981),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1981),
.Y(n_2111)
);

OAI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_1963),
.A2(n_1589),
.B1(n_1566),
.B2(n_1564),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1987),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1806),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1806),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_1776),
.B(n_1770),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1810),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1987),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1810),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1813),
.Y(n_2120)
);

INVx4_ASAP7_75t_L g2121 ( 
.A(n_1954),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1843),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1813),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1792),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1809),
.B(n_1769),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1878),
.A2(n_1392),
.B(n_1406),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1868),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_1826),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1826),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1868),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1858),
.Y(n_2131)
);

BUFx2_ASAP7_75t_L g2132 ( 
.A(n_1956),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_1814),
.B(n_1737),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2004),
.B(n_1787),
.Y(n_2134)
);

OAI21xp33_ASAP7_75t_SL g2135 ( 
.A1(n_1847),
.A2(n_1627),
.B(n_1622),
.Y(n_2135)
);

OA21x2_ASAP7_75t_L g2136 ( 
.A1(n_1798),
.A2(n_1392),
.B(n_1743),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1796),
.Y(n_2137)
);

INVxp67_ASAP7_75t_L g2138 ( 
.A(n_1944),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1842),
.Y(n_2139)
);

INVx4_ASAP7_75t_L g2140 ( 
.A(n_2011),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1796),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_1956),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_1904),
.B(n_1742),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1802),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1802),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_1857),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1851),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1815),
.B(n_1751),
.Y(n_2148)
);

BUFx6f_ASAP7_75t_SL g2149 ( 
.A(n_1795),
.Y(n_2149)
);

AO21x2_ASAP7_75t_L g2150 ( 
.A1(n_1805),
.A2(n_1617),
.B(n_1755),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1812),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2004),
.B(n_1643),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_1887),
.A2(n_2014),
.B1(n_1852),
.B2(n_1847),
.Y(n_2153)
);

INVxp67_ASAP7_75t_SL g2154 ( 
.A(n_1863),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1783),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_1956),
.Y(n_2156)
);

INVxp67_ASAP7_75t_SL g2157 ( 
.A(n_1960),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1884),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1884),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1908),
.B(n_1655),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1967),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1857),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_1795),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_1793),
.Y(n_2164)
);

OAI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_1788),
.A2(n_1619),
.B1(n_1589),
.B2(n_1566),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1850),
.B(n_1655),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2007),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_1827),
.A2(n_1687),
.B(n_1550),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1990),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1990),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1913),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1822),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1874),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_1793),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1913),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1874),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1919),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1919),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1993),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2008),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1993),
.Y(n_2181)
);

OA21x2_ASAP7_75t_L g2182 ( 
.A1(n_1771),
.A2(n_1436),
.B(n_1462),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1875),
.B(n_1566),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1993),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1850),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1929),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1929),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1876),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2001),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_1967),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2001),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1876),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1924),
.Y(n_2193)
);

BUFx10_ASAP7_75t_L g2194 ( 
.A(n_1844),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_1787),
.B(n_1643),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_1840),
.A2(n_1550),
.B(n_1436),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1924),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_1997),
.B(n_1727),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1877),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_1916),
.Y(n_2200)
);

OAI21x1_ASAP7_75t_L g2201 ( 
.A1(n_1840),
.A2(n_1485),
.B(n_1462),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1877),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1925),
.Y(n_2203)
);

AOI21x1_ASAP7_75t_L g2204 ( 
.A1(n_1900),
.A2(n_1749),
.B(n_1466),
.Y(n_2204)
);

OAI22xp33_ASAP7_75t_SL g2205 ( 
.A1(n_1849),
.A2(n_1676),
.B1(n_1759),
.B2(n_1645),
.Y(n_2205)
);

OR2x6_ASAP7_75t_L g2206 ( 
.A(n_2000),
.B(n_1676),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_1967),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1773),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1925),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1999),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1999),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1946),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1946),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1822),
.Y(n_2214)
);

AO21x2_ASAP7_75t_L g2215 ( 
.A1(n_1867),
.A2(n_1749),
.B(n_1463),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1946),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_1815),
.B(n_1749),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1953),
.B(n_1727),
.Y(n_2218)
);

OAI21x1_ASAP7_75t_L g2219 ( 
.A1(n_1840),
.A2(n_1485),
.B(n_1463),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1974),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1974),
.Y(n_2221)
);

INVx3_ASAP7_75t_L g2222 ( 
.A(n_1974),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1935),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1999),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1789),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1998),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1789),
.Y(n_2227)
);

OAI21x1_ASAP7_75t_L g2228 ( 
.A1(n_1947),
.A2(n_1466),
.B(n_1492),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_1773),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_L g2230 ( 
.A1(n_1988),
.A2(n_1492),
.B(n_1759),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1998),
.Y(n_2231)
);

INVx4_ASAP7_75t_SL g2232 ( 
.A(n_1820),
.Y(n_2232)
);

BUFx4f_ASAP7_75t_SL g2233 ( 
.A(n_1917),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_1838),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1949),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1838),
.B(n_1718),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1949),
.Y(n_2237)
);

OAI21xp5_ASAP7_75t_SL g2238 ( 
.A1(n_1945),
.A2(n_1589),
.B(n_1619),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_1931),
.Y(n_2239)
);

INVxp67_ASAP7_75t_L g2240 ( 
.A(n_1883),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1949),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1952),
.B(n_1718),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1838),
.Y(n_2243)
);

INVx1_ASAP7_75t_SL g2244 ( 
.A(n_1918),
.Y(n_2244)
);

AOI211xp5_ASAP7_75t_L g2245 ( 
.A1(n_1785),
.A2(n_1589),
.B(n_1624),
.C(n_1619),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_1931),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1998),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_1853),
.A2(n_1765),
.B(n_1760),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_1918),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1952),
.B(n_1652),
.Y(n_2250)
);

INVx1_ASAP7_75t_SL g2251 ( 
.A(n_2011),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1978),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1978),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1978),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1898),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1934),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1937),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1934),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1939),
.Y(n_2259)
);

BUFx3_ASAP7_75t_L g2260 ( 
.A(n_1883),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1939),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1938),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1969),
.Y(n_2263)
);

INVx2_ASAP7_75t_SL g2264 ( 
.A(n_1883),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1969),
.Y(n_2265)
);

INVx3_ASAP7_75t_L g2266 ( 
.A(n_1915),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1828),
.B(n_1652),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1970),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1970),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_1883),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_1828),
.B(n_1666),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_2005),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_1849),
.A2(n_1676),
.B1(n_1634),
.B2(n_1564),
.Y(n_2273)
);

BUFx2_ASAP7_75t_L g2274 ( 
.A(n_1959),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_1927),
.Y(n_2275)
);

OR2x6_ASAP7_75t_L g2276 ( 
.A(n_1781),
.B(n_1728),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_1833),
.B(n_1973),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1971),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1973),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1833),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1942),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_1915),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1893),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1942),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1834),
.B(n_1765),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1905),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1985),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2015),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2015),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2179),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2193),
.B(n_1994),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2179),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2277),
.B(n_1871),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2154),
.B(n_1855),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2181),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2277),
.B(n_1871),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2274),
.B(n_1866),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2274),
.B(n_1959),
.Y(n_2298)
);

BUFx2_ASAP7_75t_L g2299 ( 
.A(n_2140),
.Y(n_2299)
);

HB1xp67_ASAP7_75t_L g2300 ( 
.A(n_2275),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2181),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2184),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2105),
.B(n_2253),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2184),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_2061),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2129),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2193),
.B(n_2003),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2105),
.B(n_1959),
.Y(n_2308)
);

NAND4xp25_ASAP7_75t_L g2309 ( 
.A(n_2095),
.B(n_1892),
.C(n_1856),
.D(n_1865),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2253),
.B(n_1961),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2129),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2199),
.Y(n_2312)
);

OAI21xp5_ASAP7_75t_SL g2313 ( 
.A1(n_2238),
.A2(n_1781),
.B(n_1859),
.Y(n_2313)
);

BUFx2_ASAP7_75t_L g2314 ( 
.A(n_2140),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2199),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_2059),
.A2(n_1972),
.B1(n_1797),
.B2(n_1984),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2146),
.B(n_1961),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2016),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2185),
.B(n_1784),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2016),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2185),
.B(n_1950),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2155),
.B(n_1862),
.Y(n_2322)
);

NAND2x1_ASAP7_75t_L g2323 ( 
.A(n_2140),
.B(n_2059),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2020),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2202),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2155),
.B(n_1903),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2255),
.B(n_1835),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2202),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2209),
.B(n_2162),
.Y(n_2329)
);

BUFx2_ASAP7_75t_L g2330 ( 
.A(n_2140),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_2234),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2120),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2120),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2209),
.B(n_2162),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2020),
.Y(n_2335)
);

AO31x2_ASAP7_75t_L g2336 ( 
.A1(n_2210),
.A2(n_1872),
.A3(n_1951),
.B(n_2012),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2265),
.B(n_1950),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2265),
.B(n_1950),
.Y(n_2338)
);

CKINVDCx6p67_ASAP7_75t_R g2339 ( 
.A(n_2017),
.Y(n_2339)
);

AOI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_2059),
.A2(n_1972),
.B1(n_1917),
.B2(n_1977),
.Y(n_2340)
);

BUFx3_ASAP7_75t_L g2341 ( 
.A(n_2061),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_2276),
.B(n_1786),
.Y(n_2342)
);

INVx4_ASAP7_75t_L g2343 ( 
.A(n_2232),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2279),
.B(n_1899),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_2070),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2123),
.Y(n_2346)
);

BUFx3_ASAP7_75t_L g2347 ( 
.A(n_2070),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2022),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2123),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_2197),
.B(n_1829),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2022),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2279),
.B(n_1899),
.Y(n_2352)
);

NOR2x1_ASAP7_75t_R g2353 ( 
.A(n_2059),
.B(n_1842),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_SL g2354 ( 
.A1(n_2121),
.A2(n_1808),
.B1(n_1836),
.B2(n_1864),
.Y(n_2354)
);

OR2x6_ASAP7_75t_SL g2355 ( 
.A(n_2273),
.B(n_1922),
.Y(n_2355)
);

AOI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_2121),
.A2(n_1794),
.B1(n_2006),
.B2(n_1915),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2256),
.B(n_1879),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2127),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2127),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2256),
.B(n_1879),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2130),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2255),
.B(n_1911),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2130),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2258),
.B(n_1816),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_2121),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2034),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2258),
.B(n_1816),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2034),
.Y(n_2368)
);

AO31x2_ASAP7_75t_L g2369 ( 
.A1(n_2210),
.A2(n_1951),
.A3(n_1941),
.B(n_1885),
.Y(n_2369)
);

CKINVDCx20_ASAP7_75t_R g2370 ( 
.A(n_2017),
.Y(n_2370)
);

NAND2x1_ASAP7_75t_L g2371 ( 
.A(n_2121),
.B(n_1844),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2259),
.B(n_2013),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2023),
.Y(n_2373)
);

HB1xp67_ASAP7_75t_L g2374 ( 
.A(n_2072),
.Y(n_2374)
);

AOI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_2153),
.A2(n_2026),
.B1(n_2099),
.B2(n_2046),
.Y(n_2375)
);

BUFx3_ASAP7_75t_L g2376 ( 
.A(n_2172),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2056),
.A2(n_1794),
.B1(n_1846),
.B2(n_1634),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2259),
.B(n_2013),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2037),
.Y(n_2379)
);

AOI22xp33_ASAP7_75t_L g2380 ( 
.A1(n_2056),
.A2(n_1957),
.B1(n_1619),
.B2(n_1544),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2081),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2037),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2023),
.Y(n_2383)
);

AOI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_2056),
.A2(n_1566),
.B1(n_1544),
.B2(n_1564),
.Y(n_2384)
);

BUFx2_ASAP7_75t_SL g2385 ( 
.A(n_2149),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2031),
.Y(n_2386)
);

AO31x2_ASAP7_75t_L g2387 ( 
.A1(n_2211),
.A2(n_1932),
.A3(n_1882),
.B(n_1880),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2098),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2098),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_2139),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2257),
.B(n_1854),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2040),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_2032),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2257),
.B(n_1832),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2040),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2261),
.B(n_2186),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2024),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2031),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2024),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2261),
.B(n_2005),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2276),
.A2(n_1564),
.B1(n_1624),
.B2(n_1982),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2038),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2188),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2188),
.Y(n_2404)
);

AO31x2_ASAP7_75t_L g2405 ( 
.A1(n_2211),
.A2(n_1869),
.A3(n_2002),
.B(n_1933),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2186),
.B(n_1976),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2192),
.Y(n_2407)
);

AO31x2_ASAP7_75t_L g2408 ( 
.A1(n_2224),
.A2(n_2002),
.A3(n_1933),
.B(n_1905),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2192),
.Y(n_2409)
);

BUFx3_ASAP7_75t_L g2410 ( 
.A(n_2172),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2187),
.B(n_1976),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2187),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2197),
.B(n_1905),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2025),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2203),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_2032),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_2203),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2276),
.A2(n_2042),
.B1(n_2083),
.B2(n_2165),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2225),
.B(n_1933),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2173),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2171),
.B(n_2010),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2262),
.B(n_2283),
.Y(n_2422)
);

BUFx2_ASAP7_75t_SL g2423 ( 
.A(n_2149),
.Y(n_2423)
);

INVx3_ASAP7_75t_L g2424 ( 
.A(n_2234),
.Y(n_2424)
);

OR2x2_ASAP7_75t_L g2425 ( 
.A(n_2225),
.B(n_1819),
.Y(n_2425)
);

OR2x2_ASAP7_75t_L g2426 ( 
.A(n_2227),
.B(n_1819),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2251),
.A2(n_1864),
.B1(n_1786),
.B2(n_1906),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2173),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2171),
.B(n_1819),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2195),
.B(n_1624),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2175),
.B(n_1819),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2169),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2169),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_2205),
.B(n_1936),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2175),
.B(n_1888),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2025),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2280),
.B(n_1888),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2280),
.B(n_2252),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2167),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2139),
.Y(n_2440)
);

HB1xp67_ASAP7_75t_L g2441 ( 
.A(n_2167),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2252),
.B(n_1881),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2029),
.Y(n_2443)
);

OR2x2_ASAP7_75t_L g2444 ( 
.A(n_2227),
.B(n_1892),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_2038),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2170),
.Y(n_2446)
);

INVx2_ASAP7_75t_SL g2447 ( 
.A(n_2038),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2254),
.B(n_1881),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_2177),
.B(n_1895),
.Y(n_2449)
);

BUFx12f_ASAP7_75t_L g2450 ( 
.A(n_2278),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2029),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2254),
.B(n_1704),
.Y(n_2452)
);

AO221x2_ASAP7_75t_L g2453 ( 
.A1(n_2238),
.A2(n_1830),
.B1(n_1983),
.B2(n_1920),
.C(n_1971),
.Y(n_2453)
);

HB1xp67_ASAP7_75t_L g2454 ( 
.A(n_2147),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2030),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2030),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2124),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2124),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2177),
.B(n_1895),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2062),
.Y(n_2460)
);

INVx3_ASAP7_75t_L g2461 ( 
.A(n_2234),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2262),
.B(n_1921),
.Y(n_2462)
);

BUFx2_ASAP7_75t_L g2463 ( 
.A(n_2084),
.Y(n_2463)
);

AOI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_2276),
.A2(n_1624),
.B1(n_1760),
.B2(n_1757),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2062),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2147),
.Y(n_2466)
);

OAI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2276),
.A2(n_1907),
.B1(n_1687),
.B2(n_1745),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2084),
.B(n_1704),
.Y(n_2468)
);

OAI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2100),
.A2(n_1745),
.B1(n_1907),
.B2(n_1979),
.Y(n_2469)
);

OAI21xp5_ASAP7_75t_SL g2470 ( 
.A1(n_2134),
.A2(n_2168),
.B(n_2100),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2170),
.Y(n_2471)
);

OA21x2_ASAP7_75t_L g2472 ( 
.A1(n_2286),
.A2(n_1930),
.B(n_1914),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2084),
.B(n_1666),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2051),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2094),
.A2(n_2135),
.B1(n_2083),
.B2(n_2048),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2283),
.B(n_1909),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2064),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2243),
.B(n_1757),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2087),
.B(n_1704),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2064),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2051),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2060),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2060),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2087),
.B(n_1704),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2066),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2087),
.B(n_1666),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2066),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2263),
.B(n_1666),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2263),
.B(n_1979),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2151),
.B(n_1983),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2172),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2151),
.B(n_2009),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2074),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2074),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2135),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2077),
.Y(n_2496)
);

OR2x2_ASAP7_75t_L g2497 ( 
.A(n_2178),
.B(n_1745),
.Y(n_2497)
);

NOR2x1_ASAP7_75t_L g2498 ( 
.A(n_2094),
.B(n_1745),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2268),
.B(n_1349),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2268),
.B(n_1349),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2287),
.B(n_1163),
.Y(n_2501)
);

BUFx3_ASAP7_75t_L g2502 ( 
.A(n_2214),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2278),
.Y(n_2503)
);

BUFx2_ASAP7_75t_SL g2504 ( 
.A(n_2149),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2128),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2077),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2223),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2080),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2269),
.B(n_1099),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2080),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2088),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2269),
.B(n_2235),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2088),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2090),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2090),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2091),
.Y(n_2516)
);

INVx3_ASAP7_75t_L g2517 ( 
.A(n_2161),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2091),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_2161),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2287),
.B(n_2028),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2214),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2235),
.B(n_2237),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2132),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2132),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2237),
.B(n_2241),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2142),
.Y(n_2526)
);

OAI222xp33_ASAP7_75t_L g2527 ( 
.A1(n_2138),
.A2(n_2157),
.B1(n_2125),
.B2(n_2163),
.C1(n_2206),
.C2(n_2104),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2050),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2101),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2101),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2106),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2214),
.Y(n_2532)
);

INVxp67_ASAP7_75t_L g2533 ( 
.A(n_2092),
.Y(n_2533)
);

INVx5_ASAP7_75t_L g2534 ( 
.A(n_2206),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2241),
.B(n_2166),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2178),
.B(n_2103),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2223),
.B(n_2285),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2106),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2142),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2108),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2018),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2166),
.B(n_2267),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2108),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2103),
.B(n_2109),
.Y(n_2544)
);

INVx4_ASAP7_75t_L g2545 ( 
.A(n_2232),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2243),
.B(n_2039),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2224),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2293),
.B(n_2266),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2293),
.B(n_2266),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2392),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2300),
.Y(n_2551)
);

OR2x2_ASAP7_75t_SL g2552 ( 
.A(n_2476),
.B(n_2503),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2296),
.B(n_2266),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2288),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2296),
.B(n_2282),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2323),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2547),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2288),
.Y(n_2558)
);

INVx2_ASAP7_75t_R g2559 ( 
.A(n_2534),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2547),
.Y(n_2560)
);

INVxp67_ASAP7_75t_SL g2561 ( 
.A(n_2495),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2392),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2395),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2547),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2395),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2507),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2462),
.B(n_2102),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2444),
.B(n_2131),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2302),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2302),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_2305),
.B(n_2233),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2304),
.Y(n_2572)
);

AND2x4_ASAP7_75t_SL g2573 ( 
.A(n_2339),
.B(n_2206),
.Y(n_2573)
);

INVx5_ASAP7_75t_L g2574 ( 
.A(n_2343),
.Y(n_2574)
);

INVxp67_ASAP7_75t_SL g2575 ( 
.A(n_2495),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2289),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2289),
.Y(n_2577)
);

INVxp67_ASAP7_75t_L g2578 ( 
.A(n_2374),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2304),
.Y(n_2579)
);

OR2x2_ASAP7_75t_L g2580 ( 
.A(n_2444),
.B(n_2131),
.Y(n_2580)
);

CKINVDCx20_ASAP7_75t_R g2581 ( 
.A(n_2370),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2318),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2454),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2290),
.Y(n_2584)
);

BUFx3_ASAP7_75t_L g2585 ( 
.A(n_2305),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2388),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2290),
.Y(n_2587)
);

NOR2xp67_ASAP7_75t_SL g2588 ( 
.A(n_2343),
.B(n_2278),
.Y(n_2588)
);

AND2x4_ASAP7_75t_SL g2589 ( 
.A(n_2339),
.B(n_2206),
.Y(n_2589)
);

OAI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2354),
.A2(n_2245),
.B1(n_2206),
.B2(n_2112),
.Y(n_2590)
);

AOI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2309),
.A2(n_2094),
.B1(n_2039),
.B2(n_2217),
.Y(n_2591)
);

INVxp67_ASAP7_75t_SL g2592 ( 
.A(n_2475),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2492),
.B(n_2200),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2323),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2371),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2318),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2320),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2342),
.B(n_2039),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2320),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2324),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2324),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2316),
.A2(n_2245),
.B1(n_2079),
.B2(n_2039),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2292),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2335),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2546),
.B(n_2282),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2546),
.B(n_2282),
.Y(n_2606)
);

BUFx6f_ASAP7_75t_L g2607 ( 
.A(n_2503),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2371),
.Y(n_2608)
);

AND2x4_ASAP7_75t_L g2609 ( 
.A(n_2342),
.B(n_2212),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2335),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2546),
.B(n_2212),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2348),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2466),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2292),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2517),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2517),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2348),
.Y(n_2617)
);

HB1xp67_ASAP7_75t_L g2618 ( 
.A(n_2439),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2305),
.Y(n_2619)
);

OAI221xp5_ASAP7_75t_SL g2620 ( 
.A1(n_2475),
.A2(n_2216),
.B1(n_2213),
.B2(n_2116),
.C(n_2133),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2351),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2295),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2441),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2295),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2351),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2341),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2301),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2387),
.B(n_2109),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2366),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2366),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2546),
.B(n_2364),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2301),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2368),
.Y(n_2633)
);

INVx2_ASAP7_75t_SL g2634 ( 
.A(n_2517),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2368),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2364),
.B(n_2213),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2403),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2403),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2379),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2309),
.A2(n_2217),
.B1(n_2205),
.B2(n_2076),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2379),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2382),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2342),
.B(n_2216),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2404),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2382),
.Y(n_2645)
);

BUFx2_ASAP7_75t_L g2646 ( 
.A(n_2353),
.Y(n_2646)
);

NAND2x1p5_ASAP7_75t_L g2647 ( 
.A(n_2498),
.B(n_2093),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2381),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2388),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2389),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2387),
.B(n_2425),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2389),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2404),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2397),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2397),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2407),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2326),
.B(n_2122),
.Y(n_2657)
);

HB1xp67_ASAP7_75t_L g2658 ( 
.A(n_2505),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2399),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2490),
.B(n_2122),
.Y(n_2660)
);

INVx11_ASAP7_75t_L g2661 ( 
.A(n_2450),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2457),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2367),
.B(n_2217),
.Y(n_2663)
);

OR2x2_ASAP7_75t_L g2664 ( 
.A(n_2387),
.B(n_2114),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2457),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2407),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2517),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2399),
.Y(n_2668)
);

OR2x2_ASAP7_75t_L g2669 ( 
.A(n_2387),
.B(n_2425),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2367),
.B(n_2217),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2414),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2303),
.B(n_2299),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2303),
.B(n_2148),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2299),
.B(n_2148),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2314),
.B(n_2148),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2414),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2341),
.B(n_2232),
.Y(n_2677)
);

AOI22xp33_ASAP7_75t_L g2678 ( 
.A1(n_2375),
.A2(n_2314),
.B1(n_2365),
.B2(n_2330),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2330),
.B(n_2148),
.Y(n_2679)
);

OAI33xp33_ASAP7_75t_L g2680 ( 
.A1(n_2426),
.A2(n_2180),
.A3(n_2045),
.B1(n_2055),
.B2(n_2054),
.B3(n_2053),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2353),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2436),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2365),
.B(n_2236),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2463),
.B(n_2236),
.Y(n_2684)
);

NOR2x1_ASAP7_75t_SL g2685 ( 
.A(n_2342),
.B(n_2076),
.Y(n_2685)
);

BUFx3_ASAP7_75t_L g2686 ( 
.A(n_2341),
.Y(n_2686)
);

INVx3_ASAP7_75t_L g2687 ( 
.A(n_2519),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2436),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2460),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2519),
.Y(n_2690)
);

BUFx3_ASAP7_75t_L g2691 ( 
.A(n_2345),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2520),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2463),
.B(n_2236),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2308),
.B(n_2236),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2308),
.B(n_2158),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2342),
.B(n_2033),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2460),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2465),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2533),
.B(n_2085),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2465),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2409),
.Y(n_2701)
);

INVxp67_ASAP7_75t_SL g2702 ( 
.A(n_2498),
.Y(n_2702)
);

INVx1_ASAP7_75t_SL g2703 ( 
.A(n_2541),
.Y(n_2703)
);

OA21x2_ASAP7_75t_L g2704 ( 
.A1(n_2419),
.A2(n_2286),
.B(n_2231),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2409),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2477),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2519),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2387),
.B(n_2114),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2536),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2458),
.Y(n_2710)
);

NAND3xp33_ASAP7_75t_L g2711 ( 
.A(n_2313),
.B(n_2470),
.C(n_2418),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2298),
.B(n_2158),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2536),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2544),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2458),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2298),
.B(n_2159),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2343),
.B(n_2232),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2358),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2358),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2544),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2359),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2534),
.B(n_2033),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2359),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2361),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2443),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2361),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2387),
.B(n_2115),
.Y(n_2727)
);

INVx3_ASAP7_75t_L g2728 ( 
.A(n_2519),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2345),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2419),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2294),
.B(n_2085),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2363),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2363),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2373),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2477),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2373),
.Y(n_2736)
);

INVxp67_ASAP7_75t_L g2737 ( 
.A(n_2422),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2480),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2480),
.Y(n_2739)
);

INVx2_ASAP7_75t_SL g2740 ( 
.A(n_2376),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2443),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2426),
.B(n_2115),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2451),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2451),
.Y(n_2744)
);

BUFx2_ASAP7_75t_L g2745 ( 
.A(n_2393),
.Y(n_2745)
);

INVx2_ASAP7_75t_SL g2746 ( 
.A(n_2376),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2534),
.B(n_2052),
.Y(n_2747)
);

INVxp33_ASAP7_75t_L g2748 ( 
.A(n_2430),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2362),
.B(n_2391),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2383),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2321),
.B(n_2535),
.Y(n_2751)
);

AOI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2313),
.A2(n_2180),
.B1(n_2054),
.B2(n_2058),
.C(n_2055),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2455),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2383),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2386),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2321),
.B(n_2159),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2535),
.B(n_2267),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2386),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2455),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2337),
.B(n_2271),
.Y(n_2760)
);

OAI222xp33_ASAP7_75t_L g2761 ( 
.A1(n_2427),
.A2(n_2244),
.B1(n_2041),
.B2(n_2183),
.C1(n_2052),
.C2(n_2097),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2337),
.B(n_2271),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2456),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2398),
.Y(n_2764)
);

AOI221xp5_ASAP7_75t_L g2765 ( 
.A1(n_2470),
.A2(n_2058),
.B1(n_2053),
.B2(n_2049),
.C(n_2045),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2456),
.Y(n_2766)
);

HB1xp67_ASAP7_75t_L g2767 ( 
.A(n_2412),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2327),
.B(n_2394),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2482),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2338),
.B(n_2156),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2398),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2482),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2338),
.B(n_2156),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_L g2774 ( 
.A1(n_2453),
.A2(n_2076),
.B1(n_2047),
.B2(n_2150),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2357),
.B(n_2190),
.Y(n_2775)
);

AND2x6_ASAP7_75t_L g2776 ( 
.A(n_2503),
.B(n_2278),
.Y(n_2776)
);

HB1xp67_ASAP7_75t_L g2777 ( 
.A(n_2415),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2752),
.B(n_2355),
.Y(n_2778)
);

AND2x4_ASAP7_75t_L g2779 ( 
.A(n_2574),
.B(n_2534),
.Y(n_2779)
);

OR2x2_ASAP7_75t_L g2780 ( 
.A(n_2568),
.B(n_2291),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2550),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2574),
.B(n_2534),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2574),
.B(n_2534),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2631),
.B(n_2561),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2631),
.B(n_2575),
.Y(n_2785)
);

OR2x2_ASAP7_75t_L g2786 ( 
.A(n_2568),
.B(n_2291),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2663),
.B(n_2355),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2765),
.B(n_2344),
.Y(n_2788)
);

AOI21xp33_ASAP7_75t_L g2789 ( 
.A1(n_2711),
.A2(n_2469),
.B(n_2434),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2745),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2562),
.Y(n_2791)
);

INVxp67_ASAP7_75t_SL g2792 ( 
.A(n_2551),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2660),
.B(n_2344),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2563),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2565),
.Y(n_2795)
);

INVxp67_ASAP7_75t_SL g2796 ( 
.A(n_2648),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2663),
.B(n_2331),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2586),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2649),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2650),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2745),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2670),
.B(n_2331),
.Y(n_2802)
);

OAI21xp33_ASAP7_75t_L g2803 ( 
.A1(n_2591),
.A2(n_2774),
.B(n_2592),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2670),
.B(n_2331),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2557),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2598),
.B(n_2331),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2598),
.B(n_2424),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2652),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2598),
.B(n_2424),
.Y(n_2809)
);

OR2x2_ASAP7_75t_L g2810 ( 
.A(n_2731),
.B(n_2537),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2605),
.B(n_2606),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2715),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2692),
.B(n_2352),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2715),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2662),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2605),
.B(n_2424),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2665),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2606),
.B(n_2424),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2567),
.Y(n_2819)
);

INVx2_ASAP7_75t_SL g2820 ( 
.A(n_2661),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2593),
.B(n_2578),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2768),
.B(n_2749),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2672),
.B(n_2461),
.Y(n_2823)
);

CKINVDCx5p33_ASAP7_75t_R g2824 ( 
.A(n_2581),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2710),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2554),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2574),
.B(n_2343),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2672),
.B(n_2461),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2554),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2611),
.B(n_2461),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2611),
.B(n_2461),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2557),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2558),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2747),
.B(n_2542),
.Y(n_2834)
);

NAND2x1_ASAP7_75t_L g2835 ( 
.A(n_2595),
.B(n_2393),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2558),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2646),
.A2(n_2453),
.B1(n_2545),
.B2(n_2423),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2560),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2747),
.B(n_2542),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2747),
.B(n_2548),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2580),
.B(n_2116),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2576),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2560),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2737),
.B(n_2657),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2595),
.Y(n_2845)
);

HB1xp67_ASAP7_75t_L g2846 ( 
.A(n_2658),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2548),
.B(n_2357),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2564),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2549),
.B(n_2360),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2678),
.B(n_2352),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2576),
.Y(n_2851)
);

AND2x4_ASAP7_75t_L g2852 ( 
.A(n_2574),
.B(n_2545),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2577),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2549),
.B(n_2360),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2699),
.B(n_2522),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2577),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2582),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2556),
.B(n_2594),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2553),
.B(n_2522),
.Y(n_2859)
);

INVx5_ASAP7_75t_L g2860 ( 
.A(n_2776),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2564),
.Y(n_2861)
);

AOI22xp33_ASAP7_75t_L g2862 ( 
.A1(n_2640),
.A2(n_2602),
.B1(n_2453),
.B2(n_2646),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2628),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2553),
.B(n_2525),
.Y(n_2864)
);

OR2x2_ASAP7_75t_L g2865 ( 
.A(n_2580),
.B(n_2307),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2555),
.B(n_2525),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2628),
.Y(n_2867)
);

OR2x2_ASAP7_75t_L g2868 ( 
.A(n_2709),
.B(n_2307),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2555),
.B(n_2317),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2683),
.B(n_2317),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2683),
.B(n_2468),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2566),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2582),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2596),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2581),
.Y(n_2875)
);

BUFx2_ASAP7_75t_L g2876 ( 
.A(n_2585),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2596),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2684),
.B(n_2468),
.Y(n_2878)
);

NOR2xp33_ASAP7_75t_L g2879 ( 
.A(n_2585),
.B(n_2345),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2619),
.B(n_2421),
.Y(n_2880)
);

BUFx2_ASAP7_75t_L g2881 ( 
.A(n_2619),
.Y(n_2881)
);

AND2x4_ASAP7_75t_L g2882 ( 
.A(n_2556),
.B(n_2545),
.Y(n_2882)
);

INVx2_ASAP7_75t_SL g2883 ( 
.A(n_2661),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2597),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2684),
.B(n_2473),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2681),
.A2(n_2453),
.B1(n_2545),
.B2(n_2423),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2693),
.B(n_2473),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2626),
.B(n_2421),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2693),
.B(n_2674),
.Y(n_2889)
);

BUFx2_ASAP7_75t_L g2890 ( 
.A(n_2626),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2664),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2686),
.B(n_2322),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2664),
.Y(n_2893)
);

INVx2_ASAP7_75t_SL g2894 ( 
.A(n_2556),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2597),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2599),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2599),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2674),
.B(n_2675),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2600),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2686),
.B(n_2319),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2600),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2601),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2675),
.B(n_2479),
.Y(n_2903)
);

INVx3_ASAP7_75t_L g2904 ( 
.A(n_2595),
.Y(n_2904)
);

BUFx2_ASAP7_75t_L g2905 ( 
.A(n_2691),
.Y(n_2905)
);

OAI21xp5_ASAP7_75t_SL g2906 ( 
.A1(n_2681),
.A2(n_2340),
.B(n_2527),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2601),
.Y(n_2907)
);

INVx2_ASAP7_75t_SL g2908 ( 
.A(n_2594),
.Y(n_2908)
);

NAND2x1p5_ASAP7_75t_L g2909 ( 
.A(n_2588),
.B(n_2376),
.Y(n_2909)
);

NAND2x1_ASAP7_75t_L g2910 ( 
.A(n_2608),
.B(n_2594),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2604),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2708),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2691),
.B(n_2319),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2729),
.B(n_2310),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2583),
.B(n_2350),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2604),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_2608),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2613),
.B(n_2350),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2679),
.B(n_2479),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2729),
.B(n_2310),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2708),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2610),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2727),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2727),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2610),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2612),
.Y(n_2926)
);

OR2x2_ASAP7_75t_L g2927 ( 
.A(n_2709),
.B(n_2429),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2612),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2679),
.B(n_2484),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2751),
.Y(n_2930)
);

HB1xp67_ASAP7_75t_L g2931 ( 
.A(n_2618),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2571),
.Y(n_2932)
);

AND2x4_ASAP7_75t_L g2933 ( 
.A(n_2608),
.B(n_2410),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2751),
.Y(n_2934)
);

AOI22xp33_ASAP7_75t_L g2935 ( 
.A1(n_2590),
.A2(n_2047),
.B1(n_2086),
.B2(n_2347),
.Y(n_2935)
);

NAND4xp25_ASAP7_75t_L g2936 ( 
.A(n_2620),
.B(n_2401),
.C(n_2384),
.D(n_2377),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2673),
.B(n_2775),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2617),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2617),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2621),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2748),
.B(n_2435),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2573),
.B(n_2410),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2673),
.B(n_2484),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2775),
.B(n_2486),
.Y(n_2944)
);

AND2x4_ASAP7_75t_L g2945 ( 
.A(n_2573),
.B(n_2589),
.Y(n_2945)
);

AND2x4_ASAP7_75t_L g2946 ( 
.A(n_2589),
.B(n_2410),
.Y(n_2946)
);

OR2x2_ASAP7_75t_L g2947 ( 
.A(n_2623),
.B(n_2198),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2694),
.B(n_2636),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2694),
.B(n_2486),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2621),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2569),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2636),
.B(n_2385),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2609),
.B(n_2385),
.Y(n_2953)
);

INVxp67_ASAP7_75t_L g2954 ( 
.A(n_2767),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2609),
.B(n_2643),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2569),
.Y(n_2956)
);

HB1xp67_ASAP7_75t_L g2957 ( 
.A(n_2777),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2625),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2570),
.Y(n_2959)
);

AND2x2_ASAP7_75t_SL g2960 ( 
.A(n_2677),
.B(n_2356),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2740),
.B(n_2435),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2625),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2570),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_SL g2964 ( 
.A(n_2607),
.B(n_2503),
.Y(n_2964)
);

AND2x4_ASAP7_75t_L g2965 ( 
.A(n_2696),
.B(n_2491),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2572),
.Y(n_2966)
);

NOR2x1p5_ASAP7_75t_L g2967 ( 
.A(n_2702),
.B(n_2347),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2629),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2629),
.Y(n_2969)
);

INVxp67_ASAP7_75t_L g2970 ( 
.A(n_2740),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2609),
.B(n_2504),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2630),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2630),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2746),
.B(n_2297),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2633),
.Y(n_2975)
);

OR2x6_ASAP7_75t_L g2976 ( 
.A(n_2717),
.B(n_2504),
.Y(n_2976)
);

INVxp67_ASAP7_75t_SL g2977 ( 
.A(n_2790),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2952),
.B(n_2760),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2860),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2812),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2819),
.B(n_2746),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2814),
.Y(n_2982)
);

OAI322xp33_ASAP7_75t_L g2983 ( 
.A1(n_2778),
.A2(n_2669),
.A3(n_2651),
.B1(n_2730),
.B2(n_2647),
.C1(n_2713),
.C2(n_2720),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2952),
.B(n_2760),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2826),
.Y(n_2985)
);

AOI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2862),
.A2(n_2047),
.B1(n_2043),
.B2(n_2021),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2784),
.Y(n_2987)
);

AOI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2862),
.A2(n_2043),
.B1(n_2021),
.B2(n_2093),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2784),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2785),
.Y(n_2990)
);

AOI221xp5_ASAP7_75t_L g2991 ( 
.A1(n_2803),
.A2(n_2761),
.B1(n_2680),
.B2(n_2730),
.C(n_2714),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2785),
.B(n_2953),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2876),
.B(n_2757),
.Y(n_2993)
);

OA21x2_ASAP7_75t_L g2994 ( 
.A1(n_2964),
.A2(n_2579),
.B(n_2572),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2953),
.B(n_2762),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2829),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2833),
.Y(n_2997)
);

HB1xp67_ASAP7_75t_L g2998 ( 
.A(n_2846),
.Y(n_2998)
);

OAI211xp5_ASAP7_75t_SL g2999 ( 
.A1(n_2789),
.A2(n_2703),
.B(n_2651),
.C(n_2669),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2971),
.B(n_2762),
.Y(n_3000)
);

AO21x2_ASAP7_75t_L g3001 ( 
.A1(n_2964),
.A2(n_2685),
.B(n_2552),
.Y(n_3001)
);

OAI22xp5_ASAP7_75t_SL g3002 ( 
.A1(n_2837),
.A2(n_2552),
.B1(n_2347),
.B2(n_2440),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2813),
.B(n_2713),
.Y(n_3003)
);

OAI31xp33_ASAP7_75t_L g3004 ( 
.A1(n_2906),
.A2(n_2647),
.A3(n_2696),
.B(n_2722),
.Y(n_3004)
);

BUFx2_ASAP7_75t_L g3005 ( 
.A(n_2976),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2847),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2836),
.Y(n_3007)
);

AO21x2_ASAP7_75t_L g3008 ( 
.A1(n_2790),
.A2(n_2685),
.B(n_2635),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2842),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2847),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2851),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2853),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2849),
.Y(n_3013)
);

OR2x2_ASAP7_75t_L g3014 ( 
.A(n_2793),
.B(n_2714),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2856),
.Y(n_3015)
);

INVx2_ASAP7_75t_SL g3016 ( 
.A(n_2875),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2857),
.Y(n_3017)
);

HB1xp67_ASAP7_75t_L g3018 ( 
.A(n_2872),
.Y(n_3018)
);

AOI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2850),
.A2(n_2021),
.B1(n_2472),
.B2(n_2086),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2873),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2874),
.Y(n_3021)
);

AND4x1_ASAP7_75t_L g3022 ( 
.A(n_2886),
.B(n_2588),
.C(n_2152),
.D(n_2464),
.Y(n_3022)
);

AND2x4_ASAP7_75t_L g3023 ( 
.A(n_2967),
.B(n_2696),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_R g3024 ( 
.A(n_2820),
.B(n_2390),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2971),
.B(n_2757),
.Y(n_3025)
);

OAI31xp33_ASAP7_75t_SL g3026 ( 
.A1(n_2787),
.A2(n_2722),
.A3(n_2467),
.B(n_2643),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2877),
.Y(n_3027)
);

AOI22xp5_ASAP7_75t_L g3028 ( 
.A1(n_2788),
.A2(n_2776),
.B1(n_2643),
.B2(n_2450),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2884),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2801),
.Y(n_3030)
);

OAI221xp5_ASAP7_75t_L g3031 ( 
.A1(n_2935),
.A2(n_2647),
.B1(n_2380),
.B2(n_2528),
.C(n_2503),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2935),
.A2(n_2722),
.B(n_2607),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2976),
.A2(n_2607),
.B1(n_2528),
.B2(n_2502),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2881),
.B(n_2890),
.Y(n_3034)
);

AOI221xp5_ASAP7_75t_L g3035 ( 
.A1(n_2954),
.A2(n_2720),
.B1(n_2706),
.B2(n_2668),
.C(n_2700),
.Y(n_3035)
);

AOI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_2960),
.A2(n_2776),
.B1(n_2607),
.B2(n_2442),
.Y(n_3036)
);

A2O1A1Ixp33_ASAP7_75t_L g3037 ( 
.A1(n_2960),
.A2(n_2044),
.B(n_2502),
.C(n_2491),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2895),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2896),
.Y(n_3039)
);

AOI211xp5_ASAP7_75t_L g3040 ( 
.A1(n_2936),
.A2(n_2607),
.B(n_2502),
.C(n_2521),
.Y(n_3040)
);

HB1xp67_ASAP7_75t_L g3041 ( 
.A(n_2931),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2849),
.Y(n_3042)
);

OA21x2_ASAP7_75t_L g3043 ( 
.A1(n_2801),
.A2(n_2579),
.B(n_2584),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2844),
.B(n_2198),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2897),
.Y(n_3045)
);

INVx4_ASAP7_75t_SL g3046 ( 
.A(n_2820),
.Y(n_3046)
);

OR2x2_ASAP7_75t_L g3047 ( 
.A(n_2810),
.B(n_2821),
.Y(n_3047)
);

AND2x4_ASAP7_75t_L g3048 ( 
.A(n_2976),
.B(n_2776),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2840),
.B(n_2770),
.Y(n_3049)
);

INVx2_ASAP7_75t_SL g3050 ( 
.A(n_2875),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2932),
.A2(n_2472),
.B1(n_2086),
.B2(n_2559),
.Y(n_3051)
);

BUFx3_ASAP7_75t_L g3052 ( 
.A(n_2905),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2899),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2901),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2854),
.Y(n_3055)
);

OA21x2_ASAP7_75t_L g3056 ( 
.A1(n_2970),
.A2(n_2587),
.B(n_2584),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2902),
.Y(n_3057)
);

AOI221xp5_ASAP7_75t_L g3058 ( 
.A1(n_2792),
.A2(n_2659),
.B1(n_2698),
.B2(n_2697),
.C(n_2655),
.Y(n_3058)
);

NOR2x1_ASAP7_75t_L g3059 ( 
.A(n_2932),
.B(n_2615),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2907),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2796),
.B(n_2695),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_L g3062 ( 
.A1(n_2787),
.A2(n_2472),
.B1(n_2086),
.B2(n_2559),
.Y(n_3062)
);

HB1xp67_ASAP7_75t_L g3063 ( 
.A(n_2957),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_2883),
.A2(n_2472),
.B1(n_2559),
.B2(n_2776),
.Y(n_3064)
);

OAI221xp5_ASAP7_75t_L g3065 ( 
.A1(n_2976),
.A2(n_2491),
.B1(n_2521),
.B2(n_2532),
.C(n_2707),
.Y(n_3065)
);

BUFx2_ASAP7_75t_L g3066 ( 
.A(n_2945),
.Y(n_3066)
);

BUFx2_ASAP7_75t_L g3067 ( 
.A(n_2945),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2911),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2916),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2922),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2854),
.Y(n_3071)
);

NOR3xp33_ASAP7_75t_L g3072 ( 
.A(n_2879),
.B(n_2501),
.C(n_2044),
.Y(n_3072)
);

AOI221xp5_ASAP7_75t_L g3073 ( 
.A1(n_2822),
.A2(n_2654),
.B1(n_2688),
.B2(n_2689),
.C(n_2738),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2898),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_SL g3075 ( 
.A1(n_2909),
.A2(n_2776),
.B1(n_2150),
.B2(n_2523),
.Y(n_3075)
);

HB1xp67_ASAP7_75t_L g3076 ( 
.A(n_2925),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2898),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2926),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2928),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2889),
.Y(n_3080)
);

INVx1_ASAP7_75t_SL g3081 ( 
.A(n_2824),
.Y(n_3081)
);

NAND3xp33_ASAP7_75t_L g3082 ( 
.A(n_2815),
.B(n_2431),
.C(n_2429),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2938),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2892),
.B(n_2879),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2939),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2940),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2883),
.B(n_2763),
.Y(n_3087)
);

OAI33xp33_ASAP7_75t_L g3088 ( 
.A1(n_2817),
.A2(n_2738),
.A3(n_2671),
.B1(n_2676),
.B2(n_2682),
.B3(n_2633),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2950),
.Y(n_3089)
);

BUFx6f_ASAP7_75t_L g3090 ( 
.A(n_2827),
.Y(n_3090)
);

OA21x2_ASAP7_75t_L g3091 ( 
.A1(n_2882),
.A2(n_2852),
.B(n_2827),
.Y(n_3091)
);

HB1xp67_ASAP7_75t_L g3092 ( 
.A(n_2958),
.Y(n_3092)
);

OR2x6_ASAP7_75t_L g3093 ( 
.A(n_2827),
.B(n_2278),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2860),
.Y(n_3094)
);

BUFx3_ASAP7_75t_L g3095 ( 
.A(n_2824),
.Y(n_3095)
);

OAI221xp5_ASAP7_75t_L g3096 ( 
.A1(n_2909),
.A2(n_2532),
.B1(n_2521),
.B2(n_2690),
.C(n_2707),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2962),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2889),
.Y(n_3098)
);

INVx1_ASAP7_75t_SL g3099 ( 
.A(n_2945),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2968),
.Y(n_3100)
);

AOI211xp5_ASAP7_75t_L g3101 ( 
.A1(n_2779),
.A2(n_2532),
.B(n_2431),
.C(n_2448),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2840),
.B(n_2770),
.Y(n_3102)
);

BUFx2_ASAP7_75t_L g3103 ( 
.A(n_2852),
.Y(n_3103)
);

OR2x2_ASAP7_75t_L g3104 ( 
.A(n_2915),
.B(n_2742),
.Y(n_3104)
);

HB1xp67_ASAP7_75t_L g3105 ( 
.A(n_2969),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2972),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2973),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2975),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_2825),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2937),
.B(n_2834),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2880),
.B(n_2695),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2781),
.Y(n_3112)
);

OR2x2_ASAP7_75t_L g3113 ( 
.A(n_2918),
.B(n_2742),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2791),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2794),
.Y(n_3115)
);

AOI221xp5_ASAP7_75t_L g3116 ( 
.A1(n_2930),
.A2(n_2739),
.B1(n_2682),
.B2(n_2676),
.C(n_2635),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2795),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2798),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2937),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2888),
.B(n_2712),
.Y(n_3120)
);

BUFx3_ASAP7_75t_L g3121 ( 
.A(n_2852),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2859),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2859),
.Y(n_3123)
);

INVxp67_ASAP7_75t_L g3124 ( 
.A(n_2799),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2864),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2834),
.B(n_2773),
.Y(n_3126)
);

AOI22xp33_ASAP7_75t_L g3127 ( 
.A1(n_2941),
.A2(n_2776),
.B1(n_2509),
.B2(n_2150),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2900),
.B(n_2712),
.Y(n_3128)
);

INVx3_ASAP7_75t_L g3129 ( 
.A(n_2860),
.Y(n_3129)
);

NAND3xp33_ASAP7_75t_L g3130 ( 
.A(n_2860),
.B(n_2782),
.C(n_2779),
.Y(n_3130)
);

INVx4_ASAP7_75t_L g3131 ( 
.A(n_2860),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2882),
.Y(n_3132)
);

AOI22xp5_ASAP7_75t_L g3133 ( 
.A1(n_2942),
.A2(n_2442),
.B1(n_2448),
.B2(n_2437),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2800),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2808),
.Y(n_3135)
);

NOR3xp33_ASAP7_75t_SL g3136 ( 
.A(n_2913),
.B(n_2218),
.C(n_2769),
.Y(n_3136)
);

INVx2_ASAP7_75t_SL g3137 ( 
.A(n_2942),
.Y(n_3137)
);

INVx4_ASAP7_75t_L g3138 ( 
.A(n_2779),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2839),
.B(n_2773),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2951),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2944),
.B(n_2914),
.Y(n_3141)
);

AOI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_2942),
.A2(n_2437),
.B1(n_2509),
.B2(n_2478),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2839),
.B(n_2716),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2951),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2956),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2956),
.Y(n_3146)
);

OR2x2_ASAP7_75t_L g3147 ( 
.A(n_2987),
.B(n_2930),
.Y(n_3147)
);

BUFx2_ASAP7_75t_L g3148 ( 
.A(n_3024),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2992),
.B(n_2946),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_3016),
.B(n_2948),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2998),
.Y(n_3151)
);

OR2x2_ASAP7_75t_L g3152 ( 
.A(n_2987),
.B(n_2934),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2998),
.Y(n_3153)
);

NOR2xp67_ASAP7_75t_L g3154 ( 
.A(n_3131),
.B(n_2946),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_3059),
.B(n_3052),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3018),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3018),
.Y(n_3157)
);

BUFx3_ASAP7_75t_L g3158 ( 
.A(n_3095),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3041),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_3050),
.B(n_2948),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3041),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3063),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_3095),
.B(n_2946),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3063),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_3091),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3076),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3076),
.Y(n_3167)
);

INVxp67_ASAP7_75t_SL g3168 ( 
.A(n_3052),
.Y(n_3168)
);

AND3x2_ASAP7_75t_L g3169 ( 
.A(n_3040),
.B(n_2783),
.C(n_2782),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_3132),
.B(n_2882),
.Y(n_3170)
);

OR2x2_ASAP7_75t_L g3171 ( 
.A(n_2989),
.B(n_2934),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3092),
.Y(n_3172)
);

OR2x2_ASAP7_75t_L g3173 ( 
.A(n_2989),
.B(n_2780),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_3091),
.Y(n_3174)
);

OR2x2_ASAP7_75t_L g3175 ( 
.A(n_2990),
.B(n_2780),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_3066),
.B(n_2944),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_3067),
.B(n_2955),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3110),
.B(n_2955),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3092),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3105),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2995),
.B(n_2933),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3099),
.B(n_2903),
.Y(n_3182)
);

AND2x2_ASAP7_75t_L g3183 ( 
.A(n_3000),
.B(n_2933),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_2978),
.B(n_2933),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_3091),
.Y(n_3185)
);

OR2x2_ASAP7_75t_L g3186 ( 
.A(n_2990),
.B(n_3061),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3087),
.B(n_2903),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3105),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_2984),
.B(n_2965),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2994),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_3087),
.B(n_2919),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2977),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2977),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_3132),
.B(n_2782),
.Y(n_3194)
);

OR2x2_ASAP7_75t_L g3195 ( 
.A(n_3006),
.B(n_2786),
.Y(n_3195)
);

HB1xp67_ASAP7_75t_L g3196 ( 
.A(n_3030),
.Y(n_3196)
);

INVx1_ASAP7_75t_SL g3197 ( 
.A(n_3024),
.Y(n_3197)
);

NAND2x1_ASAP7_75t_L g3198 ( 
.A(n_3048),
.B(n_2845),
.Y(n_3198)
);

INVxp33_ASAP7_75t_L g3199 ( 
.A(n_3002),
.Y(n_3199)
);

AOI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_2999),
.A2(n_2783),
.B1(n_2965),
.B2(n_2920),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3030),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_3025),
.B(n_2919),
.Y(n_3202)
);

INVx2_ASAP7_75t_SL g3203 ( 
.A(n_3090),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2994),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3034),
.B(n_2929),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3109),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3109),
.B(n_3081),
.Y(n_3207)
);

HB1xp67_ASAP7_75t_L g3208 ( 
.A(n_3006),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2980),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3137),
.B(n_3049),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3103),
.B(n_2929),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_3102),
.B(n_2943),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3084),
.B(n_2869),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_3022),
.B(n_2783),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_3023),
.B(n_3074),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2994),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2982),
.Y(n_3217)
);

BUFx6f_ASAP7_75t_SL g3218 ( 
.A(n_3048),
.Y(n_3218)
);

NOR2xp67_ASAP7_75t_L g3219 ( 
.A(n_3131),
.B(n_2965),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2985),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2996),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3023),
.B(n_2943),
.Y(n_3222)
);

INVx2_ASAP7_75t_SL g3223 ( 
.A(n_3090),
.Y(n_3223)
);

HB1xp67_ASAP7_75t_L g3224 ( 
.A(n_3010),
.Y(n_3224)
);

OR2x2_ASAP7_75t_L g3225 ( 
.A(n_3010),
.B(n_2786),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2997),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_3004),
.B(n_2858),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3007),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3023),
.B(n_2949),
.Y(n_3229)
);

OR2x2_ASAP7_75t_L g3230 ( 
.A(n_3013),
.B(n_2865),
.Y(n_3230)
);

NAND2x1_ASAP7_75t_L g3231 ( 
.A(n_2979),
.B(n_2845),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3009),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_3074),
.B(n_2949),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2981),
.B(n_2869),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3043),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_3126),
.B(n_2811),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3139),
.B(n_2811),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_3121),
.B(n_3138),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3047),
.B(n_2871),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2993),
.B(n_2871),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3011),
.Y(n_3241)
);

INVx2_ASAP7_75t_SL g3242 ( 
.A(n_3090),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3143),
.B(n_2806),
.Y(n_3243)
);

AND2x4_ASAP7_75t_L g3244 ( 
.A(n_3121),
.B(n_3138),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3077),
.B(n_2974),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_3043),
.Y(n_3246)
);

OR2x2_ASAP7_75t_L g3247 ( 
.A(n_3013),
.B(n_2865),
.Y(n_3247)
);

OR2x2_ASAP7_75t_L g3248 ( 
.A(n_3042),
.B(n_2841),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3005),
.B(n_2806),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3012),
.Y(n_3250)
);

OR2x2_ASAP7_75t_L g3251 ( 
.A(n_3042),
.B(n_2855),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3077),
.B(n_2870),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3043),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3015),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3017),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3080),
.B(n_2870),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3020),
.Y(n_3257)
);

AND2x4_ASAP7_75t_L g3258 ( 
.A(n_3130),
.B(n_2858),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3080),
.B(n_2864),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3093),
.B(n_2807),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3021),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3027),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3008),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3029),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3098),
.B(n_2878),
.Y(n_3265)
);

AOI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_2986),
.A2(n_2963),
.B1(n_2966),
.B2(n_2959),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3098),
.B(n_2878),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3055),
.B(n_2885),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3008),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3055),
.B(n_2866),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3071),
.B(n_2885),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_3071),
.B(n_3141),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3038),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_3056),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3056),
.Y(n_3275)
);

INVxp67_ASAP7_75t_L g3276 ( 
.A(n_3090),
.Y(n_3276)
);

BUFx2_ASAP7_75t_L g3277 ( 
.A(n_3093),
.Y(n_3277)
);

OR2x2_ASAP7_75t_L g3278 ( 
.A(n_3128),
.B(n_2868),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3039),
.Y(n_3279)
);

OR2x2_ASAP7_75t_L g3280 ( 
.A(n_3111),
.B(n_2868),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3119),
.B(n_2866),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3045),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3053),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3093),
.B(n_2807),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3054),
.Y(n_3285)
);

INVx2_ASAP7_75t_SL g3286 ( 
.A(n_2979),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3119),
.B(n_2887),
.Y(n_3287)
);

INVx1_ASAP7_75t_SL g3288 ( 
.A(n_3046),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3057),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3124),
.B(n_2887),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3046),
.B(n_2809),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3026),
.B(n_2809),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3046),
.B(n_2797),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3124),
.B(n_2961),
.Y(n_3294)
);

INVxp33_ASAP7_75t_L g3295 ( 
.A(n_3036),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3060),
.Y(n_3296)
);

OR2x2_ASAP7_75t_L g3297 ( 
.A(n_3120),
.B(n_2947),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3068),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3122),
.B(n_3123),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3056),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3136),
.B(n_2823),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3069),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_3001),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3070),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3122),
.B(n_2797),
.Y(n_3305)
);

AOI32xp33_ASAP7_75t_L g3306 ( 
.A1(n_3199),
.A2(n_2991),
.A3(n_2986),
.B1(n_3075),
.B2(n_3031),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_3148),
.B(n_3028),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3196),
.Y(n_3308)
);

OAI21xp33_ASAP7_75t_L g3309 ( 
.A1(n_3295),
.A2(n_2988),
.B(n_3019),
.Y(n_3309)
);

OR2x2_ASAP7_75t_L g3310 ( 
.A(n_3207),
.B(n_3003),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3168),
.B(n_3112),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3168),
.B(n_3114),
.Y(n_3312)
);

OR2x2_ASAP7_75t_L g3313 ( 
.A(n_3213),
.B(n_3123),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_L g3314 ( 
.A(n_3197),
.B(n_3096),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3155),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3199),
.A2(n_3136),
.B1(n_2988),
.B2(n_3037),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3276),
.B(n_3115),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_3177),
.B(n_3125),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3196),
.Y(n_3319)
);

NOR2x1_ASAP7_75t_R g3320 ( 
.A(n_3158),
.B(n_3094),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_3231),
.Y(n_3321)
);

INVx1_ASAP7_75t_SL g3322 ( 
.A(n_3158),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3155),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3208),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3276),
.B(n_3117),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3208),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3224),
.Y(n_3327)
);

INVx4_ASAP7_75t_L g3328 ( 
.A(n_3238),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3224),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3192),
.Y(n_3330)
);

A2O1A1Ixp33_ASAP7_75t_L g3331 ( 
.A1(n_3214),
.A2(n_3037),
.B(n_3032),
.C(n_3075),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3177),
.B(n_3125),
.Y(n_3332)
);

HB1xp67_ASAP7_75t_L g3333 ( 
.A(n_3165),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3193),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3176),
.B(n_3133),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3149),
.B(n_3142),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3203),
.B(n_3118),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3293),
.B(n_3001),
.Y(n_3338)
);

NAND2x1p5_ASAP7_75t_L g3339 ( 
.A(n_3155),
.B(n_3094),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3165),
.Y(n_3340)
);

INVxp67_ASAP7_75t_SL g3341 ( 
.A(n_3274),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3201),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3291),
.B(n_3129),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_3174),
.Y(n_3344)
);

INVx2_ASAP7_75t_SL g3345 ( 
.A(n_3238),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3206),
.Y(n_3346)
);

AND2x4_ASAP7_75t_L g3347 ( 
.A(n_3219),
.B(n_3129),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3189),
.B(n_2802),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3189),
.B(n_2802),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3203),
.B(n_3223),
.Y(n_3350)
);

NOR3xp33_ASAP7_75t_L g3351 ( 
.A(n_3214),
.B(n_2983),
.C(n_3088),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3223),
.B(n_3134),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3181),
.B(n_2804),
.Y(n_3353)
);

HB1xp67_ASAP7_75t_L g3354 ( 
.A(n_3174),
.Y(n_3354)
);

OR2x2_ASAP7_75t_L g3355 ( 
.A(n_3239),
.B(n_3014),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3242),
.B(n_3135),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3185),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_3163),
.B(n_3065),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3242),
.B(n_3035),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3181),
.B(n_3101),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3151),
.Y(n_3361)
);

OR2x2_ASAP7_75t_L g3362 ( 
.A(n_3182),
.B(n_3044),
.Y(n_3362)
);

HB1xp67_ASAP7_75t_L g3363 ( 
.A(n_3185),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3183),
.B(n_2804),
.Y(n_3364)
);

BUFx2_ASAP7_75t_L g3365 ( 
.A(n_3238),
.Y(n_3365)
);

NOR3xp33_ASAP7_75t_L g3366 ( 
.A(n_3153),
.B(n_3088),
.C(n_3033),
.Y(n_3366)
);

INVx3_ASAP7_75t_SL g3367 ( 
.A(n_3288),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3156),
.Y(n_3368)
);

INVxp67_ASAP7_75t_L g3369 ( 
.A(n_3163),
.Y(n_3369)
);

OR2x2_ASAP7_75t_L g3370 ( 
.A(n_3290),
.B(n_3104),
.Y(n_3370)
);

INVxp67_ASAP7_75t_SL g3371 ( 
.A(n_3274),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3157),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3159),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3161),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3183),
.B(n_3184),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3162),
.Y(n_3376)
);

AOI322xp5_ASAP7_75t_L g3377 ( 
.A1(n_3200),
.A2(n_3058),
.A3(n_3019),
.B1(n_3127),
.B2(n_3073),
.C1(n_3116),
.C2(n_3064),
.Y(n_3377)
);

AOI21xp5_ASAP7_75t_L g3378 ( 
.A1(n_3227),
.A2(n_3127),
.B(n_3064),
.Y(n_3378)
);

AOI211xp5_ASAP7_75t_L g3379 ( 
.A1(n_3295),
.A2(n_3072),
.B(n_3079),
.C(n_3078),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3184),
.B(n_2823),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3164),
.B(n_3150),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3160),
.B(n_3083),
.Y(n_3382)
);

OR2x2_ASAP7_75t_L g3383 ( 
.A(n_3287),
.B(n_3113),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3166),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3167),
.Y(n_3385)
);

OR2x2_ASAP7_75t_L g3386 ( 
.A(n_3211),
.B(n_3085),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3210),
.B(n_3086),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3172),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_3244),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3240),
.B(n_3089),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3179),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_3252),
.B(n_3097),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3180),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3222),
.B(n_2828),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_3229),
.B(n_2828),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3188),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3244),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3299),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3147),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3249),
.B(n_3100),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3244),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3190),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3190),
.Y(n_3403)
);

INVx3_ASAP7_75t_L g3404 ( 
.A(n_3170),
.Y(n_3404)
);

BUFx2_ASAP7_75t_L g3405 ( 
.A(n_3170),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3152),
.Y(n_3406)
);

INVxp67_ASAP7_75t_L g3407 ( 
.A(n_3286),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3171),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3249),
.B(n_3215),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3205),
.B(n_3106),
.Y(n_3410)
);

OR2x2_ASAP7_75t_L g3411 ( 
.A(n_3256),
.B(n_3107),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3204),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3178),
.B(n_3108),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3178),
.B(n_2858),
.Y(n_3414)
);

BUFx2_ASAP7_75t_L g3415 ( 
.A(n_3170),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3209),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3217),
.Y(n_3417)
);

OR2x2_ASAP7_75t_L g3418 ( 
.A(n_3272),
.B(n_3140),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3220),
.Y(n_3419)
);

HB1xp67_ASAP7_75t_L g3420 ( 
.A(n_3204),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3187),
.B(n_3072),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3191),
.B(n_3144),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3221),
.Y(n_3423)
);

NOR2xp33_ASAP7_75t_L g3424 ( 
.A(n_3218),
.B(n_2835),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3216),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3216),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3226),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3292),
.B(n_2816),
.Y(n_3428)
);

INVx2_ASAP7_75t_SL g3429 ( 
.A(n_3198),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3236),
.B(n_3145),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3292),
.B(n_2816),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3228),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3232),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3258),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3236),
.B(n_2818),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3237),
.B(n_2818),
.Y(n_3436)
);

HB1xp67_ASAP7_75t_L g3437 ( 
.A(n_3275),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3241),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_3237),
.B(n_2830),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3250),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3254),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3265),
.B(n_3146),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_3322),
.B(n_3218),
.Y(n_3443)
);

INVx1_ASAP7_75t_SL g3444 ( 
.A(n_3367),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3375),
.B(n_3258),
.Y(n_3445)
);

NAND3xp33_ASAP7_75t_SL g3446 ( 
.A(n_3351),
.B(n_3306),
.C(n_3378),
.Y(n_3446)
);

OR2x2_ASAP7_75t_L g3447 ( 
.A(n_3409),
.B(n_3186),
.Y(n_3447)
);

INVx2_ASAP7_75t_SL g3448 ( 
.A(n_3404),
.Y(n_3448)
);

INVxp67_ASAP7_75t_L g3449 ( 
.A(n_3320),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3367),
.B(n_3277),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3369),
.B(n_3258),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3333),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3333),
.Y(n_3453)
);

HB1xp67_ASAP7_75t_L g3454 ( 
.A(n_3405),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3354),
.Y(n_3455)
);

OR2x2_ASAP7_75t_L g3456 ( 
.A(n_3310),
.B(n_3234),
.Y(n_3456)
);

NAND2xp33_ASAP7_75t_R g3457 ( 
.A(n_3365),
.B(n_3169),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3354),
.Y(n_3458)
);

AND2x4_ASAP7_75t_L g3459 ( 
.A(n_3404),
.B(n_3154),
.Y(n_3459)
);

NOR2x1_ASAP7_75t_R g3460 ( 
.A(n_3328),
.B(n_3227),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3363),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3363),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3369),
.B(n_3194),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3437),
.Y(n_3464)
);

NAND4xp25_ASAP7_75t_L g3465 ( 
.A(n_3351),
.B(n_3200),
.C(n_3266),
.D(n_3303),
.Y(n_3465)
);

OAI21xp33_ASAP7_75t_L g3466 ( 
.A1(n_3309),
.A2(n_3245),
.B(n_3294),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3389),
.B(n_3267),
.Y(n_3467)
);

AND2x4_ASAP7_75t_L g3468 ( 
.A(n_3404),
.B(n_3194),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3437),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3318),
.B(n_3202),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3318),
.B(n_3332),
.Y(n_3471)
);

OR2x2_ASAP7_75t_L g3472 ( 
.A(n_3400),
.B(n_3297),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3414),
.B(n_3212),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3339),
.Y(n_3474)
);

OR2x2_ASAP7_75t_L g3475 ( 
.A(n_3381),
.B(n_3259),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3339),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3420),
.Y(n_3477)
);

OR2x2_ASAP7_75t_L g3478 ( 
.A(n_3398),
.B(n_3281),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3415),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3414),
.B(n_3194),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3328),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3360),
.B(n_3260),
.Y(n_3482)
);

AND4x1_ASAP7_75t_L g3483 ( 
.A(n_3314),
.B(n_3266),
.C(n_3284),
.D(n_3260),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3308),
.B(n_3255),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3420),
.Y(n_3485)
);

HB1xp67_ASAP7_75t_L g3486 ( 
.A(n_3345),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3319),
.B(n_3257),
.Y(n_3487)
);

INVxp67_ASAP7_75t_L g3488 ( 
.A(n_3424),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3413),
.B(n_3173),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3341),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_3328),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3331),
.A2(n_3286),
.B(n_3303),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3341),
.Y(n_3493)
);

NAND2xp33_ASAP7_75t_R g3494 ( 
.A(n_3347),
.B(n_3169),
.Y(n_3494)
);

HB1xp67_ASAP7_75t_L g3495 ( 
.A(n_3345),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3360),
.B(n_3284),
.Y(n_3496)
);

NAND2xp33_ASAP7_75t_SL g3497 ( 
.A(n_3429),
.B(n_3175),
.Y(n_3497)
);

OR2x2_ASAP7_75t_L g3498 ( 
.A(n_3359),
.B(n_3278),
.Y(n_3498)
);

AND2x2_ASAP7_75t_SL g3499 ( 
.A(n_3314),
.B(n_3261),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3428),
.B(n_3268),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_3358),
.B(n_3280),
.Y(n_3501)
);

NAND2xp33_ASAP7_75t_L g3502 ( 
.A(n_3331),
.B(n_3316),
.Y(n_3502)
);

NAND4xp25_ASAP7_75t_L g3503 ( 
.A(n_3377),
.B(n_3264),
.C(n_3273),
.D(n_3262),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3371),
.Y(n_3504)
);

INVx3_ASAP7_75t_SL g3505 ( 
.A(n_3397),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3324),
.B(n_3279),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3431),
.B(n_3336),
.Y(n_3507)
);

NAND2x1p5_ASAP7_75t_L g3508 ( 
.A(n_3347),
.B(n_3282),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3343),
.B(n_3271),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3371),
.Y(n_3510)
);

AOI21xp33_ASAP7_75t_L g3511 ( 
.A1(n_3379),
.A2(n_3269),
.B(n_3263),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3430),
.B(n_3270),
.Y(n_3512)
);

NAND3xp33_ASAP7_75t_L g3513 ( 
.A(n_3366),
.B(n_3285),
.C(n_3283),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3321),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3370),
.B(n_3195),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3343),
.B(n_3335),
.Y(n_3516)
);

OAI211xp5_ASAP7_75t_SL g3517 ( 
.A1(n_3358),
.A2(n_3296),
.B(n_3298),
.C(n_3289),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3307),
.B(n_3233),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3340),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3434),
.B(n_3302),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3394),
.B(n_3243),
.Y(n_3521)
);

NAND3xp33_ASAP7_75t_L g3522 ( 
.A(n_3366),
.B(n_3304),
.C(n_3269),
.Y(n_3522)
);

INVx1_ASAP7_75t_SL g3523 ( 
.A(n_3347),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_SL g3524 ( 
.A(n_3424),
.B(n_3301),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3429),
.B(n_3225),
.Y(n_3525)
);

NAND4xp25_ASAP7_75t_L g3526 ( 
.A(n_3350),
.B(n_3311),
.C(n_3312),
.D(n_3361),
.Y(n_3526)
);

INVx1_ASAP7_75t_SL g3527 ( 
.A(n_3315),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3340),
.Y(n_3528)
);

NAND2xp33_ASAP7_75t_R g3529 ( 
.A(n_3315),
.B(n_3230),
.Y(n_3529)
);

INVx2_ASAP7_75t_SL g3530 ( 
.A(n_3321),
.Y(n_3530)
);

BUFx2_ASAP7_75t_L g3531 ( 
.A(n_3407),
.Y(n_3531)
);

OR2x2_ASAP7_75t_L g3532 ( 
.A(n_3383),
.B(n_3247),
.Y(n_3532)
);

OR2x2_ASAP7_75t_L g3533 ( 
.A(n_3434),
.B(n_3248),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_3362),
.B(n_3251),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3395),
.B(n_3243),
.Y(n_3535)
);

OAI31xp33_ASAP7_75t_L g3536 ( 
.A1(n_3368),
.A2(n_3263),
.A3(n_3300),
.B(n_3275),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3326),
.B(n_3305),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3327),
.B(n_3300),
.Y(n_3538)
);

INVx1_ASAP7_75t_SL g3539 ( 
.A(n_3323),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3344),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3329),
.B(n_3235),
.Y(n_3541)
);

OR2x2_ASAP7_75t_L g3542 ( 
.A(n_3313),
.B(n_3082),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3397),
.B(n_3062),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3380),
.B(n_2830),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3401),
.B(n_3062),
.Y(n_3545)
);

NAND2x1_ASAP7_75t_L g3546 ( 
.A(n_3323),
.B(n_2845),
.Y(n_3546)
);

INVx2_ASAP7_75t_SL g3547 ( 
.A(n_3401),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3344),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3357),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3407),
.B(n_2831),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3357),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3402),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3348),
.B(n_2831),
.Y(n_3553)
);

NOR3xp33_ASAP7_75t_SL g3554 ( 
.A(n_3317),
.B(n_3246),
.C(n_3235),
.Y(n_3554)
);

AOI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_3349),
.A2(n_3051),
.B1(n_2917),
.B2(n_2908),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3402),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3403),
.Y(n_3557)
);

OR2x2_ASAP7_75t_L g3558 ( 
.A(n_3387),
.B(n_2927),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3353),
.B(n_2917),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3403),
.Y(n_3560)
);

INVx2_ASAP7_75t_SL g3561 ( 
.A(n_3468),
.Y(n_3561)
);

INVx5_ASAP7_75t_L g3562 ( 
.A(n_3491),
.Y(n_3562)
);

INVxp67_ASAP7_75t_SL g3563 ( 
.A(n_3508),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3444),
.B(n_3399),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3454),
.Y(n_3565)
);

AOI22xp33_ASAP7_75t_SL g3566 ( 
.A1(n_3502),
.A2(n_3421),
.B1(n_3338),
.B2(n_3373),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3508),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_L g3568 ( 
.A(n_3444),
.B(n_3372),
.Y(n_3568)
);

INVxp33_ASAP7_75t_L g3569 ( 
.A(n_3460),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3516),
.B(n_3364),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3523),
.B(n_3406),
.Y(n_3571)
);

INVxp67_ASAP7_75t_L g3572 ( 
.A(n_3486),
.Y(n_3572)
);

NOR2x1_ASAP7_75t_L g3573 ( 
.A(n_3491),
.B(n_3412),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3523),
.B(n_3408),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_3499),
.B(n_3338),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3507),
.B(n_3435),
.Y(n_3576)
);

INVxp67_ASAP7_75t_L g3577 ( 
.A(n_3495),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3452),
.Y(n_3578)
);

INVx1_ASAP7_75t_SL g3579 ( 
.A(n_3497),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3445),
.B(n_3436),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3480),
.B(n_3439),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3453),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3471),
.B(n_3374),
.Y(n_3583)
);

NAND2x1p5_ASAP7_75t_L g3584 ( 
.A(n_3531),
.B(n_3330),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3509),
.B(n_3376),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3505),
.B(n_3346),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_3468),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3470),
.B(n_3384),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3459),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3479),
.B(n_3355),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3455),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3482),
.B(n_3385),
.Y(n_3592)
);

OR2x2_ASAP7_75t_L g3593 ( 
.A(n_3467),
.B(n_3386),
.Y(n_3593)
);

OR2x2_ASAP7_75t_L g3594 ( 
.A(n_3451),
.B(n_3442),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3496),
.B(n_3388),
.Y(n_3595)
);

INVx2_ASAP7_75t_SL g3596 ( 
.A(n_3459),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3473),
.B(n_3391),
.Y(n_3597)
);

INVx2_ASAP7_75t_SL g3598 ( 
.A(n_3448),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3458),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3518),
.B(n_3500),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3461),
.Y(n_3601)
);

NAND2xp33_ASAP7_75t_SL g3602 ( 
.A(n_3554),
.B(n_3412),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3521),
.B(n_3393),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3462),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3464),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_SL g3606 ( 
.A(n_3522),
.B(n_3425),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3469),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3530),
.B(n_3396),
.Y(n_3608)
);

OR2x2_ASAP7_75t_L g3609 ( 
.A(n_3533),
.B(n_3325),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3477),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3485),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3535),
.B(n_3334),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3522),
.B(n_3425),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3514),
.B(n_3342),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_3490),
.Y(n_3615)
);

INVx6_ASAP7_75t_L g3616 ( 
.A(n_3515),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3493),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3504),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3510),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3546),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3449),
.B(n_3410),
.Y(n_3621)
);

INVx6_ASAP7_75t_L g3622 ( 
.A(n_3532),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3547),
.B(n_3337),
.Y(n_3623)
);

NOR2xp67_ASAP7_75t_L g3624 ( 
.A(n_3450),
.B(n_3474),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3443),
.B(n_3390),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3527),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3463),
.B(n_3352),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3527),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_SL g3629 ( 
.A(n_3483),
.B(n_3426),
.Y(n_3629)
);

HB1xp67_ASAP7_75t_L g3630 ( 
.A(n_3539),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3559),
.B(n_3382),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3481),
.B(n_3356),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3476),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3488),
.B(n_3544),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3553),
.B(n_3422),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_3526),
.B(n_3392),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3525),
.B(n_3411),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3539),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3534),
.B(n_3418),
.Y(n_3639)
);

OR2x2_ASAP7_75t_L g3640 ( 
.A(n_3526),
.B(n_3537),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3519),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3492),
.B(n_3416),
.Y(n_3642)
);

BUFx2_ASAP7_75t_L g3643 ( 
.A(n_3549),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3528),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3540),
.Y(n_3645)
);

INVx2_ASAP7_75t_SL g3646 ( 
.A(n_3548),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3501),
.B(n_3417),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3551),
.Y(n_3648)
);

NAND2x1p5_ASAP7_75t_L g3649 ( 
.A(n_3552),
.B(n_3426),
.Y(n_3649)
);

OAI31xp33_ASAP7_75t_L g3650 ( 
.A1(n_3465),
.A2(n_3423),
.A3(n_3427),
.B(n_3419),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3447),
.B(n_3432),
.Y(n_3651)
);

HB1xp67_ASAP7_75t_L g3652 ( 
.A(n_3529),
.Y(n_3652)
);

OR2x2_ASAP7_75t_L g3653 ( 
.A(n_3537),
.B(n_3433),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_L g3654 ( 
.A(n_3446),
.B(n_3438),
.Y(n_3654)
);

HB1xp67_ASAP7_75t_L g3655 ( 
.A(n_3556),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3557),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3498),
.B(n_3440),
.Y(n_3657)
);

INVxp67_ASAP7_75t_L g3658 ( 
.A(n_3652),
.Y(n_3658)
);

OAI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3652),
.A2(n_3513),
.B1(n_3472),
.B2(n_3456),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3630),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3569),
.B(n_3524),
.Y(n_3661)
);

AOI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_3602),
.A2(n_3465),
.B1(n_3457),
.B2(n_3494),
.Y(n_3662)
);

OAI31xp33_ASAP7_75t_L g3663 ( 
.A1(n_3602),
.A2(n_3513),
.A3(n_3503),
.B(n_3517),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3630),
.Y(n_3664)
);

HB1xp67_ASAP7_75t_L g3665 ( 
.A(n_3562),
.Y(n_3665)
);

AOI221xp5_ASAP7_75t_L g3666 ( 
.A1(n_3629),
.A2(n_3503),
.B1(n_3511),
.B2(n_3466),
.C(n_3545),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3570),
.B(n_3581),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3616),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3561),
.B(n_3560),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3561),
.B(n_3489),
.Y(n_3670)
);

OAI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_3566),
.A2(n_3542),
.B1(n_3555),
.B2(n_3475),
.Y(n_3671)
);

OAI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3575),
.A2(n_3511),
.B(n_3536),
.Y(n_3672)
);

INVxp67_ASAP7_75t_L g3673 ( 
.A(n_3563),
.Y(n_3673)
);

OAI21xp33_ASAP7_75t_L g3674 ( 
.A1(n_3569),
.A2(n_3550),
.B(n_3543),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3649),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3616),
.Y(n_3676)
);

OAI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3629),
.A2(n_3536),
.B(n_3520),
.Y(n_3677)
);

AOI22xp33_ASAP7_75t_SL g3678 ( 
.A1(n_3616),
.A2(n_3538),
.B1(n_3541),
.B2(n_3487),
.Y(n_3678)
);

OAI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_3575),
.A2(n_3538),
.B(n_3487),
.Y(n_3679)
);

OR2x2_ASAP7_75t_L g3680 ( 
.A(n_3571),
.B(n_3512),
.Y(n_3680)
);

HB1xp67_ASAP7_75t_L g3681 ( 
.A(n_3562),
.Y(n_3681)
);

OAI32xp33_ASAP7_75t_L g3682 ( 
.A1(n_3579),
.A2(n_3541),
.A3(n_3478),
.B1(n_3484),
.B2(n_3506),
.Y(n_3682)
);

NAND4xp25_ASAP7_75t_SL g3683 ( 
.A(n_3566),
.B(n_3484),
.C(n_3506),
.D(n_3558),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3622),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3596),
.B(n_3441),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3622),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3622),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3649),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3576),
.B(n_2894),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3600),
.B(n_2894),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3596),
.B(n_2908),
.Y(n_3691)
);

NAND2xp33_ASAP7_75t_L g3692 ( 
.A(n_3584),
.B(n_3246),
.Y(n_3692)
);

AOI21xp33_ASAP7_75t_L g3693 ( 
.A1(n_3563),
.A2(n_3253),
.B(n_2910),
.Y(n_3693)
);

AOI22xp5_ASAP7_75t_L g3694 ( 
.A1(n_3654),
.A2(n_3253),
.B1(n_3051),
.B2(n_2904),
.Y(n_3694)
);

AOI21xp5_ASAP7_75t_L g3695 ( 
.A1(n_3606),
.A2(n_2904),
.B(n_2959),
.Y(n_3695)
);

OAI22xp33_ASAP7_75t_L g3696 ( 
.A1(n_3640),
.A2(n_2904),
.B1(n_2867),
.B2(n_2891),
.Y(n_3696)
);

AOI21xp33_ASAP7_75t_SL g3697 ( 
.A1(n_3584),
.A2(n_3613),
.B(n_3606),
.Y(n_3697)
);

A2O1A1Ixp33_ASAP7_75t_L g3698 ( 
.A1(n_3654),
.A2(n_3613),
.B(n_3642),
.C(n_3650),
.Y(n_3698)
);

OAI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3636),
.A2(n_3628),
.B1(n_3638),
.B2(n_3626),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3573),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3580),
.B(n_2927),
.Y(n_3701)
);

OAI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3572),
.A2(n_2867),
.B1(n_2891),
.B2(n_2863),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3597),
.B(n_2966),
.Y(n_3703)
);

OAI322xp33_ASAP7_75t_L g3704 ( 
.A1(n_3572),
.A2(n_2924),
.A3(n_2923),
.B1(n_2921),
.B2(n_2912),
.C1(n_2893),
.C2(n_2863),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3655),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3567),
.B(n_2963),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_SL g3707 ( 
.A1(n_3637),
.A2(n_3639),
.B1(n_3568),
.B2(n_3565),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3655),
.Y(n_3708)
);

XNOR2x1_ASAP7_75t_L g3709 ( 
.A(n_3634),
.B(n_2065),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3603),
.B(n_2805),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3574),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3562),
.Y(n_3712)
);

INVx2_ASAP7_75t_SL g3713 ( 
.A(n_3562),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3567),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3564),
.Y(n_3715)
);

AO22x1_ASAP7_75t_L g3716 ( 
.A1(n_3587),
.A2(n_2912),
.B1(n_2921),
.B2(n_2893),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3595),
.Y(n_3717)
);

OR2x2_ASAP7_75t_L g3718 ( 
.A(n_3587),
.B(n_2805),
.Y(n_3718)
);

NOR2xp67_ASAP7_75t_L g3719 ( 
.A(n_3577),
.B(n_2832),
.Y(n_3719)
);

INVx2_ASAP7_75t_SL g3720 ( 
.A(n_3598),
.Y(n_3720)
);

AOI22xp33_ASAP7_75t_L g3721 ( 
.A1(n_3621),
.A2(n_2924),
.B1(n_2923),
.B2(n_2838),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3598),
.B(n_2832),
.Y(n_3722)
);

NOR4xp25_ASAP7_75t_L g3723 ( 
.A(n_3577),
.B(n_3646),
.C(n_3615),
.D(n_3610),
.Y(n_3723)
);

NAND3xp33_ASAP7_75t_SL g3724 ( 
.A(n_3590),
.B(n_2843),
.C(n_2838),
.Y(n_3724)
);

NAND2xp33_ASAP7_75t_SL g3725 ( 
.A(n_3609),
.B(n_2616),
.Y(n_3725)
);

OAI221xp5_ASAP7_75t_L g3726 ( 
.A1(n_3624),
.A2(n_2861),
.B1(n_2848),
.B2(n_2843),
.C(n_2616),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3568),
.B(n_2848),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3589),
.B(n_2861),
.Y(n_3728)
);

XNOR2xp5_ASAP7_75t_L g3729 ( 
.A(n_3631),
.B(n_2249),
.Y(n_3729)
);

OAI21xp33_ASAP7_75t_L g3730 ( 
.A1(n_3625),
.A2(n_2067),
.B(n_2065),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3592),
.B(n_3586),
.Y(n_3731)
);

NOR2x1_ASAP7_75t_L g3732 ( 
.A(n_3589),
.B(n_2615),
.Y(n_3732)
);

INVxp67_ASAP7_75t_L g3733 ( 
.A(n_3643),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3620),
.B(n_2615),
.Y(n_3734)
);

AOI322xp5_ASAP7_75t_L g3735 ( 
.A1(n_3647),
.A2(n_2725),
.A3(n_2719),
.B1(n_2721),
.B2(n_2766),
.C1(n_2723),
.C2(n_2759),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3612),
.Y(n_3736)
);

INVxp67_ASAP7_75t_L g3737 ( 
.A(n_3623),
.Y(n_3737)
);

AOI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3627),
.A2(n_2690),
.B(n_2634),
.Y(n_3738)
);

INVxp67_ASAP7_75t_L g3739 ( 
.A(n_3608),
.Y(n_3739)
);

AOI22xp5_ASAP7_75t_L g3740 ( 
.A1(n_3635),
.A2(n_2097),
.B1(n_2634),
.B2(n_2067),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3633),
.B(n_2639),
.Y(n_3741)
);

INVxp67_ASAP7_75t_SL g3742 ( 
.A(n_3620),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3585),
.Y(n_3743)
);

NOR3xp33_ASAP7_75t_L g3744 ( 
.A(n_3632),
.B(n_2687),
.C(n_2667),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3667),
.B(n_3651),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3668),
.B(n_3633),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3676),
.B(n_3617),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3665),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3681),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3672),
.B(n_3615),
.Y(n_3750)
);

AOI221xp5_ASAP7_75t_L g3751 ( 
.A1(n_3697),
.A2(n_3618),
.B1(n_3619),
.B2(n_3578),
.C(n_3599),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3684),
.B(n_3588),
.Y(n_3752)
);

INVxp67_ASAP7_75t_L g3753 ( 
.A(n_3686),
.Y(n_3753)
);

A2O1A1Ixp33_ASAP7_75t_L g3754 ( 
.A1(n_3663),
.A2(n_3610),
.B(n_3605),
.C(n_3646),
.Y(n_3754)
);

HB1xp67_ASAP7_75t_L g3755 ( 
.A(n_3687),
.Y(n_3755)
);

NAND2x1_ASAP7_75t_L g3756 ( 
.A(n_3675),
.B(n_3605),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3690),
.B(n_3593),
.Y(n_3757)
);

OR2x2_ASAP7_75t_L g3758 ( 
.A(n_3720),
.B(n_3583),
.Y(n_3758)
);

INVxp67_ASAP7_75t_SL g3759 ( 
.A(n_3692),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3689),
.B(n_3594),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_3674),
.B(n_3657),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3713),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3707),
.B(n_3582),
.Y(n_3763)
);

INVxp67_ASAP7_75t_L g3764 ( 
.A(n_3661),
.Y(n_3764)
);

OAI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_3662),
.A2(n_3653),
.B1(n_3601),
.B2(n_3604),
.Y(n_3765)
);

OAI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3672),
.A2(n_3607),
.B(n_3591),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3742),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3678),
.B(n_3611),
.Y(n_3768)
);

AO22x1_ASAP7_75t_L g3769 ( 
.A1(n_3677),
.A2(n_3656),
.B1(n_3641),
.B2(n_3645),
.Y(n_3769)
);

INVxp67_ASAP7_75t_L g3770 ( 
.A(n_3660),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3658),
.B(n_3614),
.Y(n_3771)
);

AND2x4_ASAP7_75t_L g3772 ( 
.A(n_3688),
.B(n_3656),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3705),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3673),
.B(n_3644),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3664),
.B(n_3648),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3708),
.Y(n_3776)
);

NAND2xp33_ASAP7_75t_L g3777 ( 
.A(n_3698),
.B(n_2667),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3717),
.B(n_2667),
.Y(n_3778)
);

INVx1_ASAP7_75t_SL g3779 ( 
.A(n_3700),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3723),
.B(n_2639),
.Y(n_3780)
);

AOI211x1_ASAP7_75t_L g3781 ( 
.A1(n_3679),
.A2(n_2641),
.B(n_2645),
.C(n_2642),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3719),
.Y(n_3782)
);

HB1xp67_ASAP7_75t_L g3783 ( 
.A(n_3732),
.Y(n_3783)
);

INVx1_ASAP7_75t_SL g3784 ( 
.A(n_3680),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3712),
.Y(n_3785)
);

NOR2xp33_ASAP7_75t_L g3786 ( 
.A(n_3682),
.B(n_2687),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3670),
.B(n_2718),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3736),
.B(n_3663),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3669),
.Y(n_3789)
);

HB1xp67_ASAP7_75t_L g3790 ( 
.A(n_3723),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3714),
.B(n_2687),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3685),
.Y(n_3792)
);

NOR3xp33_ASAP7_75t_L g3793 ( 
.A(n_3659),
.B(n_2728),
.C(n_2240),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3715),
.B(n_2716),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3722),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3722),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_3733),
.B(n_2728),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3703),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3718),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3711),
.B(n_2756),
.Y(n_3800)
);

NAND2x1p5_ASAP7_75t_L g3801 ( 
.A(n_3731),
.B(n_2728),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3710),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3706),
.Y(n_3803)
);

NAND2x1_ASAP7_75t_L g3804 ( 
.A(n_3734),
.B(n_2718),
.Y(n_3804)
);

OAI22x1_ASAP7_75t_L g3805 ( 
.A1(n_3683),
.A2(n_2524),
.B1(n_2539),
.B2(n_2526),
.Y(n_3805)
);

OR2x2_ASAP7_75t_L g3806 ( 
.A(n_3691),
.B(n_2719),
.Y(n_3806)
);

NOR2x1_ASAP7_75t_L g3807 ( 
.A(n_3679),
.B(n_2641),
.Y(n_3807)
);

NAND4xp25_ASAP7_75t_L g3808 ( 
.A(n_3666),
.B(n_2489),
.C(n_2260),
.D(n_2459),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3706),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3699),
.B(n_2019),
.Y(n_3810)
);

OR2x2_ASAP7_75t_L g3811 ( 
.A(n_3671),
.B(n_2721),
.Y(n_3811)
);

INVx1_ASAP7_75t_SL g3812 ( 
.A(n_3725),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3728),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_3739),
.B(n_2734),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3701),
.Y(n_3815)
);

CKINVDCx5p33_ASAP7_75t_R g3816 ( 
.A(n_3737),
.Y(n_3816)
);

NOR2xp33_ASAP7_75t_L g3817 ( 
.A(n_3709),
.B(n_2734),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3729),
.B(n_2642),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3727),
.B(n_2645),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3743),
.B(n_2671),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3741),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3734),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3695),
.A2(n_2750),
.B(n_2736),
.Y(n_3823)
);

NOR2x1_ASAP7_75t_R g3824 ( 
.A(n_3693),
.B(n_2019),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3745),
.B(n_3757),
.Y(n_3825)
);

OAI21xp33_ASAP7_75t_L g3826 ( 
.A1(n_3808),
.A2(n_3730),
.B(n_3694),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3756),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3760),
.B(n_3740),
.Y(n_3828)
);

CKINVDCx20_ASAP7_75t_R g3829 ( 
.A(n_3816),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3782),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3746),
.Y(n_3831)
);

HB1xp67_ASAP7_75t_L g3832 ( 
.A(n_3790),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3755),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3795),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3796),
.Y(n_3835)
);

NAND3xp33_ASAP7_75t_L g3836 ( 
.A(n_3754),
.B(n_3744),
.C(n_3721),
.Y(n_3836)
);

NOR2xp33_ASAP7_75t_L g3837 ( 
.A(n_3812),
.B(n_3724),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3803),
.Y(n_3838)
);

OR2x2_ASAP7_75t_L g3839 ( 
.A(n_3784),
.B(n_3702),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3809),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3762),
.B(n_3716),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3822),
.Y(n_3842)
);

CKINVDCx14_ASAP7_75t_R g3843 ( 
.A(n_3763),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3748),
.B(n_3696),
.Y(n_3844)
);

OR2x2_ASAP7_75t_L g3845 ( 
.A(n_3784),
.B(n_3726),
.Y(n_3845)
);

OR2x2_ASAP7_75t_L g3846 ( 
.A(n_3758),
.B(n_3738),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3749),
.Y(n_3847)
);

NOR3xp33_ASAP7_75t_SL g3848 ( 
.A(n_3765),
.B(n_3704),
.C(n_3735),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_3812),
.B(n_3735),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3783),
.Y(n_3850)
);

INVx2_ASAP7_75t_SL g3851 ( 
.A(n_3772),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3752),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3767),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3807),
.Y(n_3854)
);

NAND3xp33_ASAP7_75t_L g3855 ( 
.A(n_3750),
.B(n_3704),
.C(n_2772),
.Y(n_3855)
);

O2A1O1Ixp33_ASAP7_75t_L g3856 ( 
.A1(n_3750),
.A2(n_2735),
.B(n_2739),
.C(n_2726),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3772),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3769),
.B(n_2736),
.Y(n_3858)
);

AOI32xp33_ASAP7_75t_L g3859 ( 
.A1(n_3777),
.A2(n_2416),
.A3(n_2523),
.B1(n_2524),
.B2(n_2539),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_3779),
.B(n_2019),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3815),
.B(n_2756),
.Y(n_3861)
);

CKINVDCx5p33_ASAP7_75t_R g3862 ( 
.A(n_3764),
.Y(n_3862)
);

NOR2x1p5_ASAP7_75t_SL g3863 ( 
.A(n_3811),
.B(n_2735),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3785),
.B(n_2750),
.Y(n_3864)
);

OR2x2_ASAP7_75t_L g3865 ( 
.A(n_3768),
.B(n_2723),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3779),
.B(n_2019),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3753),
.B(n_2297),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3794),
.B(n_3800),
.Y(n_3868)
);

NOR3xp33_ASAP7_75t_SL g3869 ( 
.A(n_3765),
.B(n_2772),
.C(n_2769),
.Y(n_3869)
);

HB1xp67_ASAP7_75t_L g3870 ( 
.A(n_3801),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_L g3871 ( 
.A(n_3770),
.B(n_2754),
.Y(n_3871)
);

NOR3xp33_ASAP7_75t_SL g3872 ( 
.A(n_3788),
.B(n_2726),
.C(n_2724),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3761),
.B(n_2754),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3759),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3747),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3798),
.Y(n_3876)
);

OAI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3780),
.A2(n_2416),
.B1(n_2526),
.B2(n_2208),
.Y(n_3877)
);

NAND2x1_ASAP7_75t_L g3878 ( 
.A(n_3799),
.B(n_2724),
.Y(n_3878)
);

INVxp67_ASAP7_75t_L g3879 ( 
.A(n_3824),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3802),
.B(n_2771),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3771),
.B(n_2755),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3780),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3766),
.B(n_3789),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3774),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3773),
.B(n_2771),
.Y(n_3885)
);

OR2x2_ASAP7_75t_L g3886 ( 
.A(n_3775),
.B(n_3778),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3776),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3766),
.Y(n_3888)
);

AOI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3793),
.A2(n_2489),
.B1(n_2264),
.B2(n_2019),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3786),
.A2(n_2264),
.B1(n_2208),
.B2(n_2229),
.Y(n_3890)
);

INVxp67_ASAP7_75t_L g3891 ( 
.A(n_3825),
.Y(n_3891)
);

NOR3x1_ASAP7_75t_L g3892 ( 
.A(n_3836),
.B(n_3810),
.C(n_3792),
.Y(n_3892)
);

NOR2x1_ASAP7_75t_L g3893 ( 
.A(n_3839),
.B(n_3813),
.Y(n_3893)
);

NOR2xp33_ASAP7_75t_SL g3894 ( 
.A(n_3851),
.B(n_3797),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3867),
.B(n_3817),
.Y(n_3895)
);

AOI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3832),
.A2(n_3805),
.B(n_3751),
.Y(n_3896)
);

OAI21xp5_ASAP7_75t_SL g3897 ( 
.A1(n_3843),
.A2(n_3818),
.B(n_3814),
.Y(n_3897)
);

NAND4xp25_ASAP7_75t_L g3898 ( 
.A(n_3826),
.B(n_3791),
.C(n_3820),
.D(n_3787),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3857),
.Y(n_3899)
);

NAND4xp25_ASAP7_75t_L g3900 ( 
.A(n_3837),
.B(n_3821),
.C(n_3806),
.D(n_3819),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_L g3901 ( 
.A(n_3831),
.B(n_3801),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3833),
.B(n_3781),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3863),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3827),
.B(n_3804),
.Y(n_3904)
);

OR2x2_ASAP7_75t_L g3905 ( 
.A(n_3841),
.B(n_3823),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3829),
.Y(n_3906)
);

NAND4xp25_ASAP7_75t_L g3907 ( 
.A(n_3828),
.B(n_2260),
.C(n_2459),
.D(n_2449),
.Y(n_3907)
);

OAI21xp5_ASAP7_75t_SL g3908 ( 
.A1(n_3879),
.A2(n_2270),
.B(n_2208),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3848),
.B(n_2107),
.Y(n_3909)
);

NAND4xp25_ASAP7_75t_L g3910 ( 
.A(n_3844),
.B(n_2449),
.C(n_2041),
.D(n_2497),
.Y(n_3910)
);

NOR4xp25_ASAP7_75t_L g3911 ( 
.A(n_3888),
.B(n_2766),
.C(n_2753),
.D(n_2744),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3861),
.B(n_2755),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3868),
.B(n_2758),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3842),
.B(n_2758),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3874),
.B(n_2764),
.Y(n_3915)
);

NAND4xp25_ASAP7_75t_L g3916 ( 
.A(n_3852),
.B(n_2497),
.C(n_2452),
.D(n_2406),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3847),
.B(n_2764),
.Y(n_3917)
);

AOI22xp5_ASAP7_75t_L g3918 ( 
.A1(n_3862),
.A2(n_2272),
.B1(n_2107),
.B2(n_2229),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3841),
.Y(n_3919)
);

NAND3xp33_ASAP7_75t_L g3920 ( 
.A(n_3848),
.B(n_2704),
.C(n_2732),
.Y(n_3920)
);

OAI211xp5_ASAP7_75t_L g3921 ( 
.A1(n_3849),
.A2(n_2759),
.B(n_2753),
.C(n_2732),
.Y(n_3921)
);

AOI221xp5_ASAP7_75t_L g3922 ( 
.A1(n_3883),
.A2(n_2744),
.B1(n_2743),
.B2(n_2741),
.C(n_2733),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3834),
.B(n_3835),
.Y(n_3923)
);

NOR2x1_ASAP7_75t_L g3924 ( 
.A(n_3854),
.B(n_2733),
.Y(n_3924)
);

NAND4xp75_ASAP7_75t_L g3925 ( 
.A(n_3844),
.B(n_2704),
.C(n_2743),
.D(n_2741),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3882),
.A2(n_2603),
.B(n_2587),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3838),
.B(n_2603),
.Y(n_3927)
);

BUFx3_ASAP7_75t_L g3928 ( 
.A(n_3840),
.Y(n_3928)
);

NOR3xp33_ASAP7_75t_L g3929 ( 
.A(n_3830),
.B(n_2272),
.C(n_2614),
.Y(n_3929)
);

OAI211xp5_ASAP7_75t_SL g3930 ( 
.A1(n_3845),
.A2(n_2632),
.B(n_2614),
.C(n_2622),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3870),
.A2(n_2624),
.B(n_2622),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3878),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3850),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3876),
.B(n_2624),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3846),
.Y(n_3935)
);

AOI221x1_ASAP7_75t_L g3936 ( 
.A1(n_3853),
.A2(n_2627),
.B1(n_2632),
.B2(n_2666),
.C(n_2701),
.Y(n_3936)
);

AND2x2_ASAP7_75t_L g3937 ( 
.A(n_3879),
.B(n_2637),
.Y(n_3937)
);

NOR2xp67_ASAP7_75t_L g3938 ( 
.A(n_3855),
.B(n_2627),
.Y(n_3938)
);

NAND3xp33_ASAP7_75t_L g3939 ( 
.A(n_3887),
.B(n_2704),
.C(n_2638),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3858),
.Y(n_3940)
);

OAI211xp5_ASAP7_75t_L g3941 ( 
.A1(n_3860),
.A2(n_3866),
.B(n_3858),
.C(n_3875),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3873),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_SL g3943 ( 
.A(n_3884),
.B(n_3886),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3891),
.B(n_3872),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3906),
.B(n_3869),
.Y(n_3945)
);

NAND3xp33_ASAP7_75t_SL g3946 ( 
.A(n_3896),
.B(n_3859),
.C(n_3865),
.Y(n_3946)
);

NOR2x1_ASAP7_75t_L g3947 ( 
.A(n_3893),
.B(n_3864),
.Y(n_3947)
);

NOR4xp75_ASAP7_75t_L g3948 ( 
.A(n_3909),
.B(n_3864),
.C(n_3885),
.D(n_3880),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3899),
.B(n_3871),
.Y(n_3949)
);

OAI33xp33_ASAP7_75t_L g3950 ( 
.A1(n_3919),
.A2(n_3877),
.A3(n_3885),
.B1(n_3880),
.B2(n_3856),
.B3(n_3881),
.Y(n_3950)
);

NOR3xp33_ASAP7_75t_L g3951 ( 
.A(n_3897),
.B(n_3889),
.C(n_3890),
.Y(n_3951)
);

AOI211xp5_ASAP7_75t_L g3952 ( 
.A1(n_3921),
.A2(n_3856),
.B(n_2208),
.C(n_2229),
.Y(n_3952)
);

NAND3xp33_ASAP7_75t_L g3953 ( 
.A(n_3894),
.B(n_2208),
.C(n_2107),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_L g3954 ( 
.A(n_3928),
.B(n_2637),
.Y(n_3954)
);

A2O1A1Ixp33_ASAP7_75t_L g3955 ( 
.A1(n_3920),
.A2(n_2705),
.B(n_2701),
.C(n_2638),
.Y(n_3955)
);

NAND2x1_ASAP7_75t_SL g3956 ( 
.A(n_3903),
.B(n_3932),
.Y(n_3956)
);

O2A1O1Ixp33_ASAP7_75t_L g3957 ( 
.A1(n_3904),
.A2(n_2705),
.B(n_2644),
.C(n_2666),
.Y(n_3957)
);

NOR4xp25_ASAP7_75t_SL g3958 ( 
.A(n_3940),
.B(n_2190),
.C(n_2483),
.D(n_2487),
.Y(n_3958)
);

NOR3xp33_ASAP7_75t_L g3959 ( 
.A(n_3900),
.B(n_2174),
.C(n_2164),
.Y(n_3959)
);

NAND4xp25_ASAP7_75t_L g3960 ( 
.A(n_3892),
.B(n_2452),
.C(n_2406),
.D(n_2411),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3942),
.B(n_2644),
.Y(n_3961)
);

AND2x4_ASAP7_75t_L g3962 ( 
.A(n_3895),
.B(n_3935),
.Y(n_3962)
);

NOR3xp33_ASAP7_75t_L g3963 ( 
.A(n_3898),
.B(n_3923),
.C(n_3941),
.Y(n_3963)
);

NOR2x1_ASAP7_75t_L g3964 ( 
.A(n_3905),
.B(n_2653),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3933),
.B(n_2653),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3943),
.A2(n_2656),
.B(n_2704),
.Y(n_3966)
);

AOI211xp5_ASAP7_75t_L g3967 ( 
.A1(n_3901),
.A2(n_2229),
.B(n_2107),
.C(n_2239),
.Y(n_3967)
);

NAND3xp33_ASAP7_75t_SL g3968 ( 
.A(n_3902),
.B(n_2656),
.C(n_2246),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3924),
.Y(n_3969)
);

NOR3xp33_ASAP7_75t_L g3970 ( 
.A(n_3908),
.B(n_2250),
.C(n_2411),
.Y(n_3970)
);

OAI21xp33_ASAP7_75t_L g3971 ( 
.A1(n_3907),
.A2(n_2402),
.B(n_2447),
.Y(n_3971)
);

NAND4xp25_ASAP7_75t_L g3972 ( 
.A(n_3915),
.B(n_3937),
.C(n_3927),
.D(n_3914),
.Y(n_3972)
);

NOR4xp75_ASAP7_75t_L g3973 ( 
.A(n_3925),
.B(n_2445),
.C(n_2402),
.D(n_2447),
.Y(n_3973)
);

AOI211xp5_ASAP7_75t_L g3974 ( 
.A1(n_3920),
.A2(n_2107),
.B(n_2229),
.C(n_2478),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3913),
.B(n_2445),
.Y(n_3975)
);

NAND3xp33_ASAP7_75t_L g3976 ( 
.A(n_3929),
.B(n_2049),
.C(n_2478),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3938),
.B(n_2478),
.Y(n_3977)
);

NAND3x1_ASAP7_75t_L g3978 ( 
.A(n_3917),
.B(n_2488),
.C(n_2400),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3934),
.B(n_2483),
.Y(n_3979)
);

NAND3x1_ASAP7_75t_L g3980 ( 
.A(n_3918),
.B(n_3912),
.C(n_3931),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3934),
.B(n_2512),
.Y(n_3981)
);

OAI21xp33_ASAP7_75t_SL g3982 ( 
.A1(n_3910),
.A2(n_2438),
.B(n_2378),
.Y(n_3982)
);

NAND3xp33_ASAP7_75t_L g3983 ( 
.A(n_3939),
.B(n_2082),
.C(n_2096),
.Y(n_3983)
);

AOI21xp5_ASAP7_75t_L g3984 ( 
.A1(n_3926),
.A2(n_2543),
.B(n_2540),
.Y(n_3984)
);

NOR3xp33_ASAP7_75t_L g3985 ( 
.A(n_3930),
.B(n_2250),
.C(n_2207),
.Y(n_3985)
);

AND4x1_ASAP7_75t_L g3986 ( 
.A(n_3911),
.B(n_2488),
.C(n_2220),
.D(n_2221),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3916),
.B(n_2417),
.Y(n_3987)
);

NOR2x1_ASAP7_75t_L g3988 ( 
.A(n_3939),
.B(n_2487),
.Y(n_3988)
);

NOR3xp33_ASAP7_75t_L g3989 ( 
.A(n_3916),
.B(n_2207),
.C(n_2222),
.Y(n_3989)
);

O2A1O1Ixp33_ASAP7_75t_SL g3990 ( 
.A1(n_3922),
.A2(n_2413),
.B(n_2540),
.C(n_2538),
.Y(n_3990)
);

NAND5xp2_ASAP7_75t_L g3991 ( 
.A(n_3936),
.B(n_2242),
.C(n_2221),
.D(n_2220),
.E(n_2378),
.Y(n_3991)
);

AOI221xp5_ASAP7_75t_L g3992 ( 
.A1(n_3946),
.A2(n_3963),
.B1(n_3950),
.B2(n_3953),
.C(n_3951),
.Y(n_3992)
);

NAND3x1_ASAP7_75t_SL g3993 ( 
.A(n_3947),
.B(n_2400),
.C(n_2372),
.Y(n_3993)
);

NOR2xp33_ASAP7_75t_L g3994 ( 
.A(n_3962),
.B(n_2493),
.Y(n_3994)
);

OR2x2_ASAP7_75t_L g3995 ( 
.A(n_3960),
.B(n_2369),
.Y(n_3995)
);

CKINVDCx5p33_ASAP7_75t_R g3996 ( 
.A(n_3962),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3956),
.Y(n_3997)
);

AOI221x1_ASAP7_75t_L g3998 ( 
.A1(n_3969),
.A2(n_2543),
.B1(n_2538),
.B2(n_2531),
.C(n_2530),
.Y(n_3998)
);

AOI22xp33_ASAP7_75t_L g3999 ( 
.A1(n_3959),
.A2(n_3987),
.B1(n_3944),
.B2(n_3989),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3954),
.B(n_3952),
.Y(n_4000)
);

A2O1A1Ixp33_ASAP7_75t_SL g4001 ( 
.A1(n_3949),
.A2(n_2485),
.B(n_2481),
.C(n_2474),
.Y(n_4001)
);

OAI221xp5_ASAP7_75t_SL g4002 ( 
.A1(n_3945),
.A2(n_2413),
.B1(n_2438),
.B2(n_2372),
.C(n_2512),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3964),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3971),
.A2(n_2161),
.B1(n_2207),
.B2(n_2222),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3965),
.B(n_2493),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3948),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3981),
.B(n_2494),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_L g4008 ( 
.A(n_3974),
.B(n_2494),
.Y(n_4008)
);

AOI221xp5_ASAP7_75t_L g4009 ( 
.A1(n_3968),
.A2(n_2531),
.B1(n_2530),
.B2(n_2529),
.C(n_2518),
.Y(n_4009)
);

HB1xp67_ASAP7_75t_L g4010 ( 
.A(n_3973),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3961),
.Y(n_4011)
);

OAI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3980),
.A2(n_3972),
.B(n_3966),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3977),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3979),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3975),
.B(n_3967),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3986),
.B(n_2496),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3970),
.B(n_2496),
.Y(n_4017)
);

INVxp67_ASAP7_75t_SL g4018 ( 
.A(n_3988),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3958),
.B(n_2506),
.Y(n_4019)
);

OAI211xp5_ASAP7_75t_L g4020 ( 
.A1(n_3960),
.A2(n_2529),
.B(n_2518),
.C(n_2506),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3978),
.B(n_2510),
.Y(n_4021)
);

NOR2x1_ASAP7_75t_L g4022 ( 
.A(n_3991),
.B(n_2510),
.Y(n_4022)
);

XOR2x2_ASAP7_75t_L g4023 ( 
.A(n_3985),
.B(n_2242),
.Y(n_4023)
);

HB1xp67_ASAP7_75t_L g4024 ( 
.A(n_3983),
.Y(n_4024)
);

AOI22xp5_ASAP7_75t_L g4025 ( 
.A1(n_3982),
.A2(n_2396),
.B1(n_2511),
.B2(n_2513),
.Y(n_4025)
);

AOI222xp33_ASAP7_75t_L g4026 ( 
.A1(n_3976),
.A2(n_2511),
.B1(n_2513),
.B2(n_2082),
.C1(n_2078),
.C2(n_2096),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3996),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_4012),
.A2(n_3957),
.B(n_3984),
.Y(n_4028)
);

NAND2x1p5_ASAP7_75t_SL g4029 ( 
.A(n_4022),
.B(n_3990),
.Y(n_4029)
);

NAND4xp75_ASAP7_75t_L g4030 ( 
.A(n_3992),
.B(n_3955),
.C(n_2396),
.D(n_2160),
.Y(n_4030)
);

NAND3xp33_ASAP7_75t_SL g4031 ( 
.A(n_3997),
.B(n_2063),
.C(n_2515),
.Y(n_4031)
);

NOR3xp33_ASAP7_75t_L g4032 ( 
.A(n_4006),
.B(n_2222),
.C(n_2248),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3993),
.Y(n_4033)
);

AND2x4_ASAP7_75t_L g4034 ( 
.A(n_4013),
.B(n_2474),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_4010),
.B(n_2329),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_SL g4036 ( 
.A(n_4012),
.B(n_2481),
.Y(n_4036)
);

OR2x2_ASAP7_75t_L g4037 ( 
.A(n_4000),
.B(n_2485),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_SL g4038 ( 
.A(n_4003),
.B(n_2508),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3999),
.B(n_2508),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_4018),
.Y(n_4040)
);

NOR2x1_ASAP7_75t_L g4041 ( 
.A(n_4011),
.B(n_2514),
.Y(n_4041)
);

NOR2x1p5_ASAP7_75t_L g4042 ( 
.A(n_4015),
.B(n_2063),
.Y(n_4042)
);

NOR2x1_ASAP7_75t_SL g4043 ( 
.A(n_4019),
.B(n_4014),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_4024),
.Y(n_4044)
);

AND2x2_ASAP7_75t_SL g4045 ( 
.A(n_3994),
.B(n_2133),
.Y(n_4045)
);

INVxp67_ASAP7_75t_SL g4046 ( 
.A(n_4019),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_4023),
.B(n_4005),
.Y(n_4047)
);

NOR2xp67_ASAP7_75t_L g4048 ( 
.A(n_4021),
.B(n_2514),
.Y(n_4048)
);

NAND3xp33_ASAP7_75t_L g4049 ( 
.A(n_4008),
.B(n_2078),
.C(n_2075),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_4016),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3995),
.Y(n_4051)
);

NOR3xp33_ASAP7_75t_L g4052 ( 
.A(n_4017),
.B(n_2248),
.C(n_2230),
.Y(n_4052)
);

OAI21xp33_ASAP7_75t_SL g4053 ( 
.A1(n_4009),
.A2(n_2068),
.B(n_2073),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_4007),
.Y(n_4054)
);

CKINVDCx16_ASAP7_75t_R g4055 ( 
.A(n_4025),
.Y(n_4055)
);

OAI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_4033),
.A2(n_4002),
.B1(n_4004),
.B2(n_4020),
.Y(n_4056)
);

INVx1_ASAP7_75t_SL g4057 ( 
.A(n_4035),
.Y(n_4057)
);

AND3x4_ASAP7_75t_L g4058 ( 
.A(n_4034),
.B(n_4001),
.C(n_3998),
.Y(n_4058)
);

AOI211xp5_ASAP7_75t_L g4059 ( 
.A1(n_4040),
.A2(n_4026),
.B(n_2075),
.C(n_2068),
.Y(n_4059)
);

AND3x2_ASAP7_75t_L g4060 ( 
.A(n_4046),
.B(n_2073),
.C(n_2071),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_4029),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_4043),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_4042),
.B(n_2329),
.Y(n_4063)
);

OAI321xp33_ASAP7_75t_L g4064 ( 
.A1(n_4044),
.A2(n_2071),
.A3(n_2069),
.B1(n_2204),
.B2(n_2160),
.C(n_2516),
.Y(n_4064)
);

NAND4xp75_ASAP7_75t_L g4065 ( 
.A(n_4027),
.B(n_2069),
.C(n_2334),
.D(n_2515),
.Y(n_4065)
);

BUFx2_ASAP7_75t_L g4066 ( 
.A(n_4034),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_4030),
.Y(n_4067)
);

BUFx2_ASAP7_75t_L g4068 ( 
.A(n_4041),
.Y(n_4068)
);

XOR2x1_ASAP7_75t_L g4069 ( 
.A(n_4051),
.B(n_2516),
.Y(n_4069)
);

AOI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_4032),
.A2(n_2194),
.B1(n_2050),
.B2(n_2226),
.Y(n_4070)
);

XOR2x1_ASAP7_75t_L g4071 ( 
.A(n_4050),
.B(n_2420),
.Y(n_4071)
);

AND4x1_ASAP7_75t_L g4072 ( 
.A(n_4054),
.B(n_2057),
.C(n_2089),
.D(n_2334),
.Y(n_4072)
);

INVx1_ASAP7_75t_SL g4073 ( 
.A(n_4047),
.Y(n_4073)
);

AOI221xp5_ASAP7_75t_L g4074 ( 
.A1(n_4036),
.A2(n_2306),
.B1(n_2471),
.B2(n_2446),
.C(n_2433),
.Y(n_4074)
);

OR2x6_ASAP7_75t_L g4075 ( 
.A(n_4028),
.B(n_2036),
.Y(n_4075)
);

NAND4xp75_ASAP7_75t_L g4076 ( 
.A(n_4041),
.B(n_2089),
.C(n_2057),
.D(n_2500),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_4055),
.B(n_2369),
.Y(n_4077)
);

AOI211xp5_ASAP7_75t_L g4078 ( 
.A1(n_4039),
.A2(n_2349),
.B(n_2471),
.C(n_2332),
.Y(n_4078)
);

INVxp67_ASAP7_75t_L g4079 ( 
.A(n_4038),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_L g4080 ( 
.A(n_4045),
.B(n_2369),
.Y(n_4080)
);

NOR4xp75_ASAP7_75t_L g4081 ( 
.A(n_4031),
.B(n_2204),
.C(n_2500),
.D(n_2499),
.Y(n_4081)
);

AOI22xp33_ASAP7_75t_L g4082 ( 
.A1(n_4061),
.A2(n_4037),
.B1(n_4052),
.B2(n_4048),
.Y(n_4082)
);

OAI211xp5_ASAP7_75t_L g4083 ( 
.A1(n_4062),
.A2(n_4048),
.B(n_4053),
.C(n_4049),
.Y(n_4083)
);

NAND2x1_ASAP7_75t_L g4084 ( 
.A(n_4066),
.B(n_2428),
.Y(n_4084)
);

INVx3_ASAP7_75t_L g4085 ( 
.A(n_4057),
.Y(n_4085)
);

XOR2xp5_ASAP7_75t_L g4086 ( 
.A(n_4056),
.B(n_2143),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4068),
.Y(n_4087)
);

HB1xp67_ASAP7_75t_L g4088 ( 
.A(n_4058),
.Y(n_4088)
);

AOI22xp5_ASAP7_75t_SL g4089 ( 
.A1(n_4079),
.A2(n_2312),
.B1(n_2315),
.B2(n_2325),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_SL g4090 ( 
.A(n_4073),
.B(n_2349),
.Y(n_4090)
);

INVxp67_ASAP7_75t_L g4091 ( 
.A(n_4067),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_4063),
.B(n_2369),
.Y(n_4092)
);

AND2x4_ASAP7_75t_L g4093 ( 
.A(n_4060),
.B(n_2346),
.Y(n_4093)
);

BUFx2_ASAP7_75t_L g4094 ( 
.A(n_4075),
.Y(n_4094)
);

INVx1_ASAP7_75t_SL g4095 ( 
.A(n_4069),
.Y(n_4095)
);

INVxp67_ASAP7_75t_L g4096 ( 
.A(n_4071),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_4059),
.B(n_2369),
.Y(n_4097)
);

AOI221x1_ASAP7_75t_L g4098 ( 
.A1(n_4080),
.A2(n_2226),
.B1(n_2247),
.B2(n_2231),
.C(n_2312),
.Y(n_4098)
);

XNOR2x1_ASAP7_75t_L g4099 ( 
.A(n_4077),
.B(n_2143),
.Y(n_4099)
);

OR2x2_ASAP7_75t_L g4100 ( 
.A(n_4075),
.B(n_4065),
.Y(n_4100)
);

OA22x2_ASAP7_75t_L g4101 ( 
.A1(n_4081),
.A2(n_2328),
.B1(n_2420),
.B2(n_2428),
.Y(n_4101)
);

AOI221x1_ASAP7_75t_L g4102 ( 
.A1(n_4070),
.A2(n_2247),
.B1(n_2325),
.B2(n_2328),
.C(n_2315),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_4072),
.B(n_2369),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_4076),
.B(n_2336),
.Y(n_4104)
);

NOR2x1_ASAP7_75t_L g4105 ( 
.A(n_4085),
.B(n_4064),
.Y(n_4105)
);

NAND4xp25_ASAP7_75t_L g4106 ( 
.A(n_4091),
.B(n_4078),
.C(n_4074),
.D(n_2499),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_4094),
.Y(n_4107)
);

AOI22xp5_ASAP7_75t_L g4108 ( 
.A1(n_4088),
.A2(n_2446),
.B1(n_2433),
.B2(n_2432),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4087),
.B(n_2336),
.Y(n_4109)
);

AO22x2_ASAP7_75t_L g4110 ( 
.A1(n_4095),
.A2(n_2432),
.B1(n_2346),
.B2(n_2333),
.Y(n_4110)
);

XOR2xp5_ASAP7_75t_L g4111 ( 
.A(n_4086),
.B(n_2281),
.Y(n_4111)
);

OAI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_4104),
.A2(n_2306),
.B1(n_2311),
.B2(n_2332),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4100),
.Y(n_4113)
);

OAI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_4090),
.A2(n_2036),
.B(n_2027),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_4083),
.A2(n_2333),
.B1(n_2311),
.B2(n_2050),
.Y(n_4115)
);

OAI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_4082),
.A2(n_2176),
.B1(n_2119),
.B2(n_2117),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_4096),
.B(n_2050),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_4093),
.Y(n_4118)
);

INVx2_ASAP7_75t_SL g4119 ( 
.A(n_4084),
.Y(n_4119)
);

OAI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_4103),
.A2(n_2176),
.B1(n_2119),
.B2(n_2117),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_4093),
.Y(n_4121)
);

INVx1_ASAP7_75t_SL g4122 ( 
.A(n_4099),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4101),
.Y(n_4123)
);

CKINVDCx20_ASAP7_75t_R g4124 ( 
.A(n_4097),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_4092),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4107),
.Y(n_4126)
);

AOI221xp5_ASAP7_75t_L g4127 ( 
.A1(n_4113),
.A2(n_4098),
.B1(n_4102),
.B2(n_4089),
.C(n_2111),
.Y(n_4127)
);

NAND4xp25_ASAP7_75t_L g4128 ( 
.A(n_4105),
.B(n_2035),
.C(n_2137),
.D(n_2145),
.Y(n_4128)
);

NOR2xp67_ASAP7_75t_SL g4129 ( 
.A(n_4118),
.B(n_2281),
.Y(n_4129)
);

AOI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_4122),
.A2(n_4124),
.B1(n_4117),
.B2(n_4106),
.Y(n_4130)
);

AOI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_4123),
.A2(n_2194),
.B1(n_2215),
.B2(n_2110),
.Y(n_4131)
);

AND3x4_ASAP7_75t_L g4132 ( 
.A(n_4121),
.B(n_2284),
.C(n_2191),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4119),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_4111),
.B(n_2194),
.Y(n_4134)
);

AOI221xp5_ASAP7_75t_L g4135 ( 
.A1(n_4112),
.A2(n_2113),
.B1(n_2118),
.B2(n_2110),
.C(n_2111),
.Y(n_4135)
);

OAI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_4109),
.A2(n_2230),
.B(n_2027),
.Y(n_4136)
);

AOI221xp5_ASAP7_75t_L g4137 ( 
.A1(n_4120),
.A2(n_2113),
.B1(n_2118),
.B2(n_2145),
.C(n_2141),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_4125),
.A2(n_2215),
.B(n_2284),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4110),
.Y(n_4139)
);

BUFx2_ASAP7_75t_L g4140 ( 
.A(n_4110),
.Y(n_4140)
);

NOR3xp33_ASAP7_75t_L g4141 ( 
.A(n_4126),
.B(n_4115),
.C(n_4116),
.Y(n_4141)
);

AOI22xp5_ASAP7_75t_L g4142 ( 
.A1(n_4133),
.A2(n_4108),
.B1(n_4114),
.B2(n_2194),
.Y(n_4142)
);

NAND5xp2_ASAP7_75t_L g4143 ( 
.A(n_4130),
.B(n_2336),
.C(n_2137),
.D(n_2141),
.E(n_2035),
.Y(n_4143)
);

NOR3xp33_ASAP7_75t_L g4144 ( 
.A(n_4140),
.B(n_2189),
.C(n_2191),
.Y(n_4144)
);

AOI22xp5_ASAP7_75t_L g4145 ( 
.A1(n_4134),
.A2(n_2215),
.B1(n_2189),
.B2(n_2144),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_4127),
.B(n_2336),
.Y(n_4146)
);

AOI221xp5_ASAP7_75t_L g4147 ( 
.A1(n_4139),
.A2(n_2144),
.B1(n_2405),
.B2(n_2336),
.C(n_2408),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_4132),
.Y(n_4148)
);

OR4x1_ASAP7_75t_L g4149 ( 
.A(n_4129),
.B(n_2408),
.C(n_2405),
.D(n_2336),
.Y(n_4149)
);

NAND5xp2_ASAP7_75t_L g4150 ( 
.A(n_4131),
.B(n_2405),
.C(n_2408),
.D(n_2136),
.E(n_2196),
.Y(n_4150)
);

AOI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_4128),
.A2(n_2136),
.B1(n_2182),
.B2(n_2196),
.Y(n_4151)
);

OAI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_4141),
.A2(n_4138),
.B(n_4136),
.Y(n_4152)
);

AO21x1_ASAP7_75t_L g4153 ( 
.A1(n_4148),
.A2(n_4137),
.B(n_4135),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_SL g4154 ( 
.A(n_4142),
.B(n_4146),
.Y(n_4154)
);

HB1xp67_ASAP7_75t_L g4155 ( 
.A(n_4144),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4143),
.Y(n_4156)
);

OAI22xp5_ASAP7_75t_SL g4157 ( 
.A1(n_4149),
.A2(n_2136),
.B1(n_2182),
.B2(n_2405),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4155),
.Y(n_4158)
);

XNOR2xp5_ASAP7_75t_L g4159 ( 
.A(n_4156),
.B(n_4145),
.Y(n_4159)
);

NOR3xp33_ASAP7_75t_L g4160 ( 
.A(n_4154),
.B(n_4150),
.C(n_4147),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_4152),
.Y(n_4161)
);

OAI22x1_ASAP7_75t_L g4162 ( 
.A1(n_4159),
.A2(n_4153),
.B1(n_4151),
.B2(n_4157),
.Y(n_4162)
);

XOR2xp5_ASAP7_75t_L g4163 ( 
.A(n_4158),
.B(n_2136),
.Y(n_4163)
);

OAI22xp5_ASAP7_75t_L g4164 ( 
.A1(n_4161),
.A2(n_2182),
.B1(n_2408),
.B2(n_2405),
.Y(n_4164)
);

XOR2xp5_ASAP7_75t_L g4165 ( 
.A(n_4162),
.B(n_4163),
.Y(n_4165)
);

AOI22xp5_ASAP7_75t_L g4166 ( 
.A1(n_4164),
.A2(n_4160),
.B1(n_2182),
.B2(n_2126),
.Y(n_4166)
);

AOI21xp33_ASAP7_75t_L g4167 ( 
.A1(n_4165),
.A2(n_2228),
.B(n_2126),
.Y(n_4167)
);

AOI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_4166),
.A2(n_2228),
.B(n_2219),
.Y(n_4168)
);

INVxp67_ASAP7_75t_L g4169 ( 
.A(n_4168),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4167),
.Y(n_4170)
);

OR2x6_ASAP7_75t_L g4171 ( 
.A(n_4170),
.B(n_2201),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_4171),
.A2(n_4169),
.B(n_2219),
.Y(n_4172)
);

AOI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_4172),
.A2(n_2408),
.B1(n_2405),
.B2(n_2201),
.Y(n_4173)
);


endmodule