module fake_jpeg_15243_n_163 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_15),
.B(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_36),
.A2(n_40),
.B1(n_43),
.B2(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_20),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_38),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_3),
.C(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_20),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_6),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_7),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_16),
.A2(n_12),
.B1(n_25),
.B2(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_16),
.B(n_25),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_31),
.C(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_53),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_18),
.Y(n_53)
);

NOR2x1p5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_34),
.B(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_35),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_93),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_62),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_90),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_52),
.A3(n_72),
.B1(n_77),
.B2(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_94),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_79),
.B1(n_65),
.B2(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_67),
.B1(n_54),
.B2(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_101),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_61),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_76),
.C(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_63),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_74),
.C(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_103),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_55),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_120),
.B1(n_102),
.B2(n_101),
.Y(n_125)
);

NAND2xp67_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_91),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_118),
.C(n_113),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_90),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_129),
.C(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_106),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_91),
.B(n_85),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_121),
.B(n_113),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_100),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_98),
.B1(n_94),
.B2(n_99),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_131),
.B1(n_117),
.B2(n_107),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_98),
.B1(n_93),
.B2(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_140),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_115),
.B1(n_108),
.B2(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_104),
.Y(n_141)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_133),
.A3(n_138),
.B1(n_137),
.B2(n_136),
.C1(n_140),
.C2(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

AO221x1_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_144),
.B1(n_128),
.B2(n_132),
.C(n_122),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_108),
.C(n_124),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_126),
.C(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_133),
.C(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_145),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_141),
.B(n_139),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_150),
.B(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_151),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.C(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_152),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_159),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_153),
.B(n_161),
.Y(n_163)
);


endmodule