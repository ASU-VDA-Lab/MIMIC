module fake_netlist_6_2328_n_2452 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_53, n_51, n_44, n_56, n_2452);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2452;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_68;
wire n_726;
wire n_2157;
wire n_2332;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_77;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_78;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_142;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_62;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_65;
wire n_230;
wire n_461;
wire n_873;
wire n_141;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_71;
wire n_229;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_112;
wire n_1280;
wire n_713;
wire n_1400;
wire n_126;
wire n_1467;
wire n_58;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_163;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_2113;
wire n_1641;
wire n_1918;
wire n_2190;
wire n_577;
wire n_166;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_92;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_102;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_121;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_61;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_117;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_134;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_136;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_88;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_170;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_91;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_63;
wire n_362;
wire n_148;
wire n_2279;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_125;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_131;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_59;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_108;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_86;
wire n_104;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_72;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_79;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_147;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_2316;
wire n_1771;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_156;
wire n_145;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_118;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_107;
wire n_1228;
wire n_417;
wire n_446;
wire n_89;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_69;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_98;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_66;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_100;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_124;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_123;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_162;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_128;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_146;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_113;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_90;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_99;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_120;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2181;
wire n_1594;
wire n_1995;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_144;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_106;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_2420;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_140;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_67;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_198;
wire n_1847;
wire n_2052;
wire n_179;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_73;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_101;
wire n_167;
wire n_1356;
wire n_1589;
wire n_127;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_133;
wire n_1320;
wire n_96;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_137;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_122;
wire n_2220;
wire n_1262;
wire n_218;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_70;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_97;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_80;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_2017;
wire n_1682;
wire n_370;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_83;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_105;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_164;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_76;
wire n_548;
wire n_1782;
wire n_94;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_139;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_157;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_138;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_85;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_75;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_151;
wire n_110;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_57;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_84;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_176;
wire n_114;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_74;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_111;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_119;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2284;
wire n_191;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_174;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_129;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_109;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_82;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_93;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_103;
wire n_1693;
wire n_1109;
wire n_185;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_132;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_130;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_116;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_95;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_115;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_158;
wire n_2107;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_87;
wire n_1890;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_207;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_81;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_64;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_135;
wire n_165;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_60;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_40),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_10),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_20),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_18),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_22),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_11),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_28),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_33),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_21),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_43),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_107),
.B1(n_61),
.B2(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_81),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_102),
.B(n_111),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_64),
.B(n_83),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_64),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_93),
.B(n_83),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_119),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_60),
.B(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx6p67_ASAP7_75t_R g162 ( 
.A(n_118),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_99),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_99),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_100),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_100),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_153),
.C(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_136),
.A2(n_107),
.B1(n_101),
.B2(n_112),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_144),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_101),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_145),
.B(n_129),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_145),
.B(n_151),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_144),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_143),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_144),
.B(n_148),
.Y(n_233)
);

NAND2x1_ASAP7_75t_L g234 ( 
.A(n_135),
.B(n_129),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_157),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_142),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_151),
.B(n_132),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_186),
.Y(n_240)
);

OR2x6_ASAP7_75t_L g241 ( 
.A(n_170),
.B(n_143),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_142),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_192),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_170),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

CKINVDCx8_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_202),
.A2(n_233),
.B1(n_204),
.B2(n_165),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_206),
.A2(n_136),
.B1(n_143),
.B2(n_142),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g256 ( 
.A(n_237),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_202),
.B(n_136),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

CKINVDCx11_ASAP7_75t_R g262 ( 
.A(n_196),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_185),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_189),
.B(n_143),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_173),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_186),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_185),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_231),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_218),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_186),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_206),
.A2(n_136),
.B1(n_143),
.B2(n_135),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_212),
.B(n_216),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_185),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_162),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_212),
.B(n_143),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_203),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_165),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_167),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_206),
.A2(n_116),
.B1(n_112),
.B2(n_66),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_167),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_235),
.B(n_143),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_203),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_203),
.B(n_162),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_233),
.A2(n_135),
.B1(n_162),
.B2(n_148),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_185),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_132),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_168),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_185),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_168),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_168),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_190),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_233),
.B(n_60),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_219),
.B(n_208),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_185),
.B(n_138),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_219),
.B(n_162),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_185),
.B(n_68),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_208),
.B(n_162),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_208),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_208),
.B(n_162),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_204),
.B(n_147),
.C(n_153),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_194),
.B(n_195),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_194),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_208),
.B(n_162),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_167),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_135),
.B1(n_148),
.B2(n_138),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_190),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_208),
.B(n_135),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_234),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_169),
.B(n_135),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_194),
.B(n_68),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_220),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_234),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_169),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_220),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_169),
.B(n_135),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_204),
.B(n_65),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_171),
.A2(n_135),
.B1(n_77),
.B2(n_147),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_171),
.B(n_65),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_238),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_194),
.B(n_69),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_171),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_175),
.B(n_178),
.C(n_176),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_175),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_175),
.B(n_135),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_176),
.B(n_116),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_176),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_178),
.B(n_69),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_178),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_238),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_182),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_194),
.B(n_71),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_182),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_182),
.A2(n_191),
.B1(n_197),
.B2(n_230),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_184),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_184),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_184),
.B(n_187),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_187),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_187),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_194),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_188),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_194),
.B(n_71),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_188),
.B(n_135),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_188),
.B(n_62),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_191),
.B(n_135),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_191),
.Y(n_368)
);

OR2x6_ASAP7_75t_L g369 ( 
.A(n_196),
.B(n_148),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_197),
.B(n_63),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_244),
.B(n_194),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_256),
.B(n_197),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_258),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_258),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_243),
.B(n_205),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_248),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_244),
.B(n_194),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_248),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_244),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_244),
.B(n_195),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_205),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_244),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_240),
.B(n_205),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_311),
.B(n_209),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_209),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_247),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_263),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_240),
.B(n_209),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_289),
.B(n_211),
.Y(n_390)
);

NOR3x1_ASAP7_75t_L g391 ( 
.A(n_304),
.B(n_104),
.C(n_87),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_247),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_268),
.B(n_270),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_263),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_249),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_251),
.B(n_211),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_249),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_259),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_244),
.B(n_195),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_257),
.B(n_195),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_L g401 ( 
.A(n_345),
.B(n_214),
.C(n_215),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_257),
.B(n_277),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_268),
.B(n_211),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_259),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_257),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_282),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_270),
.B(n_214),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_264),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_264),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_257),
.B(n_195),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_272),
.B(n_214),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_304),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_271),
.B(n_215),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_260),
.A2(n_228),
.B1(n_215),
.B2(n_230),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_271),
.B(n_217),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_254),
.B(n_246),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_283),
.B(n_255),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_305),
.B(n_217),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_260),
.A2(n_196),
.B1(n_230),
.B2(n_217),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_L g421 ( 
.A(n_257),
.B(n_195),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_305),
.B(n_228),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_272),
.B(n_228),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_260),
.A2(n_196),
.B1(n_234),
.B2(n_179),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_307),
.B(n_195),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_257),
.B(n_195),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_277),
.B(n_195),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_295),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_273),
.B(n_196),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_248),
.B(n_195),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_307),
.B(n_210),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_267),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_267),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_295),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_281),
.B(n_210),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_310),
.A2(n_275),
.B1(n_276),
.B2(n_273),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_308),
.B(n_210),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_308),
.B(n_210),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_266),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_274),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_274),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_310),
.A2(n_196),
.B1(n_172),
.B2(n_179),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_275),
.A2(n_148),
.B(n_229),
.C(n_224),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_338),
.Y(n_447)
);

AND2x4_ASAP7_75t_SL g448 ( 
.A(n_277),
.B(n_210),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_309),
.B(n_210),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_281),
.B(n_210),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_279),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_277),
.B(n_210),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_266),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_296),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_277),
.B(n_210),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_281),
.B(n_210),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_276),
.B(n_213),
.Y(n_457)
);

O2A1O1Ixp5_ASAP7_75t_L g458 ( 
.A1(n_314),
.A2(n_153),
.B(n_147),
.C(n_137),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_266),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_299),
.B(n_213),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_279),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_338),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_277),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_250),
.B(n_72),
.Y(n_464)
);

AND2x6_ASAP7_75t_SL g465 ( 
.A(n_296),
.B(n_75),
.Y(n_465)
);

AOI22x1_ASAP7_75t_L g466 ( 
.A1(n_309),
.A2(n_330),
.B1(n_322),
.B2(n_325),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_322),
.B(n_213),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_287),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_325),
.B(n_330),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_294),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_287),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_336),
.B(n_213),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_331),
.B(n_213),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_294),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_331),
.B(n_213),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_293),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_293),
.Y(n_477)
);

AOI221xp5_ASAP7_75t_L g478 ( 
.A1(n_285),
.A2(n_70),
.B1(n_67),
.B2(n_66),
.C(n_102),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_300),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_334),
.B(n_213),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_300),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_269),
.B(n_213),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_316),
.Y(n_483)
);

NOR3xp33_ASAP7_75t_L g484 ( 
.A(n_292),
.B(n_105),
.C(n_84),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_294),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_252),
.B(n_213),
.C(n_229),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_284),
.B(n_213),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_284),
.B(n_224),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_286),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_336),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_316),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_334),
.B(n_224),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_286),
.A2(n_321),
.B1(n_333),
.B2(n_350),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_369),
.B(n_172),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_297),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_265),
.B(n_224),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_318),
.B(n_153),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_261),
.B(n_224),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_297),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_297),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_369),
.B(n_172),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_373),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_373),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_374),
.Y(n_505)
);

OR2x2_ASAP7_75t_SL g506 ( 
.A(n_465),
.B(n_75),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_390),
.B(n_381),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_375),
.B(n_310),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_442),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_379),
.B(n_382),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_396),
.B(n_339),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_376),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_374),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_383),
.B(n_339),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_393),
.B(n_350),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_453),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_469),
.B(n_372),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_369),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_460),
.B(n_351),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_388),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_418),
.A2(n_285),
.B1(n_262),
.B2(n_370),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_453),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_379),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_241),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_406),
.B(n_351),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_383),
.B(n_347),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_490),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_482),
.B(n_359),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_494),
.B(n_369),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_459),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_388),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_376),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_463),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_447),
.A2(n_366),
.B1(n_337),
.B2(n_318),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_394),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_386),
.A2(n_340),
.B1(n_329),
.B2(n_353),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_498),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_489),
.B(n_291),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_386),
.A2(n_364),
.B1(n_369),
.B2(n_346),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_459),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_463),
.B(n_265),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_378),
.B(n_265),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_489),
.B(n_341),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_386),
.A2(n_368),
.B1(n_346),
.B2(n_348),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_SL g552 ( 
.A(n_478),
.B(n_70),
.C(n_67),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_500),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_470),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_470),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_241),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_470),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_464),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_378),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_386),
.Y(n_563)
);

NOR2x2_ASAP7_75t_L g564 ( 
.A(n_454),
.B(n_241),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_489),
.B(n_341),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_462),
.B(n_343),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_429),
.B(n_348),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_384),
.B(n_265),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_384),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_474),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_389),
.B(n_352),
.Y(n_571)
);

BUFx4f_ASAP7_75t_SL g572 ( 
.A(n_501),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

AO21x1_ASAP7_75t_L g574 ( 
.A1(n_493),
.A2(n_306),
.B(n_298),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_385),
.B(n_343),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_485),
.Y(n_577)
);

BUFx12f_ASAP7_75t_SL g578 ( 
.A(n_501),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_414),
.B(n_438),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_421),
.A2(n_362),
.B(n_303),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_429),
.B(n_352),
.Y(n_581)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_501),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_452),
.B(n_302),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_499),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_SL g586 ( 
.A(n_484),
.B(n_250),
.C(n_78),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_379),
.B(n_354),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_465),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_499),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_387),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_411),
.B(n_354),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_411),
.B(n_358),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_415),
.B(n_280),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_423),
.B(n_358),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_423),
.B(n_368),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_448),
.B(n_298),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_448),
.B(n_298),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_457),
.B(n_360),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_391),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_415),
.B(n_360),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_428),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_420),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_387),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_387),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_379),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_379),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_495),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_392),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_392),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_392),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_395),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_391),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_395),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_382),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_457),
.B(n_245),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_395),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_428),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_420),
.A2(n_357),
.B1(n_323),
.B2(n_361),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_404),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_486),
.A2(n_337),
.B1(n_241),
.B2(n_356),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_435),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_487),
.B(n_323),
.Y(n_625)
);

AND3x1_ASAP7_75t_SL g626 ( 
.A(n_435),
.B(n_91),
.C(n_110),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_404),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_487),
.B(n_298),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_SL g629 ( 
.A(n_401),
.B(n_106),
.C(n_79),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_488),
.B(n_306),
.Y(n_630)
);

OR2x2_ASAP7_75t_SL g631 ( 
.A(n_486),
.B(n_76),
.Y(n_631)
);

BUFx2_ASAP7_75t_SL g632 ( 
.A(n_382),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_404),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_434),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_398),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_434),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_398),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_488),
.B(n_306),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_397),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_497),
.B(n_306),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_408),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_497),
.B(n_320),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_397),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_440),
.B(n_323),
.Y(n_644)
);

NOR2x2_ASAP7_75t_L g645 ( 
.A(n_434),
.B(n_241),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_448),
.B(n_320),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_445),
.B(n_327),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_403),
.B(n_320),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_445),
.B(n_323),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_L g650 ( 
.A(n_424),
.B(n_342),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_440),
.A2(n_357),
.B1(n_361),
.B2(n_342),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_382),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_437),
.B(n_357),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_432),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_407),
.B(n_320),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_408),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_409),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_409),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_443),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_413),
.B(n_416),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_617),
.B(n_382),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_507),
.B(n_419),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_524),
.B(n_355),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_530),
.B(n_355),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_530),
.B(n_355),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_521),
.B(n_422),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_542),
.B(n_561),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_514),
.B(n_355),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_604),
.B(n_437),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_604),
.B(n_437),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_509),
.B(n_532),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_SL g672 ( 
.A(n_602),
.B(n_319),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_582),
.B(n_303),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_582),
.B(n_303),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_598),
.B(n_424),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_563),
.B(n_303),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_563),
.B(n_303),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_526),
.B(n_303),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_516),
.B(n_537),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_SL g680 ( 
.A(n_552),
.B(n_405),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_516),
.B(n_362),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_537),
.B(n_550),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_SL g683 ( 
.A(n_519),
.B(n_405),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_518),
.B(n_660),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_647),
.B(n_362),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_647),
.B(n_362),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_647),
.B(n_362),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_647),
.B(n_362),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_518),
.B(n_472),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_569),
.B(n_430),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_629),
.B(n_405),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_569),
.B(n_436),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_504),
.B(n_450),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_504),
.B(n_456),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_504),
.B(n_405),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_583),
.B(n_472),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_583),
.B(n_466),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_SL g698 ( 
.A(n_649),
.B(n_425),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_583),
.B(n_466),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_566),
.B(n_290),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_SL g701 ( 
.A(n_523),
.B(n_371),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_531),
.B(n_290),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_649),
.B(n_290),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_539),
.B(n_290),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_539),
.B(n_290),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_598),
.B(n_357),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_SL g707 ( 
.A(n_597),
.B(n_377),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_588),
.B(n_361),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_533),
.B(n_431),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_588),
.B(n_361),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_594),
.B(n_401),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_567),
.B(n_439),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_SL g713 ( 
.A(n_601),
.B(n_441),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_572),
.B(n_443),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_621),
.B(n_444),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_SL g716 ( 
.A(n_615),
.B(n_449),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_579),
.B(n_444),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_567),
.B(n_467),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_581),
.B(n_461),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_599),
.B(n_473),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_581),
.B(n_461),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_SL g722 ( 
.A(n_646),
.B(n_475),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_625),
.B(n_650),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_522),
.B(n_72),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_625),
.B(n_468),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_650),
.B(n_468),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_522),
.B(n_471),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_522),
.B(n_471),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_522),
.B(n_479),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_534),
.B(n_479),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_SL g731 ( 
.A(n_528),
.B(n_480),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_534),
.B(n_481),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_534),
.B(n_481),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_534),
.B(n_483),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_528),
.B(n_492),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_562),
.B(n_483),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_571),
.B(n_491),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_620),
.B(n_72),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_491),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_562),
.B(n_432),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_543),
.B(n_433),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_576),
.B(n_433),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_617),
.B(n_451),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_SL g744 ( 
.A(n_528),
.B(n_380),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_529),
.B(n_451),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_529),
.B(n_476),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_617),
.B(n_476),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_617),
.B(n_477),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_617),
.B(n_477),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_SL g750 ( 
.A(n_528),
.B(n_399),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_592),
.B(n_446),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_617),
.B(n_242),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_651),
.B(n_242),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_529),
.B(n_558),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_541),
.B(n_242),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_SL g756 ( 
.A(n_603),
.B(n_400),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_603),
.B(n_72),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_644),
.B(n_242),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_551),
.B(n_253),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_640),
.B(n_253),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_529),
.B(n_402),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_642),
.B(n_508),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_508),
.B(n_538),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_508),
.B(n_253),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_628),
.B(n_410),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_624),
.B(n_72),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_SL g767 ( 
.A(n_630),
.B(n_426),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_538),
.B(n_253),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_538),
.B(n_278),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_624),
.B(n_278),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_502),
.B(n_278),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_502),
.B(n_278),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_503),
.B(n_288),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_503),
.B(n_288),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_505),
.B(n_288),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_SL g776 ( 
.A(n_638),
.B(n_427),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_593),
.B(n_455),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_595),
.B(n_328),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_505),
.B(n_288),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_596),
.B(n_335),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_517),
.B(n_327),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_517),
.B(n_327),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_525),
.B(n_327),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_586),
.B(n_74),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_525),
.B(n_332),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_536),
.B(n_344),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_536),
.B(n_332),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_540),
.B(n_545),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_540),
.B(n_545),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_SL g790 ( 
.A(n_600),
.B(n_496),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_618),
.B(n_365),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_549),
.B(n_332),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_565),
.B(n_332),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_SL g794 ( 
.A(n_648),
.B(n_655),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_544),
.B(n_224),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_653),
.B(n_224),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_635),
.B(n_367),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_SL g798 ( 
.A(n_635),
.B(n_301),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_637),
.B(n_224),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_637),
.B(n_224),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_641),
.B(n_224),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_641),
.B(n_324),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_SL g803 ( 
.A(n_656),
.B(n_315),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_656),
.B(n_229),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_657),
.B(n_229),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_SL g806 ( 
.A(n_657),
.B(n_317),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_658),
.B(n_229),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_658),
.B(n_229),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_659),
.B(n_229),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_634),
.B(n_229),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_SL g811 ( 
.A(n_634),
.B(n_229),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_659),
.B(n_229),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_547),
.B(n_458),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_553),
.B(n_312),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_547),
.B(n_86),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_547),
.B(n_88),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_553),
.B(n_89),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_554),
.B(n_90),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_SL g819 ( 
.A(n_636),
.B(n_326),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_554),
.B(n_92),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_623),
.B(n_96),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_623),
.B(n_97),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_568),
.B(n_103),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_636),
.B(n_108),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_639),
.B(n_113),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_639),
.B(n_85),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_643),
.B(n_85),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_SL g828 ( 
.A(n_608),
.B(n_312),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_643),
.B(n_85),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_654),
.B(n_85),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_654),
.B(n_85),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_605),
.B(n_172),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_SL g833 ( 
.A(n_608),
.B(n_312),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_591),
.B(n_312),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_591),
.B(n_312),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_SL g836 ( 
.A(n_608),
.B(n_609),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_605),
.B(n_172),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_SL g838 ( 
.A(n_645),
.B(n_76),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_SL g839 ( 
.A(n_609),
.B(n_80),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_609),
.B(n_80),
.Y(n_840)
);

BUFx4f_ASAP7_75t_L g841 ( 
.A(n_661),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_684),
.B(n_610),
.Y(n_842)
);

XNOR2x1_ASAP7_75t_L g843 ( 
.A(n_738),
.B(n_506),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_675),
.B(n_529),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_788),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_789),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_745),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_737),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_757),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_711),
.B(n_666),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_667),
.Y(n_851)
);

NAND2x1_ASAP7_75t_L g852 ( 
.A(n_745),
.B(n_513),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_766),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_745),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_746),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_662),
.B(n_610),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_739),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_671),
.B(n_669),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_682),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_784),
.A2(n_626),
.B1(n_558),
.B2(n_587),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_696),
.B(n_631),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_661),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_679),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_670),
.B(n_613),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_SL g865 ( 
.A(n_709),
.B(n_632),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_746),
.Y(n_866)
);

BUFx12f_ASAP7_75t_L g867 ( 
.A(n_724),
.Y(n_867)
);

BUFx12f_ASAP7_75t_L g868 ( 
.A(n_746),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_675),
.B(n_558),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_719),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_675),
.B(n_558),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_721),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_821),
.A2(n_558),
.B1(n_578),
.B2(n_574),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_838),
.B(n_606),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_742),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_736),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_754),
.B(n_606),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_802),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_708),
.A2(n_506),
.B1(n_631),
.B2(n_580),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_689),
.B(n_613),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_754),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_786),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_740),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_712),
.B(n_614),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_754),
.B(n_607),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_797),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_761),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_710),
.B(n_607),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_761),
.B(n_611),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_761),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_727),
.B(n_652),
.Y(n_892)
);

AOI221x1_ASAP7_75t_L g893 ( 
.A1(n_701),
.A2(n_574),
.B1(n_612),
.B2(n_611),
.C(n_616),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_728),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_718),
.B(n_614),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_SL g896 ( 
.A1(n_751),
.A2(n_104),
.B1(n_98),
.B2(n_110),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_723),
.B(n_612),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_678),
.A2(n_587),
.B1(n_548),
.B2(n_622),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_680),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_729),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_777),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_817),
.B(n_818),
.Y(n_902)
);

CKINVDCx11_ASAP7_75t_R g903 ( 
.A(n_691),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_730),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_732),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_714),
.B(n_616),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_771),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_772),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_820),
.B(n_652),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_693),
.A2(n_632),
.B1(n_619),
.B2(n_622),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_822),
.B(n_619),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_695),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_698),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_703),
.B(n_627),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_773),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_685),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_733),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_824),
.A2(n_587),
.B1(n_172),
.B2(n_179),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_704),
.B(n_652),
.Y(n_919)
);

AND3x1_ASAP7_75t_SL g920 ( 
.A(n_713),
.B(n_109),
.C(n_98),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_774),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_734),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_705),
.B(n_555),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_775),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_825),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_694),
.A2(n_559),
.B1(n_575),
.B2(n_555),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_725),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_763),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_815),
.B(n_627),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_672),
.A2(n_564),
.B(n_557),
.C(n_559),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_716),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_770),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_779),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_816),
.Y(n_934)
);

INVxp33_ASAP7_75t_L g935 ( 
.A(n_826),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_SL g936 ( 
.A1(n_791),
.A2(n_587),
.B1(n_513),
.B2(n_91),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_697),
.B(n_633),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_717),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_726),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_672),
.A2(n_556),
.B(n_570),
.C(n_557),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_834),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_699),
.B(n_633),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_778),
.B(n_510),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_814),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_836),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_686),
.B(n_556),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_687),
.B(n_560),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_781),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_688),
.B(n_560),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_827),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_690),
.B(n_570),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_796),
.A2(n_795),
.B1(n_664),
.B2(n_665),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_764),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_663),
.B(n_575),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_829),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_835),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_830),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_706),
.B(n_577),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_756),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_782),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_692),
.B(n_577),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_831),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_783),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_673),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_785),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_674),
.B(n_584),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_787),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_780),
.B(n_510),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_681),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_823),
.B(n_511),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_762),
.B(n_511),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_715),
.B(n_512),
.Y(n_973)
);

AOI21xp33_ASAP7_75t_L g974 ( 
.A1(n_755),
.A2(n_584),
.B(n_589),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_702),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_794),
.B(n_512),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_794),
.B(n_515),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_813),
.B(n_590),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_769),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_792),
.B(n_515),
.Y(n_980)
);

NAND3xp33_ASAP7_75t_SL g981 ( 
.A(n_701),
.B(n_109),
.C(n_94),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_799),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_790),
.B(n_765),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_743),
.B(n_520),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_839),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_790),
.B(n_520),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_832),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_800),
.B(n_527),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_801),
.B(n_527),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_836),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_804),
.Y(n_991)
);

AND3x1_ASAP7_75t_SL g992 ( 
.A(n_840),
.B(n_94),
.C(n_87),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_793),
.B(n_535),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_805),
.B(n_535),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_747),
.B(n_546),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_810),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_837),
.B(n_546),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_828),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_700),
.B(n_578),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_807),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_748),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_753),
.B(n_573),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_749),
.B(n_573),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_744),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_R g1005 ( 
.A(n_707),
.B(n_513),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_668),
.B(n_585),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_808),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_765),
.A2(n_82),
.B(n_589),
.C(n_585),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_809),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_978),
.A2(n_760),
.B(n_812),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_868),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_864),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_850),
.B(n_590),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_981),
.A2(n_683),
.B(n_776),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_978),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_978),
.A2(n_676),
.B(n_677),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_878),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_868),
.Y(n_1018)
);

BUFx12f_ASAP7_75t_L g1019 ( 
.A(n_849),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_983),
.A2(n_776),
.B(n_767),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_998),
.A2(n_752),
.B(n_758),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_848),
.B(n_857),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_998),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_851),
.B(n_853),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_945),
.Y(n_1025)
);

INVx6_ASAP7_75t_L g1026 ( 
.A(n_888),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_878),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_937),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_951),
.Y(n_1029)
);

BUFx4f_ASAP7_75t_L g1030 ( 
.A(n_919),
.Y(n_1030)
);

AO21x2_ASAP7_75t_L g1031 ( 
.A1(n_940),
.A2(n_759),
.B(n_148),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_893),
.A2(n_148),
.B(n_137),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_851),
.B(n_82),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_886),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_998),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_891),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_951),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_945),
.Y(n_1038)
);

OR2x6_ASAP7_75t_L g1039 ( 
.A(n_913),
.B(n_828),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_945),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_896),
.A2(n_767),
.B1(n_707),
.B2(n_722),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_937),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_886),
.Y(n_1043)
);

BUFx12f_ASAP7_75t_L g1044 ( 
.A(n_849),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_986),
.A2(n_803),
.B(n_798),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_962),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_891),
.B(n_513),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_890),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_882),
.Y(n_1049)
);

BUFx2_ASAP7_75t_R g1050 ( 
.A(n_863),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_990),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_852),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_962),
.Y(n_1053)
);

AO21x2_ASAP7_75t_L g1054 ( 
.A1(n_930),
.A2(n_806),
.B(n_798),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_890),
.B(n_844),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_990),
.A2(n_811),
.B(n_810),
.Y(n_1056)
);

INVx2_ASAP7_75t_R g1057 ( 
.A(n_1004),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_902),
.A2(n_806),
.B(n_803),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_882),
.B(n_513),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_882),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_865),
.A2(n_137),
.B(n_138),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_990),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_976),
.A2(n_138),
.B(n_819),
.Y(n_1063)
);

CKINVDCx14_ASAP7_75t_R g1064 ( 
.A(n_859),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_977),
.A2(n_819),
.B(n_833),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_1008),
.A2(n_137),
.B(n_735),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_858),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_893),
.A2(n_941),
.B(n_852),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_958),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_913),
.B(n_865),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_941),
.A2(n_833),
.B(n_731),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_879),
.B(n_720),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_1009),
.A2(n_161),
.B(n_158),
.Y(n_1073)
);

AOI21x1_ASAP7_75t_L g1074 ( 
.A1(n_880),
.A2(n_889),
.B(n_960),
.Y(n_1074)
);

AO21x2_ASAP7_75t_L g1075 ( 
.A1(n_974),
.A2(n_811),
.B(n_750),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_888),
.B(n_513),
.Y(n_1076)
);

BUFx10_ASAP7_75t_L g1077 ( 
.A(n_931),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_941),
.A2(n_181),
.B(n_166),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_859),
.Y(n_1079)
);

BUFx4f_ASAP7_75t_L g1080 ( 
.A(n_919),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_1004),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_942),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_888),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_854),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_944),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_923),
.A2(n_181),
.B(n_166),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_923),
.A2(n_181),
.B(n_166),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_931),
.B(n_158),
.Y(n_1088)
);

BUFx12f_ASAP7_75t_L g1089 ( 
.A(n_958),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_935),
.B(n_53),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_942),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_923),
.A2(n_181),
.B(n_166),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_919),
.A2(n_193),
.B(n_177),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_879),
.B(n_587),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_996),
.B(n_587),
.Y(n_1095)
);

AOI22x1_ASAP7_75t_L g1096 ( 
.A1(n_960),
.A2(n_587),
.B1(n_513),
.B2(n_158),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_952),
.A2(n_158),
.B(n_161),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_872),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_844),
.B(n_158),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_944),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_841),
.A2(n_312),
.B(n_161),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_854),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_883),
.B(n_161),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1006),
.A2(n_193),
.B(n_236),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_847),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_901),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_916),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_863),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_847),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_947),
.A2(n_193),
.B(n_236),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_947),
.A2(n_193),
.B(n_236),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_843),
.A2(n_312),
.B1(n_161),
.B2(n_172),
.Y(n_1112)
);

INVxp67_ASAP7_75t_SL g1113 ( 
.A(n_883),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_935),
.B(n_0),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_947),
.Y(n_1115)
);

BUFx2_ASAP7_75t_SL g1116 ( 
.A(n_909),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_980),
.A2(n_236),
.B(n_226),
.Y(n_1117)
);

AOI22x1_ASAP7_75t_L g1118 ( 
.A1(n_887),
.A2(n_151),
.B1(n_154),
.B2(n_179),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_956),
.Y(n_1119)
);

BUFx2_ASAP7_75t_SL g1120 ( 
.A(n_899),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_916),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_867),
.B(n_151),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_872),
.Y(n_1123)
);

BUFx2_ASAP7_75t_SL g1124 ( 
.A(n_899),
.Y(n_1124)
);

AOI22x1_ASAP7_75t_L g1125 ( 
.A1(n_887),
.A2(n_154),
.B1(n_179),
.B2(n_223),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_1005),
.A2(n_154),
.B(n_225),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_916),
.Y(n_1127)
);

AO21x2_ASAP7_75t_L g1128 ( 
.A1(n_1009),
.A2(n_154),
.B(n_225),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_993),
.A2(n_226),
.B(n_225),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_901),
.Y(n_1130)
);

AO21x2_ASAP7_75t_L g1131 ( 
.A1(n_898),
.A2(n_154),
.B(n_225),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_897),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_869),
.B(n_0),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1002),
.A2(n_174),
.B(n_223),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_956),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_897),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_869),
.B(n_871),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_938),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_996),
.B(n_226),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_841),
.Y(n_1140)
);

AOI22x1_ASAP7_75t_L g1141 ( 
.A1(n_876),
.A2(n_179),
.B1(n_223),
.B2(n_221),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_950),
.B(n_1),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_855),
.Y(n_1143)
);

NAND2x1p5_ASAP7_75t_L g1144 ( 
.A(n_841),
.B(n_916),
.Y(n_1144)
);

BUFx12f_ASAP7_75t_L g1145 ( 
.A(n_867),
.Y(n_1145)
);

BUFx2_ASAP7_75t_R g1146 ( 
.A(n_985),
.Y(n_1146)
);

INVx3_ASAP7_75t_SL g1147 ( 
.A(n_985),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_988),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_988),
.Y(n_1149)
);

OR3x4_ASAP7_75t_SL g1150 ( 
.A(n_843),
.B(n_1),
.C(n_2),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_926),
.A2(n_174),
.B(n_223),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_871),
.B(n_3),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1142),
.A2(n_950),
.B1(n_955),
.B2(n_963),
.Y(n_1153)
);

CKINVDCx11_ASAP7_75t_R g1154 ( 
.A(n_1150),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1041),
.A2(n_955),
.B1(n_963),
.B2(n_934),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1019),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1028),
.Y(n_1157)
);

BUFx12f_ASAP7_75t_L g1158 ( 
.A(n_1145),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1108),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1081),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1028),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1138),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1033),
.A2(n_934),
.B1(n_925),
.B2(n_861),
.Y(n_1163)
);

BUFx8_ASAP7_75t_L g1164 ( 
.A(n_1019),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1079),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1081),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1058),
.A2(n_861),
.B1(n_925),
.B2(n_965),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1114),
.A2(n_916),
.B1(n_860),
.B2(n_903),
.Y(n_1168)
);

BUFx12f_ASAP7_75t_L g1169 ( 
.A(n_1145),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1019),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1020),
.A2(n_965),
.B1(n_970),
.B2(n_999),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1028),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1138),
.Y(n_1173)
);

CKINVDCx11_ASAP7_75t_R g1174 ( 
.A(n_1147),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1044),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1122),
.A2(n_965),
.B1(n_970),
.B2(n_922),
.Y(n_1176)
);

OAI21xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1140),
.A2(n_939),
.B(n_906),
.Y(n_1177)
);

BUFx4_ASAP7_75t_SL g1178 ( 
.A(n_1011),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1044),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1090),
.A2(n_1152),
.B1(n_1133),
.B2(n_1112),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1069),
.A2(n_965),
.B1(n_970),
.B2(n_911),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1133),
.A2(n_903),
.B1(n_965),
.B2(n_970),
.Y(n_1182)
);

BUFx8_ASAP7_75t_SL g1183 ( 
.A(n_1069),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_1145),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1152),
.A2(n_970),
.B1(n_874),
.B2(n_855),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1069),
.A2(n_911),
.B1(n_917),
.B2(n_904),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1148),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1064),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1042),
.B(n_866),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1042),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1067),
.B(n_866),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1101),
.A2(n_936),
.B(n_856),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1148),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1147),
.Y(n_1194)
);

INVx6_ASAP7_75t_L g1195 ( 
.A(n_1081),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1067),
.B(n_845),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1044),
.A2(n_929),
.B1(n_987),
.B2(n_900),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1089),
.A2(n_894),
.B1(n_905),
.B2(n_927),
.Y(n_1198)
);

INVx6_ASAP7_75t_L g1199 ( 
.A(n_1081),
.Y(n_1199)
);

INVx6_ASAP7_75t_L g1200 ( 
.A(n_1081),
.Y(n_1200)
);

BUFx8_ASAP7_75t_SL g1201 ( 
.A(n_1089),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1042),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1107),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1089),
.A2(n_892),
.B1(n_932),
.B2(n_875),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1081),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1079),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_SL g1207 ( 
.A(n_1147),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1120),
.A2(n_892),
.B1(n_959),
.B2(n_846),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1107),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1098),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1095),
.Y(n_1211)
);

INVx6_ASAP7_75t_L g1212 ( 
.A(n_1140),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1050),
.A2(n_975),
.B1(n_870),
.B2(n_873),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1012),
.B(n_928),
.Y(n_1214)
);

INVx6_ASAP7_75t_L g1215 ( 
.A(n_1140),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1149),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1120),
.A2(n_892),
.B1(n_959),
.B2(n_877),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1124),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1132),
.B(n_946),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1098),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1124),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1107),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1024),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1077),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1070),
.A2(n_884),
.B1(n_979),
.B2(n_948),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1146),
.A2(n_912),
.B1(n_1001),
.B2(n_968),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1011),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1149),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1099),
.A2(n_959),
.B1(n_966),
.B2(n_964),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1122),
.A2(n_918),
.B1(n_842),
.B2(n_971),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1039),
.A2(n_961),
.B1(n_933),
.B2(n_924),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1070),
.A2(n_914),
.B1(n_1007),
.B2(n_1000),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1014),
.A2(n_910),
.B1(n_920),
.B2(n_967),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1052),
.Y(n_1234)
);

INVx8_ASAP7_75t_L g1235 ( 
.A(n_1038),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1052),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1011),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1039),
.A2(n_924),
.B1(n_915),
.B2(n_933),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1099),
.A2(n_967),
.B1(n_921),
.B2(n_908),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1029),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1029),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1039),
.A2(n_967),
.B1(n_921),
.B2(n_908),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1052),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1070),
.A2(n_914),
.B1(n_991),
.B2(n_1000),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1039),
.A2(n_1018),
.B1(n_1137),
.B2(n_1095),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1018),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1077),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1098),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1018),
.A2(n_992),
.B1(n_954),
.B2(n_907),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1107),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1054),
.A2(n_946),
.B1(n_949),
.B2(n_915),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1123),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1123),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1077),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1123),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1077),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1095),
.A2(n_1144),
.B1(n_1039),
.B2(n_1088),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1107),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1113),
.B(n_949),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_SL g1260 ( 
.A(n_1140),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1037),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1038),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1137),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1055),
.B(n_953),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1084),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1137),
.A2(n_907),
.B1(n_957),
.B2(n_953),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1052),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_SL g1268 ( 
.A(n_1076),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1038),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1054),
.A2(n_957),
.B1(n_862),
.B2(n_1007),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1037),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1095),
.A2(n_881),
.B1(n_973),
.B2(n_969),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1038),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1107),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1046),
.Y(n_1275)
);

BUFx8_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1054),
.A2(n_862),
.B1(n_991),
.B2(n_982),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1116),
.A2(n_862),
.B1(n_995),
.B2(n_984),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1046),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1038),
.B(n_982),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1137),
.A2(n_995),
.B1(n_984),
.B2(n_895),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1072),
.A2(n_972),
.B1(n_994),
.B2(n_885),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1121),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1034),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1265),
.B(n_1053),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1214),
.B(n_1053),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1238),
.A2(n_1063),
.B(n_1061),
.Y(n_1287)
);

OAI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1155),
.A2(n_1022),
.B1(n_1116),
.B2(n_1144),
.C(n_1074),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1157),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1157),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1164),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1161),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1231),
.A2(n_1063),
.B(n_1061),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1162),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1173),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1192),
.A2(n_1056),
.B(n_1272),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1172),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1177),
.A2(n_1045),
.B(n_1030),
.C(n_1080),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1232),
.A2(n_1074),
.B(n_1068),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1263),
.B(n_1057),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1240),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1245),
.A2(n_1068),
.B(n_1045),
.Y(n_1303)
);

AOI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1213),
.A2(n_1013),
.B(n_1032),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1233),
.A2(n_1080),
.B(n_1030),
.C(n_1038),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1165),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1168),
.A2(n_1065),
.B(n_1071),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1172),
.B(n_1057),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1190),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1241),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1280),
.A2(n_1065),
.B(n_1117),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1190),
.Y(n_1312)
);

AOI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1282),
.A2(n_1060),
.B(n_1049),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1230),
.A2(n_1080),
.B(n_1030),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1164),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1154),
.A2(n_1097),
.B1(n_1031),
.B2(n_1066),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1225),
.A2(n_1080),
.B(n_1030),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1261),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1211),
.A2(n_1095),
.B(n_1096),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1202),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1154),
.A2(n_1097),
.B1(n_1031),
.B2(n_1066),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1171),
.A2(n_1071),
.B(n_1040),
.C(n_1051),
.Y(n_1322)
);

INVx8_ASAP7_75t_L g1323 ( 
.A(n_1158),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1271),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1235),
.B(n_1025),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1202),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1275),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1195),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1284),
.B(n_1136),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1279),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1187),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1219),
.B(n_1057),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1207),
.A2(n_1025),
.B1(n_1062),
.B2(n_1144),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1196),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1167),
.A2(n_1051),
.B(n_1040),
.C(n_1135),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1211),
.A2(n_1235),
.B(n_1096),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1211),
.B(n_1132),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1164),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1191),
.B(n_1136),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1247),
.B(n_1121),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1211),
.A2(n_1097),
.B(n_1075),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1264),
.B(n_1132),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1211),
.A2(n_1235),
.B(n_1097),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1163),
.A2(n_1062),
.B1(n_1025),
.B2(n_1026),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1235),
.A2(n_1075),
.B(n_1032),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1259),
.B(n_1193),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1234),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1273),
.B(n_1025),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1242),
.A2(n_1117),
.B(n_1129),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1280),
.A2(n_1129),
.B(n_1134),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1218),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1216),
.B(n_1082),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1210),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1228),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1204),
.A2(n_1104),
.B(n_1134),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1180),
.A2(n_1031),
.B1(n_1066),
.B2(n_1048),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1189),
.B(n_1219),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1244),
.A2(n_1015),
.B(n_1128),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1174),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1210),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1234),
.B(n_1015),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1234),
.B(n_1015),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1257),
.A2(n_1075),
.B(n_1032),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1186),
.B(n_1121),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1278),
.A2(n_1128),
.B(n_1131),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1220),
.Y(n_1366)
);

NAND2x1_ASAP7_75t_L g1367 ( 
.A(n_1273),
.B(n_1062),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1220),
.B(n_1017),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1236),
.B(n_1115),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1270),
.A2(n_1032),
.B(n_1277),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1248),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1174),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1176),
.A2(n_1141),
.B(n_1062),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1189),
.B(n_1082),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1248),
.B(n_1055),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1252),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1206),
.B(n_1091),
.Y(n_1377)
);

AOI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1197),
.A2(n_1060),
.B(n_1049),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1252),
.B(n_1091),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1253),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1253),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1255),
.A2(n_1104),
.B(n_1010),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1262),
.A2(n_1141),
.B(n_1031),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1281),
.B(n_1017),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1236),
.B(n_1115),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1255),
.A2(n_1010),
.B(n_1016),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1153),
.A2(n_1026),
.B1(n_1043),
.B2(n_1027),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1262),
.A2(n_1066),
.B(n_943),
.Y(n_1388)
);

NOR2x1_ASAP7_75t_SL g1389 ( 
.A(n_1262),
.B(n_1126),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1203),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1236),
.A2(n_1016),
.B(n_1021),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1266),
.B(n_1027),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1243),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1198),
.A2(n_1026),
.B1(n_1043),
.B2(n_1100),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1243),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1269),
.A2(n_1040),
.B(n_1051),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1243),
.B(n_1267),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1237),
.B(n_1085),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1267),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1203),
.B(n_1085),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_R g1401 ( 
.A(n_1246),
.B(n_1085),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1267),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1249),
.A2(n_1128),
.B(n_1131),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1269),
.A2(n_1040),
.B(n_1051),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1158),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1224),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1269),
.A2(n_1094),
.B(n_1139),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1222),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1222),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1185),
.A2(n_1021),
.B(n_1078),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1221),
.B(n_1084),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1251),
.A2(n_1139),
.B(n_1131),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1250),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1239),
.A2(n_1115),
.B(n_1073),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1250),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1223),
.A2(n_1218),
.B1(n_1169),
.B2(n_1184),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1205),
.B(n_1036),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1226),
.A2(n_1085),
.B(n_1119),
.C(n_1100),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1169),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1205),
.B(n_1036),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1258),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1181),
.B(n_1121),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1258),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1274),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1274),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1195),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1208),
.A2(n_1139),
.B(n_1131),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1195),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1209),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1195),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1182),
.A2(n_1106),
.B(n_1130),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1229),
.B(n_1100),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1223),
.A2(n_1100),
.B1(n_1119),
.B2(n_1135),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1297),
.A2(n_1217),
.B(n_1194),
.C(n_1188),
.Y(n_1434)
);

OAI211xp5_ASAP7_75t_L g1435 ( 
.A1(n_1370),
.A2(n_1224),
.B(n_1254),
.C(n_1256),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1356),
.A2(n_1288),
.B1(n_1321),
.B2(n_1316),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1341),
.A2(n_1128),
.B(n_1130),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1334),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1356),
.A2(n_1223),
.B1(n_1184),
.B2(n_1175),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1397),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1416),
.A2(n_1175),
.B1(n_1156),
.B2(n_1170),
.C(n_1179),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1375),
.B(n_1227),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1305),
.A2(n_1194),
.B(n_1188),
.C(n_1179),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1305),
.A2(n_1256),
.B1(n_1260),
.B2(n_1268),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1397),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1416),
.A2(n_1215),
.B1(n_1212),
.B2(n_1200),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1364),
.A2(n_1260),
.B1(n_1268),
.B2(n_1215),
.Y(n_1447)
);

OAI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1316),
.A2(n_1254),
.B(n_1119),
.C(n_1135),
.Y(n_1448)
);

OAI211xp5_ASAP7_75t_L g1449 ( 
.A1(n_1321),
.A2(n_1119),
.B(n_1135),
.C(n_1227),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1357),
.B(n_1102),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1359),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1364),
.A2(n_1344),
.B1(n_1422),
.B2(n_1394),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1375),
.B(n_1156),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1359),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1359),
.A2(n_1170),
.B1(n_1183),
.B2(n_1201),
.Y(n_1455)
);

OAI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1431),
.A2(n_1200),
.B1(n_1199),
.B2(n_1212),
.C(n_1215),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1332),
.B(n_1102),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1359),
.A2(n_1183),
.B1(n_1201),
.B2(n_1260),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1411),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1313),
.B(n_1127),
.C(n_1121),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1294),
.Y(n_1461)
);

OAI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1322),
.A2(n_1200),
.B1(n_1199),
.B2(n_1212),
.C(n_1215),
.Y(n_1462)
);

OAI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1322),
.A2(n_1200),
.B1(n_1199),
.B2(n_1212),
.C(n_1159),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1372),
.A2(n_1268),
.B1(n_1273),
.B2(n_1199),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1372),
.A2(n_1102),
.B1(n_1127),
.B2(n_1106),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1346),
.B(n_1160),
.Y(n_1466)
);

AOI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1363),
.A2(n_1166),
.B(n_1160),
.C(n_1127),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1372),
.A2(n_1127),
.B1(n_1105),
.B2(n_1109),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1332),
.B(n_1160),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1299),
.A2(n_1126),
.B(n_1115),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1306),
.A2(n_1127),
.B1(n_1143),
.B2(n_1109),
.C(n_1105),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1372),
.A2(n_1127),
.B1(n_1143),
.B2(n_1023),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1387),
.A2(n_1035),
.B1(n_1023),
.B2(n_1273),
.Y(n_1473)
);

AOI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1432),
.A2(n_1166),
.B(n_1160),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1291),
.A2(n_1023),
.B1(n_1035),
.B2(n_984),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1368),
.B(n_1166),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1291),
.A2(n_1035),
.B1(n_1023),
.B2(n_995),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1315),
.A2(n_1035),
.B1(n_1166),
.B2(n_1026),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1418),
.A2(n_1159),
.B1(n_1052),
.B2(n_1026),
.C(n_1209),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1406),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1405),
.B(n_1209),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1315),
.A2(n_1059),
.B1(n_1047),
.B2(n_1052),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1314),
.A2(n_1083),
.B1(n_1283),
.B2(n_1209),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1378),
.A2(n_1103),
.B1(n_1083),
.B2(n_6),
.C(n_7),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1286),
.B(n_1083),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1418),
.A2(n_1335),
.B1(n_1299),
.B2(n_1412),
.C(n_1345),
.Y(n_1486)
);

AOI222xp33_ASAP7_75t_L g1487 ( 
.A1(n_1422),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_9),
.C2(n_12),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1397),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1335),
.A2(n_1059),
.B1(n_1076),
.B2(n_1083),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1426),
.B(n_1283),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1347),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1405),
.B(n_1059),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1392),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.C(n_15),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1333),
.A2(n_1076),
.B1(n_1059),
.B2(n_1047),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1391),
.A2(n_1078),
.B(n_1086),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1406),
.A2(n_1076),
.B1(n_1047),
.B2(n_1003),
.Y(n_1496)
);

AOI222xp33_ASAP7_75t_L g1497 ( 
.A1(n_1384),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_21),
.C2(n_22),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1342),
.B(n_1276),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1393),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1374),
.B(n_1073),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1329),
.B(n_1073),
.Y(n_1501)
);

OAI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1351),
.A2(n_1047),
.B1(n_1178),
.B2(n_994),
.C1(n_989),
.C2(n_1118),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1338),
.A2(n_1419),
.B1(n_1405),
.B2(n_1406),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1430),
.B(n_1126),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1317),
.A2(n_997),
.B(n_989),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1343),
.B(n_1073),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1373),
.A2(n_16),
.B(n_23),
.C(n_25),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1406),
.A2(n_1118),
.B1(n_1125),
.B2(n_1276),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1295),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1419),
.A2(n_1125),
.B1(n_27),
.B2(n_29),
.C(n_30),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1391),
.A2(n_1086),
.B(n_1092),
.Y(n_1512)
);

BUFx12f_ASAP7_75t_L g1513 ( 
.A(n_1338),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1377),
.B(n_1285),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1323),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1401),
.A2(n_1276),
.B1(n_27),
.B2(n_30),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1353),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1353),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1400),
.B(n_1092),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1383),
.A2(n_1087),
.B(n_1111),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1369),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1339),
.B(n_26),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1427),
.A2(n_1151),
.B1(n_32),
.B2(n_34),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1366),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1433),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_1525)
);

OAI21xp33_ASAP7_75t_L g1526 ( 
.A1(n_1304),
.A2(n_163),
.B(n_37),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1323),
.A2(n_1151),
.B1(n_38),
.B2(n_39),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1323),
.A2(n_1087),
.B1(n_1110),
.B2(n_1111),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1323),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1328),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1417),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1403),
.A2(n_1300),
.B1(n_1365),
.B2(n_1293),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1311),
.A2(n_1388),
.B(n_1404),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_R g1534 ( 
.A(n_1307),
.B(n_42),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1331),
.B(n_45),
.Y(n_1535)
);

OAI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1433),
.A2(n_45),
.B1(n_163),
.B2(n_159),
.C(n_157),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1319),
.A2(n_1110),
.B(n_1093),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1302),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1354),
.B(n_1093),
.Y(n_1539)
);

AOI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1310),
.A2(n_159),
.B1(n_163),
.B2(n_179),
.C(n_139),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1403),
.A2(n_1300),
.B1(n_1365),
.B2(n_1293),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1318),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1389),
.A2(n_157),
.A3(n_139),
.B(n_134),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1293),
.A2(n_159),
.B1(n_163),
.B2(n_133),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1337),
.B(n_159),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1420),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1398),
.Y(n_1547)
);

AOI33xp33_ASAP7_75t_L g1548 ( 
.A1(n_1324),
.A2(n_139),
.A3(n_157),
.B1(n_149),
.B2(n_226),
.B3(n_180),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1287),
.A2(n_159),
.B1(n_163),
.B2(n_133),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1393),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1325),
.A2(n_163),
.B1(n_157),
.B2(n_159),
.Y(n_1551)
);

NOR2x1_ASAP7_75t_R g1552 ( 
.A(n_1328),
.B(n_164),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1287),
.A2(n_159),
.B1(n_163),
.B2(n_133),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1307),
.A2(n_159),
.B1(n_163),
.B2(n_133),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1369),
.B(n_159),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1395),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_SL g1557 ( 
.A(n_1336),
.B(n_1367),
.C(n_1407),
.Y(n_1557)
);

OAI211xp5_ASAP7_75t_L g1558 ( 
.A1(n_1303),
.A2(n_163),
.B(n_159),
.C(n_139),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1429),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1366),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1307),
.A2(n_159),
.B1(n_163),
.B2(n_133),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1325),
.A2(n_159),
.B1(n_133),
.B2(n_156),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1390),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1395),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1301),
.B(n_159),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1400),
.B(n_159),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1327),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1303),
.A2(n_159),
.B1(n_135),
.B2(n_164),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1347),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1330),
.B(n_159),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1360),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1371),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1371),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1301),
.B(n_139),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1325),
.A2(n_133),
.B1(n_156),
.B2(n_149),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1340),
.A2(n_149),
.B(n_156),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1289),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1413),
.B(n_156),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1352),
.A2(n_156),
.B1(n_149),
.B2(n_150),
.C(n_134),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1340),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1325),
.A2(n_156),
.B1(n_135),
.B2(n_134),
.Y(n_1581)
);

OAI221xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1348),
.A2(n_156),
.B1(n_149),
.B2(n_221),
.C(n_180),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1303),
.A2(n_134),
.B1(n_149),
.B2(n_183),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1401),
.A2(n_149),
.B1(n_134),
.B2(n_183),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1289),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1348),
.A2(n_183),
.B1(n_207),
.B2(n_201),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1428),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1410),
.A2(n_134),
.B1(n_183),
.B2(n_198),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1290),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1348),
.A2(n_134),
.B1(n_198),
.B2(n_199),
.Y(n_1590)
);

AOI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1415),
.A2(n_198),
.B(n_207),
.C(n_201),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1421),
.B(n_198),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1513),
.B(n_1428),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1517),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1445),
.B(n_1348),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1517),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1571),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1445),
.B(n_1440),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1510),
.B(n_1326),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1573),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1518),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1451),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1438),
.B(n_1500),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1518),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1563),
.B(n_1326),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1488),
.B(n_1347),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1451),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1436),
.A2(n_1369),
.B1(n_1385),
.B2(n_1337),
.Y(n_1608)
);

NAND2x1_ASAP7_75t_L g1609 ( 
.A(n_1506),
.B(n_1337),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1524),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1524),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1560),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1521),
.B(n_1469),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1560),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1461),
.B(n_1379),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1451),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1572),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1509),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1453),
.B(n_1429),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1436),
.A2(n_1385),
.B1(n_1410),
.B2(n_1358),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1491),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_1385),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1538),
.B(n_1542),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1526),
.A2(n_1396),
.B(n_1358),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1567),
.B(n_1379),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1497),
.A2(n_1410),
.B1(n_1362),
.B2(n_1361),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1547),
.B(n_1290),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1534),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1534),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1585),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1467),
.B(n_1308),
.Y(n_1633)
);

BUFx8_ASAP7_75t_L g1634 ( 
.A(n_1451),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1491),
.B(n_1308),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1501),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1569),
.B(n_1361),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1589),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1569),
.B(n_1559),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1506),
.B(n_1361),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1499),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1506),
.B(n_1362),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1559),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1550),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1514),
.B(n_1292),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1556),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1559),
.B(n_1362),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1530),
.B(n_1425),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1564),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1460),
.B(n_1402),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1574),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1515),
.B(n_1424),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1442),
.B(n_1423),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1559),
.B(n_1408),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1539),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1489),
.A2(n_1380),
.A3(n_1376),
.B(n_1381),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1565),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1487),
.A2(n_1399),
.B(n_1409),
.C(n_1414),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1533),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1533),
.B(n_1296),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1533),
.Y(n_1661)
);

BUFx2_ASAP7_75t_SL g1662 ( 
.A(n_1454),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1587),
.B(n_1296),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1459),
.B(n_1292),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1447),
.B(n_1320),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1493),
.A2(n_1414),
.B1(n_1355),
.B2(n_1349),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1480),
.Y(n_1667)
);

AND2x4_ASAP7_75t_SL g1668 ( 
.A(n_1480),
.B(n_1515),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1485),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1532),
.B(n_1541),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1507),
.A2(n_1311),
.B(n_1350),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1535),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1476),
.Y(n_1673)
);

AO31x2_ASAP7_75t_L g1674 ( 
.A1(n_1505),
.A2(n_1381),
.A3(n_1380),
.B(n_1376),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1437),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1437),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1504),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1486),
.A2(n_1386),
.B(n_1355),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1543),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1466),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1452),
.B(n_1320),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1580),
.B(n_1312),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1570),
.Y(n_1683)
);

AO21x2_ASAP7_75t_L g1684 ( 
.A1(n_1557),
.A2(n_1350),
.B(n_1312),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1543),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1480),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1531),
.B(n_1386),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1546),
.B(n_1386),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1444),
.B(n_1382),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1522),
.B(n_1382),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1450),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1457),
.B(n_1355),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1543),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1532),
.B(n_1382),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1543),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1566),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1519),
.B(n_1349),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1494),
.B(n_1349),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1592),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1495),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1495),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1495),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1454),
.Y(n_1703)
);

AO31x2_ASAP7_75t_L g1704 ( 
.A1(n_1470),
.A2(n_180),
.A3(n_207),
.B(n_201),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1490),
.B(n_221),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1512),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1578),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1464),
.B(n_221),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1449),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1474),
.B(n_180),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1512),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1456),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1541),
.B(n_177),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1439),
.B(n_207),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1481),
.B(n_177),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1480),
.Y(n_1716)
);

AO31x2_ASAP7_75t_L g1717 ( 
.A1(n_1537),
.A2(n_177),
.A3(n_200),
.B(n_199),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1512),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1515),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1515),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1520),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1443),
.B(n_174),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1690),
.B(n_1462),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1619),
.Y(n_1724)
);

AO21x2_ASAP7_75t_L g1725 ( 
.A1(n_1670),
.A2(n_1507),
.B(n_1516),
.Y(n_1725)
);

OR2x2_ASAP7_75t_SL g1726 ( 
.A(n_1630),
.B(n_1458),
.Y(n_1726)
);

NOR3xp33_ASAP7_75t_L g1727 ( 
.A(n_1658),
.B(n_1435),
.C(n_1484),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1660),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1619),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1625),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1630),
.B(n_1443),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1609),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1631),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1628),
.A2(n_1631),
.B1(n_1712),
.B2(n_1709),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1672),
.B(n_1481),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1672),
.B(n_1455),
.Y(n_1736)
);

AO31x2_ASAP7_75t_L g1737 ( 
.A1(n_1678),
.A2(n_1446),
.A3(n_1434),
.B(n_1492),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1597),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1657),
.B(n_1439),
.Y(n_1739)
);

OAI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1628),
.A2(n_1463),
.B1(n_1479),
.B2(n_1441),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1625),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1634),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1660),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1597),
.Y(n_1744)
);

AOI222xp33_ASAP7_75t_L g1745 ( 
.A1(n_1658),
.A2(n_1529),
.B1(n_1525),
.B2(n_1511),
.C1(n_1434),
.C2(n_1536),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1634),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1678),
.A2(n_1458),
.B(n_1455),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1634),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1660),
.Y(n_1749)
);

AO31x2_ASAP7_75t_L g1750 ( 
.A1(n_1675),
.A2(n_1492),
.A3(n_1496),
.B(n_1586),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1622),
.A2(n_1671),
.B(n_1670),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1600),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1600),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1615),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1615),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1668),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1627),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1666),
.A2(n_1503),
.B1(n_1523),
.B2(n_1473),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1712),
.A2(n_1523),
.B1(n_1529),
.B2(n_1503),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1594),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1709),
.B(n_1483),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1627),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_SL g1763 ( 
.A(n_1593),
.B(n_1448),
.C(n_1584),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1670),
.A2(n_1527),
.B1(n_1473),
.B2(n_1482),
.Y(n_1764)
);

AOI21xp33_ASAP7_75t_L g1765 ( 
.A1(n_1666),
.A2(n_1552),
.B(n_1545),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1594),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1657),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1694),
.A2(n_1588),
.B(n_1583),
.Y(n_1768)
);

INVx5_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1651),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1594),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1707),
.B(n_1471),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1651),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1596),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1608),
.A2(n_1482),
.B1(n_1527),
.B2(n_1478),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1671),
.A2(n_1498),
.B(n_1544),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1596),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1683),
.Y(n_1778)
);

AOI21xp33_ASAP7_75t_SL g1779 ( 
.A1(n_1681),
.A2(n_1545),
.B(n_1508),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1596),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1667),
.B(n_1716),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1601),
.Y(n_1782)
);

OA21x2_ASAP7_75t_L g1783 ( 
.A1(n_1694),
.A2(n_1588),
.B(n_1583),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_SL g1784 ( 
.A(n_1609),
.B(n_1465),
.C(n_1478),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1703),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1683),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1633),
.B(n_1465),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1691),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1626),
.A2(n_1555),
.B(n_1472),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1690),
.B(n_1544),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1659),
.A2(n_1520),
.B(n_1475),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1601),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1601),
.Y(n_1793)
);

O2A1O1Ixp5_ASAP7_75t_L g1794 ( 
.A1(n_1689),
.A2(n_1502),
.B(n_1558),
.C(n_1555),
.Y(n_1794)
);

AO21x2_ASAP7_75t_L g1795 ( 
.A1(n_1675),
.A2(n_1590),
.B(n_1576),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1602),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1703),
.Y(n_1797)
);

AO31x2_ASAP7_75t_L g1798 ( 
.A1(n_1675),
.A2(n_1676),
.A3(n_1661),
.B(n_1659),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1696),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1696),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1633),
.B(n_1472),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1633),
.B(n_1468),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1668),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1691),
.A2(n_1553),
.B1(n_1549),
.B2(n_1568),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1699),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1595),
.B(n_1468),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1604),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1604),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1604),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1698),
.A2(n_1553),
.B(n_1549),
.C(n_1561),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1668),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1664),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1707),
.B(n_1554),
.Y(n_1813)
);

INVx6_ASAP7_75t_L g1814 ( 
.A(n_1634),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1703),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1611),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1681),
.A2(n_1673),
.B1(n_1722),
.B2(n_1665),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1602),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1664),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1614),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1614),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1626),
.A2(n_1477),
.B(n_1475),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1686),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1610),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1699),
.B(n_1554),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1662),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1602),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1686),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1662),
.A2(n_1477),
.B1(n_1561),
.B2(n_1562),
.Y(n_1829)
);

AO21x2_ASAP7_75t_L g1830 ( 
.A1(n_1676),
.A2(n_1551),
.B(n_1575),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1603),
.B(n_1520),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_1607),
.Y(n_1832)
);

OAI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1659),
.A2(n_1581),
.B(n_1562),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1610),
.Y(n_1834)
);

INVx4_ASAP7_75t_SL g1835 ( 
.A(n_1607),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1798),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1742),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1733),
.Y(n_1838)
);

AO21x2_ASAP7_75t_L g1839 ( 
.A1(n_1751),
.A2(n_1661),
.B(n_1676),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1826),
.B(n_1719),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1823),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1736),
.B(n_1719),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1725),
.B(n_1673),
.Y(n_1843)
);

OAI31xp33_ASAP7_75t_L g1844 ( 
.A1(n_1731),
.A2(n_1722),
.A3(n_1689),
.B(n_1698),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1756),
.B(n_1719),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1798),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1724),
.Y(n_1847)
);

AOI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1734),
.A2(n_1727),
.B1(n_1758),
.B2(n_1740),
.C(n_1725),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1823),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1756),
.B(n_1720),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1724),
.Y(n_1851)
);

OAI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1747),
.A2(n_1636),
.B1(n_1720),
.B2(n_1655),
.C(n_1669),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1803),
.B(n_1720),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1828),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1828),
.Y(n_1855)
);

AO21x2_ASAP7_75t_L g1856 ( 
.A1(n_1725),
.A2(n_1661),
.B(n_1713),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1789),
.A2(n_1689),
.B1(n_1698),
.B2(n_1636),
.C(n_1626),
.Y(n_1857)
);

OAI33xp33_ASAP7_75t_L g1858 ( 
.A1(n_1770),
.A2(n_1773),
.A3(n_1761),
.B1(n_1741),
.B2(n_1730),
.B3(n_1790),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1803),
.B(n_1720),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1790),
.B(n_1603),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1745),
.A2(n_1626),
.B1(n_1722),
.B2(n_1698),
.Y(n_1861)
);

O2A1O1Ixp33_ASAP7_75t_SL g1862 ( 
.A1(n_1811),
.A2(n_1667),
.B(n_1716),
.C(n_1652),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1779),
.B(n_1669),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1729),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1811),
.B(n_1687),
.Y(n_1865)
);

INVx4_ASAP7_75t_L g1866 ( 
.A(n_1814),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1787),
.B(n_1687),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1759),
.A2(n_1655),
.B1(n_1716),
.B2(n_1667),
.C(n_1607),
.Y(n_1868)
);

OAI31xp33_ASAP7_75t_SL g1869 ( 
.A1(n_1784),
.A2(n_1689),
.A3(n_1688),
.B(n_1665),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1739),
.B(n_1708),
.C(n_1713),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1812),
.B(n_1677),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1769),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1812),
.B(n_1677),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1729),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1787),
.B(n_1688),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1801),
.B(n_1639),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1738),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1801),
.B(n_1639),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1732),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_L g1880 ( 
.A(n_1764),
.B(n_1794),
.C(n_1822),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1776),
.A2(n_1722),
.B1(n_1642),
.B2(n_1640),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1798),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1835),
.B(n_1640),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1781),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1819),
.B(n_1629),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1738),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1785),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1775),
.A2(n_1642),
.B(n_1640),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1802),
.B(n_1806),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1785),
.Y(n_1890)
);

AOI31xp33_ASAP7_75t_SL g1891 ( 
.A1(n_1765),
.A2(n_1629),
.A3(n_1693),
.B(n_1695),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1802),
.B(n_1639),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1744),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1806),
.B(n_1595),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1797),
.B(n_1815),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1797),
.B(n_1616),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1732),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1744),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1742),
.B(n_1616),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1781),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1752),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1798),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1815),
.B(n_1796),
.Y(n_1903)
);

NAND3xp33_ASAP7_75t_SL g1904 ( 
.A(n_1817),
.B(n_1708),
.C(n_1705),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1752),
.Y(n_1905)
);

INVx4_ASAP7_75t_L g1906 ( 
.A(n_1814),
.Y(n_1906)
);

OAI31xp33_ASAP7_75t_L g1907 ( 
.A1(n_1726),
.A2(n_1616),
.A3(n_1650),
.B(n_1714),
.Y(n_1907)
);

NAND3xp33_ASAP7_75t_L g1908 ( 
.A(n_1768),
.B(n_1710),
.C(n_1715),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1732),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1746),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1723),
.A2(n_1680),
.B1(n_1684),
.B2(n_1645),
.C(n_1692),
.Y(n_1911)
);

INVxp67_ASAP7_75t_L g1912 ( 
.A(n_1735),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1796),
.B(n_1640),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1796),
.B(n_1642),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1798),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1753),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1819),
.B(n_1645),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1818),
.B(n_1642),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1788),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1753),
.Y(n_1920)
);

BUFx2_ASAP7_75t_L g1921 ( 
.A(n_1781),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1778),
.B(n_1605),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1814),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1818),
.B(n_1598),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1728),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1835),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1818),
.B(n_1598),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1726),
.B(n_1680),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1827),
.B(n_1624),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1827),
.B(n_1624),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1835),
.B(n_1684),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1855),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1889),
.B(n_1835),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1926),
.B(n_1769),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1855),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1838),
.B(n_1723),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1884),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1838),
.B(n_1786),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1841),
.Y(n_1939)
);

OA21x2_ASAP7_75t_L g1940 ( 
.A1(n_1848),
.A2(n_1791),
.B(n_1711),
.Y(n_1940)
);

NAND2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1926),
.B(n_1746),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1889),
.B(n_1827),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1849),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1854),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1919),
.B(n_1767),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1867),
.B(n_1832),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1867),
.B(n_1832),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1860),
.B(n_1754),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1875),
.B(n_1748),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1875),
.B(n_1748),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1924),
.B(n_1769),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1861),
.B(n_1769),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1847),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1884),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1837),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1860),
.B(n_1754),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1924),
.B(n_1769),
.Y(n_1957)
);

OAI33xp33_ASAP7_75t_L g1958 ( 
.A1(n_1880),
.A2(n_1821),
.A3(n_1820),
.B1(n_1762),
.B2(n_1757),
.B3(n_1755),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1927),
.B(n_1755),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1927),
.B(n_1757),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1922),
.B(n_1762),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1894),
.B(n_1737),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1883),
.B(n_1820),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1894),
.B(n_1737),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1922),
.B(n_1805),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1892),
.B(n_1737),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1900),
.Y(n_1967)
);

INVx4_ASAP7_75t_L g1968 ( 
.A(n_1866),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1900),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1847),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1892),
.B(n_1895),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1921),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1912),
.B(n_1799),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1921),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1895),
.B(n_1737),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1836),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1851),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1836),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1836),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1928),
.B(n_1800),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1858),
.B(n_1814),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1856),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1880),
.A2(n_1768),
.B1(n_1783),
.B2(n_1772),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1843),
.B(n_1821),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1851),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1910),
.B(n_1887),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1846),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1861),
.A2(n_1763),
.B1(n_1810),
.B2(n_1783),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1876),
.B(n_1737),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1864),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1876),
.B(n_1643),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1879),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1864),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1878),
.B(n_1643),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1846),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1874),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1846),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1878),
.B(n_1643),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1887),
.B(n_1834),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1903),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1874),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1877),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1885),
.B(n_1824),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1882),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1885),
.B(n_1824),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1883),
.B(n_1834),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1903),
.B(n_1643),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1890),
.B(n_1813),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1845),
.B(n_1728),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1842),
.A2(n_1795),
.B1(n_1783),
.B2(n_1768),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1845),
.B(n_1743),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1850),
.B(n_1743),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_R g2013 ( 
.A(n_1923),
.B(n_1705),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1837),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1877),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1886),
.Y(n_2016)
);

INVx4_ASAP7_75t_L g2017 ( 
.A(n_1866),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1882),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1986),
.B(n_1863),
.Y(n_2019)
);

XNOR2xp5_ASAP7_75t_L g2020 ( 
.A(n_1988),
.B(n_1899),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1986),
.B(n_1837),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1955),
.Y(n_2022)
);

AND4x1_ASAP7_75t_L g2023 ( 
.A(n_1981),
.B(n_1907),
.C(n_1869),
.D(n_1933),
.Y(n_2023)
);

OAI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1988),
.A2(n_1907),
.B(n_1868),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1955),
.B(n_1923),
.Y(n_2025)
);

AND2x4_ASAP7_75t_SL g2026 ( 
.A(n_1971),
.B(n_1866),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_1982),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1954),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1949),
.B(n_1923),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1954),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1955),
.B(n_2014),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1949),
.B(n_1923),
.Y(n_2032)
);

NAND4xp75_ASAP7_75t_SL g2033 ( 
.A(n_1981),
.B(n_1844),
.C(n_1840),
.D(n_1859),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1932),
.B(n_1870),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1972),
.Y(n_2035)
);

NAND4xp75_ASAP7_75t_L g2036 ( 
.A(n_1952),
.B(n_2010),
.C(n_1933),
.D(n_1857),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1972),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1939),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1939),
.Y(n_2039)
);

XNOR2xp5_ASAP7_75t_L g2040 ( 
.A(n_1971),
.B(n_1888),
.Y(n_2040)
);

AND4x1_ASAP7_75t_L g2041 ( 
.A(n_2010),
.B(n_1844),
.C(n_1896),
.D(n_1881),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1932),
.B(n_1840),
.Y(n_2042)
);

XNOR2xp5_ASAP7_75t_L g2043 ( 
.A(n_1950),
.B(n_1904),
.Y(n_2043)
);

NAND4xp75_ASAP7_75t_SL g2044 ( 
.A(n_1950),
.B(n_1850),
.C(n_1859),
.D(n_1853),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1942),
.B(n_1866),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1942),
.B(n_1946),
.Y(n_2046)
);

XNOR2x2_ASAP7_75t_L g2047 ( 
.A(n_1935),
.B(n_2000),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2014),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_2008),
.B(n_1908),
.Y(n_2049)
);

XOR2xp5_ASAP7_75t_L g2050 ( 
.A(n_1983),
.B(n_1804),
.Y(n_2050)
);

INVx4_ASAP7_75t_L g2051 ( 
.A(n_1968),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1983),
.A2(n_1906),
.B1(n_1852),
.B2(n_1883),
.Y(n_2052)
);

NOR4xp25_ASAP7_75t_L g2053 ( 
.A(n_1935),
.B(n_1891),
.C(n_1911),
.D(n_1908),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1941),
.Y(n_2054)
);

NOR3xp33_ASAP7_75t_SL g2055 ( 
.A(n_2008),
.B(n_1906),
.C(n_1898),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1941),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1934),
.Y(n_2057)
);

XNOR2x1_ASAP7_75t_L g2058 ( 
.A(n_1941),
.B(n_1896),
.Y(n_2058)
);

NOR2x1_ASAP7_75t_R g2059 ( 
.A(n_1968),
.B(n_1906),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_1946),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1937),
.B(n_1856),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1937),
.B(n_1856),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1992),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1958),
.A2(n_1906),
.B1(n_1883),
.B2(n_1865),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_2000),
.B(n_1862),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1937),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_1934),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1947),
.B(n_1865),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1967),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1967),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1936),
.A2(n_1829),
.B1(n_1872),
.B2(n_1891),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1992),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_R g2073 ( 
.A(n_1943),
.B(n_1872),
.Y(n_2073)
);

XNOR2xp5_ASAP7_75t_L g2074 ( 
.A(n_1947),
.B(n_1853),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_1934),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1967),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1992),
.Y(n_2077)
);

NAND4xp75_ASAP7_75t_L g2078 ( 
.A(n_1975),
.B(n_1913),
.C(n_1914),
.D(n_1918),
.Y(n_2078)
);

INVx5_ASAP7_75t_L g2079 ( 
.A(n_1968),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1958),
.A2(n_1930),
.B1(n_1929),
.B2(n_1795),
.Y(n_2080)
);

NAND3xp33_ASAP7_75t_L g2081 ( 
.A(n_1936),
.B(n_1886),
.C(n_1901),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1969),
.Y(n_2082)
);

NAND4xp75_ASAP7_75t_L g2083 ( 
.A(n_1975),
.B(n_1914),
.C(n_1913),
.D(n_1918),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1969),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2007),
.B(n_1929),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1969),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1934),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1974),
.Y(n_2088)
);

NOR2x1_ASAP7_75t_R g2089 ( 
.A(n_1968),
.B(n_1825),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_1974),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2007),
.B(n_1991),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1974),
.B(n_1893),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_2017),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1943),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_1982),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1944),
.B(n_1945),
.Y(n_2096)
);

XOR2xp5_ASAP7_75t_L g2097 ( 
.A(n_1980),
.B(n_1930),
.Y(n_2097)
);

INVx2_ASAP7_75t_SL g2098 ( 
.A(n_1951),
.Y(n_2098)
);

NOR2xp67_ASAP7_75t_L g2099 ( 
.A(n_2022),
.B(n_2017),
.Y(n_2099)
);

OR2x6_ASAP7_75t_L g2100 ( 
.A(n_2031),
.B(n_2017),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2046),
.B(n_1991),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2048),
.B(n_1944),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2019),
.B(n_1980),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2090),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2021),
.B(n_1973),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_2053),
.B(n_2017),
.Y(n_2106)
);

INVx2_ASAP7_75t_SL g2107 ( 
.A(n_2031),
.Y(n_2107)
);

AOI32xp33_ASAP7_75t_SL g2108 ( 
.A1(n_2065),
.A2(n_1973),
.A3(n_1945),
.B1(n_1999),
.B2(n_2016),
.Y(n_2108)
);

OR2x6_ASAP7_75t_L g2109 ( 
.A(n_2051),
.B(n_1951),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2028),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2030),
.B(n_1959),
.Y(n_2111)
);

INVxp67_ASAP7_75t_SL g2112 ( 
.A(n_2047),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2042),
.B(n_1948),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2042),
.B(n_2049),
.Y(n_2114)
);

INVxp67_ASAP7_75t_SL g2115 ( 
.A(n_2089),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2035),
.Y(n_2116)
);

INVx2_ASAP7_75t_SL g2117 ( 
.A(n_2056),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2057),
.Y(n_2118)
);

OAI31xp33_ASAP7_75t_L g2119 ( 
.A1(n_2071),
.A2(n_1966),
.A3(n_1989),
.B(n_1962),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2037),
.B(n_1959),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2034),
.B(n_1948),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2095),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2029),
.B(n_2032),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2095),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2025),
.B(n_1963),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2068),
.B(n_2045),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2038),
.B(n_1960),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_2027),
.Y(n_2128)
);

OR2x6_ASAP7_75t_L g2129 ( 
.A(n_2051),
.B(n_1957),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2057),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2066),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2087),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2069),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2034),
.B(n_1956),
.Y(n_2134)
);

INVxp67_ASAP7_75t_SL g2135 ( 
.A(n_2020),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2060),
.B(n_1956),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2098),
.B(n_1999),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2070),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2076),
.Y(n_2139)
);

A2O1A1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_2024),
.A2(n_1989),
.B(n_1966),
.C(n_1962),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2096),
.B(n_1938),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2082),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2087),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2085),
.B(n_1994),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2084),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2086),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2027),
.Y(n_2147)
);

AO22x1_ASAP7_75t_L g2148 ( 
.A1(n_2024),
.A2(n_1957),
.B1(n_1963),
.B2(n_2006),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2025),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2091),
.B(n_1994),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_2063),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2039),
.B(n_1960),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2053),
.B(n_1938),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_2026),
.Y(n_2154)
);

INVx1_ASAP7_75t_SL g2155 ( 
.A(n_2058),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2096),
.B(n_2071),
.Y(n_2156)
);

NAND3xp33_ASAP7_75t_L g2157 ( 
.A(n_2041),
.B(n_1940),
.C(n_1963),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2088),
.Y(n_2158)
);

A2O1A1Ixp33_ASAP7_75t_L g2159 ( 
.A1(n_2055),
.A2(n_1964),
.B(n_1984),
.C(n_1833),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_2054),
.Y(n_2160)
);

OAI221xp5_ASAP7_75t_L g2161 ( 
.A1(n_2112),
.A2(n_2050),
.B1(n_2023),
.B2(n_2052),
.C(n_2055),
.Y(n_2161)
);

NAND2x1_ASAP7_75t_SL g2162 ( 
.A(n_2125),
.B(n_2064),
.Y(n_2162)
);

AO21x1_ASAP7_75t_L g2163 ( 
.A1(n_2112),
.A2(n_2062),
.B(n_2061),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2136),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2125),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2153),
.A2(n_2043),
.B(n_2061),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2107),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2155),
.B(n_2067),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2100),
.Y(n_2169)
);

OAI211xp5_ASAP7_75t_L g2170 ( 
.A1(n_2106),
.A2(n_2073),
.B(n_2080),
.C(n_2094),
.Y(n_2170)
);

AOI21xp5_ASAP7_75t_SL g2171 ( 
.A1(n_2106),
.A2(n_2059),
.B(n_2062),
.Y(n_2171)
);

INVxp67_ASAP7_75t_L g2172 ( 
.A(n_2128),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2128),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2147),
.Y(n_2174)
);

AOI211x1_ASAP7_75t_L g2175 ( 
.A1(n_2157),
.A2(n_2081),
.B(n_2092),
.C(n_2033),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2135),
.A2(n_2036),
.B1(n_2040),
.B2(n_2074),
.Y(n_2176)
);

O2A1O1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_2153),
.A2(n_2067),
.B(n_2075),
.C(n_2033),
.Y(n_2177)
);

OAI221xp5_ASAP7_75t_SL g2178 ( 
.A1(n_2119),
.A2(n_2097),
.B1(n_2075),
.B2(n_1964),
.C(n_1984),
.Y(n_2178)
);

INVxp67_ASAP7_75t_L g2179 ( 
.A(n_2147),
.Y(n_2179)
);

INVxp67_ASAP7_75t_SL g2180 ( 
.A(n_2099),
.Y(n_2180)
);

OAI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_2156),
.A2(n_1940),
.B1(n_1879),
.B2(n_1909),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2151),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2135),
.A2(n_1940),
.B1(n_1879),
.B2(n_1909),
.Y(n_2183)
);

OAI21xp33_ASAP7_75t_L g2184 ( 
.A1(n_2123),
.A2(n_1963),
.B(n_1998),
.Y(n_2184)
);

OAI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2140),
.A2(n_2083),
.B1(n_2078),
.B2(n_1940),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2151),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2104),
.Y(n_2187)
);

OAI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_2159),
.A2(n_2140),
.B(n_2115),
.Y(n_2188)
);

AOI21xp33_ASAP7_75t_L g2189 ( 
.A1(n_2115),
.A2(n_1940),
.B(n_2093),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_2148),
.A2(n_2092),
.B(n_2077),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2114),
.B(n_1965),
.Y(n_2191)
);

OAI21xp33_ASAP7_75t_L g2192 ( 
.A1(n_2154),
.A2(n_1998),
.B(n_2013),
.Y(n_2192)
);

OAI211xp5_ASAP7_75t_SL g2193 ( 
.A1(n_2103),
.A2(n_2093),
.B(n_2072),
.C(n_1970),
.Y(n_2193)
);

AOI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2101),
.A2(n_2009),
.B1(n_2011),
.B2(n_2012),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2122),
.Y(n_2195)
);

XNOR2xp5_ASAP7_75t_L g2196 ( 
.A(n_2126),
.B(n_2044),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2124),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2100),
.Y(n_2198)
);

NAND3xp33_ASAP7_75t_SL g2199 ( 
.A(n_2159),
.B(n_2044),
.C(n_1970),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2100),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2150),
.B(n_2079),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2144),
.B(n_2079),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2109),
.Y(n_2203)
);

A2O1A1Ixp33_ASAP7_75t_L g2204 ( 
.A1(n_2121),
.A2(n_1931),
.B(n_2079),
.C(n_2016),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2149),
.B(n_2079),
.Y(n_2205)
);

XNOR2xp5_ASAP7_75t_L g2206 ( 
.A(n_2117),
.B(n_2006),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2109),
.Y(n_2207)
);

OAI31xp33_ASAP7_75t_L g2208 ( 
.A1(n_2134),
.A2(n_1931),
.A3(n_2006),
.B(n_1897),
.Y(n_2208)
);

OA22x2_ASAP7_75t_L g2209 ( 
.A1(n_2118),
.A2(n_2006),
.B1(n_2015),
.B2(n_1985),
.Y(n_2209)
);

CKINVDCx16_ASAP7_75t_R g2210 ( 
.A(n_2109),
.Y(n_2210)
);

NOR2x1_ASAP7_75t_L g2211 ( 
.A(n_2129),
.B(n_1953),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2102),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2209),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2211),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2210),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2167),
.B(n_2130),
.Y(n_2216)
);

HB1xp67_ASAP7_75t_L g2217 ( 
.A(n_2172),
.Y(n_2217)
);

A2O1A1Ixp33_ASAP7_75t_L g2218 ( 
.A1(n_2177),
.A2(n_2141),
.B(n_2113),
.C(n_2120),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2166),
.B(n_2132),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2209),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2172),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2165),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2161),
.A2(n_2160),
.B1(n_2143),
.B2(n_2120),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2164),
.B(n_2129),
.Y(n_2224)
);

OR2x2_ASAP7_75t_L g2225 ( 
.A(n_2168),
.B(n_2111),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2173),
.Y(n_2226)
);

AOI322xp5_ASAP7_75t_L g2227 ( 
.A1(n_2199),
.A2(n_2108),
.A3(n_2110),
.B1(n_2116),
.B2(n_2102),
.C1(n_2152),
.C2(n_2127),
.Y(n_2227)
);

AOI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2177),
.A2(n_2127),
.B1(n_2152),
.B2(n_2111),
.C(n_2145),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2174),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2173),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2191),
.B(n_2137),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2166),
.B(n_2105),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2180),
.Y(n_2233)
);

OAI22xp33_ASAP7_75t_SL g2234 ( 
.A1(n_2178),
.A2(n_2129),
.B1(n_2146),
.B2(n_2142),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2187),
.B(n_2131),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2178),
.A2(n_2158),
.B1(n_2139),
.B2(n_2138),
.C(n_2133),
.Y(n_2236)
);

AOI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2175),
.A2(n_1990),
.B1(n_2015),
.B2(n_1993),
.C(n_1985),
.Y(n_2237)
);

AOI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_2176),
.A2(n_1990),
.B(n_2002),
.Y(n_2238)
);

A2O1A1Ixp33_ASAP7_75t_L g2239 ( 
.A1(n_2162),
.A2(n_2188),
.B(n_2170),
.C(n_2199),
.Y(n_2239)
);

OAI221xp5_ASAP7_75t_L g2240 ( 
.A1(n_2170),
.A2(n_1965),
.B1(n_1961),
.B2(n_1953),
.C(n_1993),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2179),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2179),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2202),
.B(n_2009),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2182),
.Y(n_2244)
);

AOI21xp33_ASAP7_75t_SL g2245 ( 
.A1(n_2185),
.A2(n_1977),
.B(n_1996),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2186),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2201),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_L g2248 ( 
.A(n_2203),
.B(n_1879),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2195),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_SL g2250 ( 
.A1(n_2189),
.A2(n_2005),
.B(n_2003),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2207),
.B(n_2011),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2197),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2190),
.A2(n_1996),
.B1(n_1977),
.B2(n_2001),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2205),
.B(n_2012),
.Y(n_2254)
);

INVxp67_ASAP7_75t_L g2255 ( 
.A(n_2190),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2192),
.A2(n_1961),
.B1(n_2002),
.B2(n_2001),
.C(n_1897),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2193),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2193),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2184),
.B(n_2003),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2163),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2206),
.B(n_1897),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2183),
.A2(n_1839),
.B1(n_1931),
.B2(n_1795),
.Y(n_2262)
);

NOR2x1_ASAP7_75t_L g2263 ( 
.A(n_2171),
.B(n_1897),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2169),
.B(n_2005),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2217),
.Y(n_2265)
);

OAI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2239),
.A2(n_2255),
.B(n_2214),
.Y(n_2266)
);

OAI21xp33_ASAP7_75t_L g2267 ( 
.A1(n_2239),
.A2(n_2215),
.B(n_2196),
.Y(n_2267)
);

OAI31xp33_ASAP7_75t_L g2268 ( 
.A1(n_2234),
.A2(n_2181),
.A3(n_2204),
.B(n_2212),
.Y(n_2268)
);

INVx1_ASAP7_75t_SL g2269 ( 
.A(n_2231),
.Y(n_2269)
);

AOI32xp33_ASAP7_75t_L g2270 ( 
.A1(n_2260),
.A2(n_2200),
.A3(n_2198),
.B1(n_1931),
.B2(n_1909),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2243),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2233),
.B(n_2194),
.Y(n_2272)
);

AOI21xp33_ASAP7_75t_SL g2273 ( 
.A1(n_2253),
.A2(n_2208),
.B(n_1839),
.Y(n_2273)
);

AOI211xp5_ASAP7_75t_L g2274 ( 
.A1(n_2253),
.A2(n_1905),
.B(n_1893),
.C(n_1898),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_2263),
.Y(n_2275)
);

OAI221xp5_ASAP7_75t_L g2276 ( 
.A1(n_2255),
.A2(n_1909),
.B1(n_1905),
.B2(n_1916),
.C(n_1920),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2217),
.Y(n_2277)
);

INVxp67_ASAP7_75t_L g2278 ( 
.A(n_2224),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2214),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2233),
.B(n_1901),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2232),
.A2(n_1839),
.B(n_2004),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2216),
.B(n_1916),
.Y(n_2282)
);

OAI21xp33_ASAP7_75t_L g2283 ( 
.A1(n_2223),
.A2(n_1925),
.B(n_1920),
.Y(n_2283)
);

OAI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2218),
.A2(n_2018),
.B1(n_2004),
.B2(n_1997),
.C(n_1995),
.Y(n_2284)
);

OAI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2219),
.A2(n_1925),
.B1(n_1917),
.B2(n_1873),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2251),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2261),
.B(n_1925),
.Y(n_2287)
);

NAND3x2_ASAP7_75t_L g2288 ( 
.A(n_2225),
.B(n_1917),
.C(n_1873),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2254),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2247),
.B(n_1871),
.Y(n_2290)
);

NOR3xp33_ASAP7_75t_L g2291 ( 
.A(n_2236),
.B(n_2228),
.C(n_2245),
.Y(n_2291)
);

XOR2x2_ASAP7_75t_L g2292 ( 
.A(n_2259),
.B(n_2264),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2222),
.B(n_1613),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2221),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2213),
.B(n_1871),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2226),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2257),
.B(n_1760),
.Y(n_2297)
);

A2O1A1Ixp33_ASAP7_75t_SL g2298 ( 
.A1(n_2230),
.A2(n_2241),
.B(n_2242),
.C(n_2258),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_SL g2299 ( 
.A(n_2220),
.B(n_1976),
.Y(n_2299)
);

OAI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2240),
.A2(n_2018),
.B1(n_2004),
.B2(n_1997),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2229),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2227),
.B(n_1749),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2244),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2269),
.B(n_2248),
.Y(n_2304)
);

AOI21xp33_ASAP7_75t_L g2305 ( 
.A1(n_2267),
.A2(n_2250),
.B(n_2248),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2278),
.B(n_2246),
.Y(n_2306)
);

OAI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2281),
.A2(n_2238),
.B(n_2237),
.Y(n_2307)
);

AOI221x1_ASAP7_75t_L g2308 ( 
.A1(n_2291),
.A2(n_2249),
.B1(n_2252),
.B2(n_2238),
.C(n_1976),
.Y(n_2308)
);

AOI211xp5_ASAP7_75t_SL g2309 ( 
.A1(n_2275),
.A2(n_2235),
.B(n_2256),
.C(n_2262),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_2278),
.B(n_2262),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2293),
.Y(n_2311)
);

NAND2xp33_ASAP7_75t_L g2312 ( 
.A(n_2270),
.B(n_1976),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2271),
.B(n_1749),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2265),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2289),
.B(n_2290),
.Y(n_2315)
);

OAI21xp33_ASAP7_75t_L g2316 ( 
.A1(n_2292),
.A2(n_2018),
.B(n_1997),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2302),
.A2(n_1995),
.B1(n_1987),
.B2(n_1979),
.Y(n_2317)
);

AOI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_2286),
.A2(n_1995),
.B1(n_1987),
.B2(n_1979),
.Y(n_2318)
);

XNOR2x1_ASAP7_75t_L g2319 ( 
.A(n_2266),
.B(n_1833),
.Y(n_2319)
);

NOR3x1_ASAP7_75t_L g2320 ( 
.A(n_2298),
.B(n_1791),
.C(n_1831),
.Y(n_2320)
);

NAND3xp33_ASAP7_75t_SL g2321 ( 
.A(n_2268),
.B(n_1987),
.C(n_1979),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2277),
.B(n_1760),
.Y(n_2322)
);

NOR2xp67_ASAP7_75t_L g2323 ( 
.A(n_2279),
.B(n_1978),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2281),
.A2(n_2299),
.B(n_2273),
.Y(n_2324)
);

BUFx2_ASAP7_75t_L g2325 ( 
.A(n_2288),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_2295),
.Y(n_2326)
);

AOI21xp33_ASAP7_75t_SL g2327 ( 
.A1(n_2285),
.A2(n_1978),
.B(n_1915),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2287),
.Y(n_2328)
);

AOI21xp33_ASAP7_75t_L g2329 ( 
.A1(n_2272),
.A2(n_1978),
.B(n_1915),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2294),
.B(n_1613),
.Y(n_2330)
);

NAND3x1_ASAP7_75t_L g2331 ( 
.A(n_2301),
.B(n_2296),
.C(n_2303),
.Y(n_2331)
);

OAI322xp33_ASAP7_75t_L g2332 ( 
.A1(n_2300),
.A2(n_2284),
.A3(n_2297),
.B1(n_2282),
.B2(n_2280),
.C1(n_2276),
.C2(n_2283),
.Y(n_2332)
);

OAI322xp33_ASAP7_75t_L g2333 ( 
.A1(n_2310),
.A2(n_2284),
.A3(n_2276),
.B1(n_1915),
.B2(n_1902),
.C1(n_1882),
.C2(n_2274),
.Y(n_2333)
);

OAI221xp5_ASAP7_75t_SL g2334 ( 
.A1(n_2316),
.A2(n_1902),
.B1(n_1831),
.B2(n_1816),
.C(n_1809),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2326),
.B(n_1766),
.Y(n_2335)
);

O2A1O1Ixp33_ASAP7_75t_L g2336 ( 
.A1(n_2307),
.A2(n_2321),
.B(n_2309),
.C(n_2324),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2330),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2304),
.Y(n_2338)
);

OAI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2307),
.A2(n_1902),
.B(n_1715),
.Y(n_2339)
);

OAI211xp5_ASAP7_75t_L g2340 ( 
.A1(n_2305),
.A2(n_1780),
.B(n_1816),
.C(n_1809),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2306),
.Y(n_2341)
);

OAI21xp5_ASAP7_75t_SL g2342 ( 
.A1(n_2309),
.A2(n_1714),
.B(n_1710),
.Y(n_2342)
);

AOI211xp5_ASAP7_75t_L g2343 ( 
.A1(n_2332),
.A2(n_1714),
.B(n_1808),
.C(n_1807),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2328),
.B(n_1766),
.Y(n_2344)
);

AOI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_2312),
.A2(n_1777),
.B(n_1808),
.Y(n_2345)
);

NAND4xp75_ASAP7_75t_L g2346 ( 
.A(n_2308),
.B(n_1780),
.C(n_1807),
.D(n_1793),
.Y(n_2346)
);

AOI211xp5_ASAP7_75t_L g2347 ( 
.A1(n_2315),
.A2(n_1774),
.B(n_1793),
.C(n_1792),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2319),
.A2(n_1771),
.B(n_1792),
.Y(n_2348)
);

OA211x2_ASAP7_75t_L g2349 ( 
.A1(n_2313),
.A2(n_1579),
.B(n_1581),
.C(n_1540),
.Y(n_2349)
);

OAI322xp33_ASAP7_75t_L g2350 ( 
.A1(n_2314),
.A2(n_1771),
.A3(n_1782),
.B1(n_1777),
.B2(n_1774),
.C1(n_1721),
.C2(n_1711),
.Y(n_2350)
);

NOR4xp25_ASAP7_75t_L g2351 ( 
.A(n_2331),
.B(n_1782),
.C(n_1721),
.D(n_1700),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2311),
.B(n_1684),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2325),
.B(n_1623),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_2323),
.A2(n_1830),
.B1(n_1684),
.B2(n_1721),
.Y(n_2354)
);

NAND4xp25_ASAP7_75t_SL g2355 ( 
.A(n_2327),
.B(n_1654),
.C(n_1692),
.D(n_1606),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2322),
.B(n_1623),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2335),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2337),
.Y(n_2358)
);

AOI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2353),
.A2(n_2338),
.B1(n_2341),
.B2(n_2355),
.Y(n_2359)
);

AO22x2_ASAP7_75t_L g2360 ( 
.A1(n_2336),
.A2(n_2317),
.B1(n_2320),
.B2(n_2329),
.Y(n_2360)
);

AOI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_2342),
.A2(n_2318),
.B1(n_1830),
.B2(n_1650),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_2356),
.A2(n_1623),
.B(n_1650),
.C(n_1700),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2346),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2344),
.Y(n_2364)
);

AOI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_2349),
.A2(n_1830),
.B1(n_1650),
.B2(n_1654),
.Y(n_2365)
);

AO22x1_ASAP7_75t_L g2366 ( 
.A1(n_2339),
.A2(n_1623),
.B1(n_1648),
.B2(n_1606),
.Y(n_2366)
);

A2O1A1Ixp33_ASAP7_75t_SL g2367 ( 
.A1(n_2334),
.A2(n_1702),
.B(n_1700),
.C(n_1701),
.Y(n_2367)
);

OAI22x1_ASAP7_75t_L g2368 ( 
.A1(n_2352),
.A2(n_1648),
.B1(n_1682),
.B2(n_1611),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2333),
.Y(n_2369)
);

AOI221xp5_ASAP7_75t_L g2370 ( 
.A1(n_2351),
.A2(n_1701),
.B1(n_1702),
.B2(n_1711),
.C(n_1706),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2343),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2340),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2348),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2347),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2345),
.Y(n_2375)
);

OAI31xp33_ASAP7_75t_L g2376 ( 
.A1(n_2345),
.A2(n_1682),
.A3(n_1697),
.B(n_1706),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2354),
.A2(n_1611),
.B1(n_1612),
.B2(n_1632),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2350),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2335),
.Y(n_2379)
);

AOI221xp5_ASAP7_75t_L g2380 ( 
.A1(n_2360),
.A2(n_1702),
.B1(n_1701),
.B2(n_1706),
.C(n_1718),
.Y(n_2380)
);

NOR3xp33_ASAP7_75t_L g2381 ( 
.A(n_2358),
.B(n_1718),
.C(n_1697),
.Y(n_2381)
);

AND4x1_ASAP7_75t_L g2382 ( 
.A(n_2359),
.B(n_1548),
.C(n_1591),
.D(n_1647),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2361),
.B(n_1612),
.Y(n_2383)
);

XNOR2xp5_ASAP7_75t_L g2384 ( 
.A(n_2360),
.B(n_1647),
.Y(n_2384)
);

AOI221xp5_ASAP7_75t_L g2385 ( 
.A1(n_2369),
.A2(n_2378),
.B1(n_2372),
.B2(n_2371),
.C(n_2363),
.Y(n_2385)
);

OAI221xp5_ASAP7_75t_SL g2386 ( 
.A1(n_2376),
.A2(n_2374),
.B1(n_2365),
.B2(n_2364),
.C(n_2373),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2368),
.B(n_1612),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2375),
.Y(n_2388)
);

OAI21xp33_ASAP7_75t_L g2389 ( 
.A1(n_2357),
.A2(n_1718),
.B(n_1647),
.Y(n_2389)
);

NAND5xp2_ASAP7_75t_L g2390 ( 
.A(n_2379),
.B(n_1582),
.C(n_1635),
.D(n_1750),
.E(n_1653),
.Y(n_2390)
);

OAI322xp33_ASAP7_75t_L g2391 ( 
.A1(n_2377),
.A2(n_1618),
.A3(n_1617),
.B1(n_1644),
.B2(n_1620),
.C1(n_1632),
.C2(n_1649),
.Y(n_2391)
);

NAND4xp25_ASAP7_75t_L g2392 ( 
.A(n_2367),
.B(n_1653),
.C(n_1635),
.D(n_1621),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_2366),
.A2(n_2362),
.B1(n_2370),
.B2(n_1635),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2358),
.B(n_1632),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2358),
.Y(n_2395)
);

AOI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_2360),
.A2(n_1620),
.B(n_1644),
.Y(n_2396)
);

A2O1A1Ixp33_ASAP7_75t_SL g2397 ( 
.A1(n_2358),
.A2(n_1620),
.B(n_1644),
.C(n_1618),
.Y(n_2397)
);

OAI221xp5_ASAP7_75t_L g2398 ( 
.A1(n_2359),
.A2(n_1638),
.B1(n_1646),
.B2(n_1641),
.C(n_1649),
.Y(n_2398)
);

OAI22xp33_ASAP7_75t_L g2399 ( 
.A1(n_2393),
.A2(n_1605),
.B1(n_1617),
.B2(n_1638),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2384),
.B(n_1750),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2395),
.B(n_1750),
.Y(n_2401)
);

OAI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2385),
.A2(n_1641),
.B(n_1646),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2386),
.A2(n_2388),
.B(n_2383),
.Y(n_2403)
);

A2O1A1Ixp33_ASAP7_75t_L g2404 ( 
.A1(n_2389),
.A2(n_1637),
.B(n_1663),
.C(n_1679),
.Y(n_2404)
);

NAND4xp25_ASAP7_75t_L g2405 ( 
.A(n_2394),
.B(n_1621),
.C(n_1599),
.D(n_1663),
.Y(n_2405)
);

AOI221xp5_ASAP7_75t_L g2406 ( 
.A1(n_2398),
.A2(n_1685),
.B1(n_1679),
.B2(n_1637),
.C(n_1693),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2387),
.Y(n_2407)
);

NAND3xp33_ASAP7_75t_L g2408 ( 
.A(n_2396),
.B(n_1685),
.C(n_1695),
.Y(n_2408)
);

BUFx2_ASAP7_75t_L g2409 ( 
.A(n_2392),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2409),
.Y(n_2410)
);

NAND2x1p5_ASAP7_75t_L g2411 ( 
.A(n_2403),
.B(n_2382),
.Y(n_2411)
);

AND2x4_ASAP7_75t_L g2412 ( 
.A(n_2402),
.B(n_2381),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2407),
.B(n_2380),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2399),
.B(n_2397),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_SL g2415 ( 
.A(n_2401),
.B(n_2400),
.C(n_2404),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2408),
.A2(n_2405),
.B1(n_2406),
.B2(n_2390),
.Y(n_2416)
);

AOI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_2403),
.A2(n_2391),
.B(n_1599),
.Y(n_2417)
);

XNOR2xp5_ASAP7_75t_L g2418 ( 
.A(n_2409),
.B(n_1637),
.Y(n_2418)
);

AOI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2399),
.A2(n_1695),
.B1(n_1693),
.B2(n_1750),
.C(n_1528),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2418),
.Y(n_2420)
);

NAND3xp33_ASAP7_75t_L g2421 ( 
.A(n_2413),
.B(n_134),
.C(n_164),
.Y(n_2421)
);

OR2x2_ASAP7_75t_L g2422 ( 
.A(n_2410),
.B(n_1750),
.Y(n_2422)
);

INVx1_ASAP7_75t_SL g2423 ( 
.A(n_2412),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2411),
.B(n_1656),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2416),
.A2(n_1656),
.B1(n_1674),
.B2(n_1704),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2417),
.B(n_1717),
.Y(n_2426)
);

NOR2x1_ASAP7_75t_L g2427 ( 
.A(n_2415),
.B(n_150),
.Y(n_2427)
);

OR2x2_ASAP7_75t_L g2428 ( 
.A(n_2414),
.B(n_1656),
.Y(n_2428)
);

NOR5xp2_ASAP7_75t_L g2429 ( 
.A(n_2421),
.B(n_2419),
.C(n_1656),
.D(n_1704),
.E(n_1674),
.Y(n_2429)
);

AND3x2_ASAP7_75t_L g2430 ( 
.A(n_2420),
.B(n_201),
.C(n_200),
.Y(n_2430)
);

NAND3xp33_ASAP7_75t_L g2431 ( 
.A(n_2427),
.B(n_164),
.C(n_150),
.Y(n_2431)
);

AOI221x1_ASAP7_75t_L g2432 ( 
.A1(n_2426),
.A2(n_150),
.B1(n_200),
.B2(n_174),
.C(n_199),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2422),
.Y(n_2433)
);

NOR3xp33_ASAP7_75t_L g2434 ( 
.A(n_2423),
.B(n_2428),
.C(n_2424),
.Y(n_2434)
);

NAND4xp25_ASAP7_75t_L g2435 ( 
.A(n_2425),
.B(n_150),
.C(n_200),
.D(n_199),
.Y(n_2435)
);

OAI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2423),
.A2(n_150),
.B(n_164),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2433),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2434),
.B(n_1656),
.Y(n_2438)
);

BUFx3_ASAP7_75t_L g2439 ( 
.A(n_2431),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2430),
.B(n_1656),
.Y(n_2440)
);

OAI22x1_ASAP7_75t_L g2441 ( 
.A1(n_2437),
.A2(n_2438),
.B1(n_2440),
.B2(n_2439),
.Y(n_2441)
);

AOI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2437),
.A2(n_2435),
.B1(n_2436),
.B2(n_2429),
.Y(n_2442)
);

AOI22xp33_ASAP7_75t_L g2443 ( 
.A1(n_2441),
.A2(n_2432),
.B1(n_150),
.B2(n_164),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2443),
.A2(n_2442),
.B1(n_164),
.B2(n_150),
.Y(n_2444)
);

OAI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_2444),
.A2(n_164),
.B1(n_150),
.B2(n_1656),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2445),
.A2(n_164),
.B1(n_150),
.B2(n_1674),
.Y(n_2446)
);

XOR2xp5_ASAP7_75t_L g2447 ( 
.A(n_2446),
.B(n_164),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2447),
.B(n_164),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2448),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2449),
.B(n_164),
.Y(n_2450)
);

AOI221xp5_ASAP7_75t_L g2451 ( 
.A1(n_2450),
.A2(n_164),
.B1(n_1674),
.B2(n_1704),
.C(n_1717),
.Y(n_2451)
);

AOI211xp5_ASAP7_75t_L g2452 ( 
.A1(n_2451),
.A2(n_164),
.B(n_1704),
.C(n_1674),
.Y(n_2452)
);


endmodule