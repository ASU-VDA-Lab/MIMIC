module real_jpeg_24630_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_35),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_84),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_84),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_84),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_33),
.B1(n_53),
.B2(n_54),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_33),
.B1(n_65),
.B2(n_66),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_22),
.B1(n_25),
.B2(n_33),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_6),
.B(n_21),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_6),
.A2(n_25),
.B(n_91),
.C(n_241),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_6),
.A2(n_22),
.B1(n_25),
.B2(n_179),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_6),
.B(n_54),
.C(n_69),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_179),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_6),
.A2(n_51),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_6),
.B(n_134),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_7),
.A2(n_64),
.B1(n_85),
.B2(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_35),
.B1(n_40),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_8),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_22),
.B1(n_25),
.B2(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_80),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_9),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_9),
.A2(n_29),
.B1(n_40),
.B2(n_170),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_170),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_170),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_11),
.A2(n_40),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_11),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_22),
.B1(n_25),
.B2(n_118),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_118),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_118),
.Y(n_269)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_13),
.A2(n_22),
.B1(n_25),
.B2(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_13),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_95),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_13),
.A2(n_40),
.B1(n_95),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_95),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_14),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_14),
.A2(n_22),
.B1(n_25),
.B2(n_39),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_16),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_16),
.A2(n_52),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_16),
.Y(n_201)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_16),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_16),
.A2(n_52),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_32),
.Y(n_20)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_27),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_21),
.A2(n_27),
.B1(n_117),
.B2(n_210),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_21),
.A2(n_27),
.B1(n_38),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx5_ASAP7_75t_SL g25 ( 
.A(n_22),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_22),
.A2(n_25),
.B1(n_91),
.B2(n_92),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_22),
.A2(n_26),
.B(n_180),
.C(n_190),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g190 ( 
.A(n_24),
.B(n_25),
.C(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_27),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_27),
.A2(n_122),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_29),
.Y(n_191)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_31),
.A2(n_79),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_31),
.B(n_83),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_31),
.A2(n_79),
.B1(n_120),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_31),
.A2(n_120),
.B1(n_142),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_31),
.A2(n_81),
.B(n_209),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_34),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_37),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_37),
.B(n_356),
.Y(n_357)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_40),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_355),
.B(n_357),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_343),
.B(n_354),
.Y(n_44)
);

OAI31xp33_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_145),
.A3(n_159),
.B(n_340),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_123),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_47),
.B(n_123),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_86),
.C(n_102),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_48),
.A2(n_86),
.B1(n_87),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_48),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_75),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_50),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_50),
.A2(n_61),
.B1(n_62),
.B2(n_76),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_58),
.B(n_60),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_51),
.A2(n_60),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_51),
.A2(n_186),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_51),
.A2(n_107),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_51),
.A2(n_269),
.B(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_52),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_54),
.B1(n_69),
.B2(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_53),
.B(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_67),
.B1(n_74),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_66),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_65),
.B(n_261),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_66),
.A2(n_92),
.B(n_179),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_67),
.A2(n_74),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_67),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_67),
.A2(n_74),
.B1(n_236),
.B2(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_72),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_72),
.A2(n_98),
.B1(n_112),
.B2(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_72),
.B(n_179),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_72),
.A2(n_175),
.B(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_74),
.B(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_85),
.B(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B(n_101),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_89),
.A2(n_90),
.B1(n_136),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_89),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_89),
.A2(n_207),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_90),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_90),
.A2(n_114),
.B(n_195),
.Y(n_319)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_98),
.A2(n_235),
.B(n_237),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_98),
.A2(n_237),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_102),
.A2(n_103),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.C(n_115),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_104),
.A2(n_105),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_106),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_108),
.B(n_179),
.Y(n_273)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_108),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_108),
.A2(n_243),
.B(n_267),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_113),
.B(n_115),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B(n_121),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_126),
.C(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_141),
.B2(n_144),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_138),
.C(n_141),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_134),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_133),
.A2(n_134),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_134),
.B(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_138),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_138),
.B(n_152),
.C(n_156),
.Y(n_353)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_144),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_141),
.B(n_148),
.C(n_151),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_146),
.A2(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_158),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_147),
.B(n_158),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_153),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_157),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_333),
.B(n_339),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_323),
.B(n_332),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_222),
.B(n_306),
.C(n_322),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_202),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_163),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_181),
.C(n_192),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_164),
.A2(n_165),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_173),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_172),
.C(n_177),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_181),
.A2(n_182),
.B1(n_192),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_188),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_192),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.C(n_199),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_201),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_211),
.B1(n_212),
.B2(n_221),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_203),
.Y(n_358)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.CI(n_208),
.CON(n_203),
.SN(n_203)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_204),
.B(n_205),
.C(n_208),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_220),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_213),
.B(n_220),
.C(n_221),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_214),
.B(n_219),
.Y(n_320)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_299),
.B(n_305),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_254),
.B(n_298),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_246),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_227),
.B(n_246),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_245),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_234),
.C(n_238),
.Y(n_304)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.C(n_251),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_248),
.A2(n_251),
.B1(n_252),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_292),
.B(n_297),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_282),
.B(n_291),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_270),
.B(n_281),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_265),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_277),
.B(n_280),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_279),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_290),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_296),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_321),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_318),
.C(n_320),
.Y(n_331)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_328),
.C(n_331),
.Y(n_338)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_338),
.Y(n_339)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_345),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_353),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_349),
.B1(n_351),
.B2(n_352),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_347),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_349),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_351),
.C(n_353),
.Y(n_356)
);


endmodule