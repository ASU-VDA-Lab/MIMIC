module fake_jpeg_21942_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_16),
.A2(n_17),
.B(n_28),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_34),
.A2(n_18),
.B(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_42),
.Y(n_70)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_15),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_27),
.B1(n_31),
.B2(n_15),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_32),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_72),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_25),
.Y(n_100)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_36),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_87),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_22),
.B1(n_25),
.B2(n_21),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_58),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_89),
.CI(n_29),
.CON(n_106),
.SN(n_106)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_5),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_5),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_6),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_50),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_54),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_66),
.B1(n_63),
.B2(n_47),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_103),
.B1(n_48),
.B2(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_111),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_63),
.B1(n_53),
.B2(n_60),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_109),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_110),
.B1(n_90),
.B2(n_23),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_6),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_93),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_7),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_85),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_122),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_77),
.B(n_75),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_75),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_96),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_128),
.B1(n_112),
.B2(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_113),
.C(n_83),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NOR4xp25_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_107),
.C(n_111),
.D(n_70),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_133),
.B(n_135),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_108),
.B(n_88),
.C(n_106),
.D(n_109),
.Y(n_133)
);

XOR2x2_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_108),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_117),
.C(n_119),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_144),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_142),
.B1(n_129),
.B2(n_128),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_107),
.B1(n_89),
.B2(n_82),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_96),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_106),
.B(n_114),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_148),
.B(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_97),
.Y(n_149)
);

OA21x2_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_152),
.B(n_154),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_142),
.B1(n_140),
.B2(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_141),
.B1(n_138),
.B2(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_157),
.B1(n_146),
.B2(n_142),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_159),
.B(n_160),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_140),
.C(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_125),
.C(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_165),
.B1(n_167),
.B2(n_155),
.Y(n_169)
);

AOI31xp67_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_158),
.A3(n_157),
.B(n_142),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_168),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_94),
.B(n_100),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_7),
.B(n_8),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_172),
.A3(n_170),
.B1(n_94),
.B2(n_76),
.C1(n_10),
.C2(n_11),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_100),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_115),
.A3(n_94),
.B1(n_11),
.B2(n_12),
.C1(n_9),
.C2(n_8),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_7),
.B(n_9),
.C(n_171),
.D(n_177),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_9),
.Y(n_179)
);


endmodule