module fake_netlist_6_1806_n_1912 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1912);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1912;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_1328;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx2_ASAP7_75t_L g494 ( 
.A(n_22),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_440),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_136),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_64),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_35),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_276),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_398),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_33),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_95),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_73),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_75),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_327),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_331),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_22),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_287),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_370),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_27),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_380),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_436),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_445),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_264),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_412),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_153),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_113),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_394),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_201),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_322),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_194),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_97),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_234),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_369),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_4),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_239),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_473),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_416),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_158),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_302),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_27),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_53),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_157),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_97),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_38),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_39),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_379),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_240),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_346),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_282),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_213),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_487),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_249),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_364),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_156),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_168),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_152),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_463),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_182),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_170),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_105),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_43),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_205),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_154),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_127),
.Y(n_557)
);

BUFx5_ASAP7_75t_L g558 ( 
.A(n_7),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_345),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_43),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_68),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_167),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_326),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_474),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_116),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_363),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_210),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_247),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_203),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_230),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_244),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_35),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_200),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_148),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_298),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_1),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_207),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_403),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_344),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_491),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_428),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_144),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_32),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_17),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_427),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_144),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_392),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_260),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_92),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_317),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_29),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_14),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_53),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_389),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_242),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_133),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_378),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_356),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_384),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_489),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_484),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_10),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_254),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_353),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_1),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_180),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_371),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_442),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_166),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_88),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_4),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_3),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_236),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_146),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_30),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_426),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_393),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_289),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_215),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_446),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_128),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_156),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_175),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_0),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_404),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_250),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_259),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_24),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_166),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_305),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_406),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_263),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_74),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_112),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_439),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_79),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_437),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_311),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_377),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_350),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_402),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_209),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_401),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_135),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_470),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_340),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_252),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_231),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_158),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_78),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_256),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_455),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_400),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_58),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_409),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_390),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_64),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_162),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_202),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_181),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_160),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_270),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_307),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_124),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_359),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_55),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_199),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_60),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_160),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_15),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_90),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_89),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_255),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_104),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_486),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_20),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_60),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_89),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_397),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_348),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_170),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_6),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_235),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_195),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_24),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_104),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_241),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_172),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

INVxp33_ASAP7_75t_SL g692 ( 
.A(n_494),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_558),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_495),
.Y(n_694)
);

INVxp33_ASAP7_75t_SL g695 ( 
.A(n_498),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_558),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_502),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_558),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_558),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_549),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_508),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_645),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_508),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_659),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_590),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_673),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_616),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_502),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_581),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_598),
.B(n_0),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_553),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_553),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_686),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_686),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_686),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_556),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_686),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_556),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_565),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_687),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_499),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_687),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_581),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_687),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_687),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_503),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_497),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_524),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_527),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_531),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_514),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_534),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_537),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_660),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_496),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_637),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_506),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_504),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_565),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_573),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_585),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_593),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_683),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_594),
.Y(n_745)
);

INVxp33_ASAP7_75t_SL g746 ( 
.A(n_505),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_608),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_614),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_538),
.Y(n_749)
);

INVxp33_ASAP7_75t_L g750 ( 
.A(n_497),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_617),
.Y(n_751)
);

INVxp33_ASAP7_75t_L g752 ( 
.A(n_626),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_631),
.Y(n_753)
);

CKINVDCx16_ASAP7_75t_R g754 ( 
.A(n_564),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_635),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_511),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_656),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_662),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_663),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_670),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_510),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_518),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_676),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_533),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_637),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_688),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_690),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_536),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_500),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_507),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_528),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_509),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_515),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_592),
.Y(n_774)
);

INVxp33_ASAP7_75t_SL g775 ( 
.A(n_548),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_516),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_525),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_694),
.B(n_513),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_721),
.Y(n_779)
);

BUFx12f_ASAP7_75t_L g780 ( 
.A(n_701),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_722),
.B(n_517),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_721),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_710),
.B(n_519),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_714),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_691),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_715),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_716),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_707),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_693),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_718),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_707),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_738),
.B(n_761),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_723),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_692),
.A2(n_550),
.B1(n_574),
.B2(n_501),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_725),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_SL g797 ( 
.A1(n_698),
.A2(n_611),
.B1(n_666),
.B2(n_592),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_696),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_726),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_737),
.B(n_598),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_732),
.B(n_528),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_765),
.B(n_579),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_699),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_746),
.B(n_521),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_700),
.Y(n_806)
);

INVx5_ASAP7_75t_L g807 ( 
.A(n_728),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_746),
.B(n_571),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_728),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_753),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_753),
.Y(n_811)
);

XNOR2x2_ASAP7_75t_L g812 ( 
.A(n_749),
.B(n_604),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_769),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_724),
.B(n_523),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_770),
.A2(n_629),
.B(n_605),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_724),
.B(n_629),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_768),
.B(n_599),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_772),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_773),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_776),
.A2(n_605),
.B(n_541),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_692),
.A2(n_550),
.B1(n_574),
.B2(n_501),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_777),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_727),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_729),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_730),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_754),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_750),
.B(n_547),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_736),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_731),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_703),
.B(n_541),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_733),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_734),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_771),
.Y(n_833)
);

BUFx8_ASAP7_75t_L g834 ( 
.A(n_708),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_801),
.B(n_711),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_827),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_786),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_827),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_823),
.Y(n_839)
);

INVxp33_ASAP7_75t_L g840 ( 
.A(n_814),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_805),
.B(n_817),
.C(n_808),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_786),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_798),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_790),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_800),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_804),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_830),
.A2(n_695),
.B1(n_671),
.B2(n_706),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_804),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_833),
.B(n_756),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_833),
.B(n_762),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_SL g851 ( 
.A(n_784),
.B(n_611),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_779),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_803),
.A2(n_695),
.B1(n_775),
.B2(n_768),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_779),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_822),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_783),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_834),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_798),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_778),
.B(n_775),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_783),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_798),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_809),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_816),
.A2(n_529),
.B(n_526),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_814),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_809),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_806),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_784),
.B(n_764),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_806),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_801),
.B(n_739),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_781),
.B(n_641),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_832),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_793),
.B(n_641),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_806),
.Y(n_873)
);

AND3x2_ASAP7_75t_L g874 ( 
.A(n_782),
.B(n_744),
.C(n_675),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_825),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_788),
.Y(n_876)
);

INVxp33_ASAP7_75t_L g877 ( 
.A(n_795),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_822),
.B(n_739),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_813),
.B(n_512),
.Y(n_879)
);

BUFx10_ASAP7_75t_L g880 ( 
.A(n_826),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_788),
.Y(n_881)
);

NOR2x1p5_ASAP7_75t_L g882 ( 
.A(n_826),
.B(n_771),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_822),
.B(n_582),
.Y(n_883)
);

BUFx6f_ASAP7_75t_SL g884 ( 
.A(n_825),
.Y(n_884)
);

BUFx6f_ASAP7_75t_SL g885 ( 
.A(n_829),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_822),
.B(n_644),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_788),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_829),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_813),
.B(n_520),
.Y(n_889)
);

AND2x6_ASAP7_75t_L g890 ( 
.A(n_813),
.B(n_644),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_822),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_788),
.Y(n_892)
);

BUFx6f_ASAP7_75t_SL g893 ( 
.A(n_810),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_788),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_785),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_832),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_789),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_832),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_832),
.B(n_675),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_807),
.Y(n_900)
);

INVxp33_ASAP7_75t_SL g901 ( 
.A(n_821),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_832),
.Y(n_902)
);

AND3x2_ASAP7_75t_L g903 ( 
.A(n_782),
.B(n_792),
.C(n_735),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_785),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_787),
.Y(n_905)
);

INVx8_ASAP7_75t_L g906 ( 
.A(n_780),
.Y(n_906)
);

NOR2x1p5_ASAP7_75t_L g907 ( 
.A(n_780),
.B(n_535),
.Y(n_907)
);

INVxp33_ASAP7_75t_SL g908 ( 
.A(n_797),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_824),
.B(n_582),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_824),
.B(n_522),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_820),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_875),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_888),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_911),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_839),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_895),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_841),
.B(n_828),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_835),
.B(n_820),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_904),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_904),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_843),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_862),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_905),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_905),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_849),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_859),
.B(n_705),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_843),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_864),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_836),
.B(n_818),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_906),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_906),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_859),
.B(n_828),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_840),
.B(n_792),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_862),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_852),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_865),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_854),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_879),
.B(n_824),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_850),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_856),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_837),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_856),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_860),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_860),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_855),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_858),
.Y(n_947)
);

AND2x6_ASAP7_75t_L g948 ( 
.A(n_911),
.B(n_582),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_840),
.B(n_802),
.Y(n_949)
);

AO21x1_ASAP7_75t_L g950 ( 
.A1(n_872),
.A2(n_539),
.B(n_532),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_869),
.B(n_698),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_842),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_867),
.B(n_750),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_861),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_866),
.B(n_831),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_838),
.B(n_709),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_868),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_873),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_906),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_897),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_880),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_842),
.Y(n_962)
);

XNOR2xp5_ASAP7_75t_L g963 ( 
.A(n_901),
.B(n_709),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_874),
.Y(n_964)
);

XOR2x2_ASAP7_75t_L g965 ( 
.A(n_908),
.B(n_901),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_844),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_844),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_872),
.B(n_717),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_845),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_846),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_848),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_909),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_909),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_877),
.B(n_752),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_886),
.Y(n_975)
);

INVx8_ASAP7_75t_L g976 ( 
.A(n_884),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_886),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_899),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_877),
.B(n_752),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_870),
.A2(n_815),
.B(n_546),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_878),
.B(n_702),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_878),
.B(n_882),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_891),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_896),
.Y(n_984)
);

AND2x2_ASAP7_75t_SL g985 ( 
.A(n_857),
.B(n_812),
.Y(n_985)
);

INVxp67_ASAP7_75t_SL g986 ( 
.A(n_855),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_898),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_880),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_902),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_870),
.B(n_831),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_907),
.B(n_819),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_876),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_880),
.B(n_704),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_884),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_853),
.B(n_717),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_881),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_903),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_889),
.B(n_712),
.Y(n_998)
);

BUFx6f_ASAP7_75t_SL g999 ( 
.A(n_908),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_881),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_871),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_890),
.B(n_831),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_851),
.B(n_812),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_892),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_910),
.B(n_713),
.Y(n_1005)
);

OR2x2_ASAP7_75t_SL g1006 ( 
.A(n_847),
.B(n_719),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_894),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_894),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_863),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_885),
.B(n_552),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_885),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_890),
.B(n_819),
.Y(n_1012)
);

INVxp33_ASAP7_75t_L g1013 ( 
.A(n_893),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_893),
.Y(n_1014)
);

INVxp33_ASAP7_75t_L g1015 ( 
.A(n_855),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_890),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_890),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_890),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_855),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_887),
.B(n_741),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_887),
.B(n_742),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_887),
.B(n_719),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_883),
.A2(n_559),
.B(n_545),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_883),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_900),
.Y(n_1025)
);

AO22x1_ASAP7_75t_L g1026 ( 
.A1(n_932),
.A2(n_834),
.B1(n_554),
.B2(n_560),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_926),
.B(n_720),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_981),
.B(n_572),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_925),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_930),
.Y(n_1030)
);

OAI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_974),
.A2(n_562),
.B1(n_575),
.B2(n_561),
.C(n_551),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_998),
.B(n_576),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_986),
.A2(n_900),
.B(n_807),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1003),
.A2(n_586),
.B1(n_615),
.B2(n_589),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1005),
.B(n_628),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_975),
.A2(n_634),
.B1(n_639),
.B2(n_632),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_SL g1037 ( 
.A1(n_963),
.A2(n_740),
.B1(n_774),
.B2(n_666),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_921),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_974),
.A2(n_642),
.B1(n_643),
.B2(n_640),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_953),
.B(n_650),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1020),
.B(n_653),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_914),
.B(n_912),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_933),
.B(n_740),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_931),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_914),
.B(n_913),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_L g1046 ( 
.A(n_959),
.B(n_743),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_921),
.B(n_811),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_960),
.Y(n_1048)
);

AND2x6_ASAP7_75t_SL g1049 ( 
.A(n_995),
.B(n_745),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1018),
.A2(n_655),
.B1(n_661),
.B2(n_654),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_940),
.B(n_669),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_949),
.A2(n_685),
.B(n_815),
.C(n_791),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_979),
.B(n_787),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_986),
.B(n_791),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_929),
.B(n_794),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_929),
.B(n_834),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_982),
.B(n_530),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_927),
.B(n_794),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_968),
.A2(n_799),
.B(n_796),
.C(n_542),
.Y(n_1059)
);

AO21x1_ASAP7_75t_L g1060 ( 
.A1(n_918),
.A2(n_799),
.B(n_796),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_SL g1061 ( 
.A(n_961),
.B(n_774),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_915),
.B(n_540),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_SL g1063 ( 
.A(n_951),
.B(n_583),
.C(n_577),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_917),
.B(n_584),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_L g1065 ( 
.A(n_988),
.B(n_747),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1021),
.B(n_543),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_1021),
.B(n_811),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_916),
.B(n_544),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_976),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_976),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_977),
.A2(n_603),
.B1(n_582),
.B2(n_667),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_919),
.B(n_555),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_920),
.B(n_563),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_976),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_993),
.B(n_566),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_1018),
.B(n_567),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_978),
.A2(n_603),
.B1(n_667),
.B2(n_568),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_923),
.B(n_569),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_942),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_924),
.B(n_947),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_954),
.B(n_570),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_928),
.B(n_748),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_969),
.B(n_578),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_970),
.B(n_580),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_928),
.B(n_587),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_950),
.A2(n_603),
.B1(n_588),
.B2(n_595),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_946),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_971),
.B(n_591),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_938),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_952),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1022),
.B(n_557),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_918),
.A2(n_600),
.B1(n_601),
.B2(n_596),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_991),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_941),
.A2(n_602),
.B1(n_609),
.B2(n_606),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_1009),
.A2(n_810),
.B(n_755),
.C(n_757),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_956),
.B(n_597),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1006),
.B(n_607),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_990),
.B(n_610),
.Y(n_1099)
);

NAND2x1_ASAP7_75t_L g1100 ( 
.A(n_957),
.B(n_751),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_991),
.B(n_618),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_990),
.B(n_619),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_948),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1010),
.B(n_684),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_943),
.B(n_620),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_985),
.B(n_612),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_944),
.B(n_621),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_939),
.B(n_622),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_964),
.Y(n_1109)
);

NOR2x1p5_ASAP7_75t_L g1110 ( 
.A(n_994),
.B(n_613),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1010),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_994),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_966),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_967),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_945),
.A2(n_633),
.B1(n_647),
.B2(n_627),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_972),
.A2(n_649),
.B1(n_657),
.B2(n_648),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_958),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_962),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_L g1119 ( 
.A(n_997),
.B(n_758),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1010),
.B(n_684),
.Y(n_1120)
);

AND2x6_ASAP7_75t_SL g1121 ( 
.A(n_999),
.B(n_759),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_1014),
.Y(n_1122)
);

AND2x6_ASAP7_75t_SL g1123 ( 
.A(n_999),
.B(n_760),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_973),
.A2(n_664),
.B1(n_665),
.B2(n_658),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_922),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1011),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_955),
.A2(n_980),
.B(n_1016),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_936),
.B(n_677),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_L g1129 ( 
.A(n_1012),
.B(n_766),
.C(n_763),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1002),
.A2(n_807),
.B(n_682),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1012),
.B(n_681),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1013),
.B(n_623),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_965),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1002),
.A2(n_767),
.B(n_689),
.C(n_625),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_937),
.A2(n_984),
.B1(n_987),
.B2(n_983),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_992),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_989),
.B(n_1024),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_996),
.A2(n_630),
.B1(n_636),
.B2(n_624),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1001),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1000),
.A2(n_646),
.B1(n_651),
.B2(n_638),
.Y(n_1140)
);

CKINVDCx16_ASAP7_75t_R g1141 ( 
.A(n_980),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1019),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1004),
.B(n_652),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_948),
.B(n_668),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1017),
.A2(n_674),
.B1(n_678),
.B2(n_672),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_948),
.A2(n_1023),
.B1(n_1025),
.B2(n_1015),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_925),
.B(n_679),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_932),
.A2(n_680),
.B1(n_807),
.B2(n_206),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_981),
.B(n_807),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_935),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_981),
.B(n_2),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_935),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_925),
.B(n_204),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_981),
.B(n_2),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_925),
.B(n_208),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_953),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_981),
.B(n_3),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_925),
.B(n_211),
.Y(n_1159)
);

BUFx8_ASAP7_75t_L g1160 ( 
.A(n_999),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_961),
.B(n_212),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_932),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_921),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_935),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_981),
.B(n_8),
.Y(n_1165)
);

AND2x6_ASAP7_75t_SL g1166 ( 
.A(n_995),
.B(n_8),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_981),
.B(n_9),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_960),
.Y(n_1168)
);

NAND2x1_ASAP7_75t_L g1169 ( 
.A(n_946),
.B(n_214),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_981),
.B(n_9),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_925),
.B(n_216),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_981),
.B(n_10),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_929),
.B(n_217),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_935),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_L g1175 ( 
.A(n_932),
.B(n_11),
.C(n_12),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_930),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_932),
.A2(n_219),
.B1(n_220),
.B2(n_218),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_981),
.B(n_11),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_932),
.B(n_12),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_932),
.B(n_13),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_934),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_953),
.B(n_14),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_925),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_981),
.B(n_15),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_932),
.B(n_16),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_932),
.B(n_16),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_925),
.B(n_221),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_R g1188 ( 
.A(n_1126),
.B(n_222),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1183),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1071),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1157),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_1160),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1042),
.B(n_1045),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1068),
.Y(n_1194)
);

OR2x2_ASAP7_75t_SL g1195 ( 
.A(n_1063),
.B(n_18),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1029),
.B(n_223),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1118),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1094),
.B(n_224),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1173),
.B(n_225),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1173),
.B(n_226),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1163),
.Y(n_1201)
);

AOI222xp33_ASAP7_75t_L g1202 ( 
.A1(n_1037),
.A2(n_1106),
.B1(n_1027),
.B2(n_1043),
.C1(n_1180),
.C2(n_1179),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1121),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1181),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1160),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1083),
.B(n_18),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1075),
.B(n_19),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1070),
.B(n_227),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1117),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1048),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1080),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1092),
.B(n_19),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1163),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1030),
.Y(n_1214)
);

AOI211xp5_ASAP7_75t_L g1215 ( 
.A1(n_1098),
.A2(n_1064),
.B(n_1186),
.C(n_1185),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1109),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1163),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1141),
.A2(n_229),
.B1(n_232),
.B2(n_228),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1070),
.B(n_233),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1070),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1090),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1053),
.B(n_21),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1088),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1182),
.B(n_23),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1086),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1097),
.B(n_23),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1028),
.B(n_25),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1044),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1176),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1040),
.B(n_1032),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1168),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1061),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1142),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1111),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1055),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1091),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1104),
.Y(n_1237)
);

CKINVDCx14_ASAP7_75t_R g1238 ( 
.A(n_1112),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1065),
.B(n_25),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1151),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1088),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1056),
.B(n_26),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1140),
.B(n_26),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1153),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1035),
.B(n_28),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1122),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1133),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1152),
.B(n_28),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1049),
.Y(n_1249)
);

CKINVDCx6p67_ASAP7_75t_R g1250 ( 
.A(n_1120),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1113),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1142),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1155),
.B(n_1158),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1165),
.B(n_29),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1137),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1142),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1144),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1164),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1119),
.B(n_237),
.Y(n_1259)
);

OR2x4_ASAP7_75t_L g1260 ( 
.A(n_1132),
.B(n_30),
.Y(n_1260)
);

BUFx10_ASAP7_75t_L g1261 ( 
.A(n_1110),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1148),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1038),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1174),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1140),
.B(n_31),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1123),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1167),
.B(n_31),
.Y(n_1267)
);

NOR3xp33_ASAP7_75t_SL g1268 ( 
.A(n_1031),
.B(n_32),
.C(n_33),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1170),
.B(n_34),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_1067),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1114),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1125),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1136),
.Y(n_1273)
);

NOR3xp33_ASAP7_75t_SL g1274 ( 
.A(n_1101),
.B(n_34),
.C(n_36),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1172),
.B(n_36),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1169),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1178),
.B(n_37),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1051),
.Y(n_1278)
);

AND3x2_ASAP7_75t_SL g1279 ( 
.A(n_1166),
.B(n_37),
.C(n_38),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1076),
.A2(n_243),
.B1(n_245),
.B2(n_238),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1081),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1139),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1184),
.B(n_246),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1096),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1100),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1127),
.A2(n_251),
.B(n_248),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1058),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1047),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1034),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1054),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1139),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1077),
.A2(n_257),
.B(n_253),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1041),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1099),
.B(n_1146),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1154),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_R g1297 ( 
.A(n_1145),
.B(n_1161),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1156),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1062),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1135),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1128),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1057),
.B(n_42),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_1046),
.B(n_44),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1039),
.B(n_44),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1175),
.B(n_45),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1159),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1069),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1039),
.B(n_45),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1082),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1073),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1066),
.B(n_1129),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1150),
.A2(n_261),
.B1(n_262),
.B2(n_258),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1074),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1171),
.B(n_265),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1079),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1105),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1084),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1085),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1187),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1059),
.B(n_46),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1107),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1116),
.B(n_1124),
.Y(n_1322)
);

NOR3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1050),
.B(n_47),
.C(n_48),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1089),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1116),
.B(n_49),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1026),
.B(n_50),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1036),
.B(n_50),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1093),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1095),
.B(n_51),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1102),
.B(n_1095),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1115),
.B(n_51),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1115),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1103),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1131),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1138),
.B(n_52),
.Y(n_1335)
);

NAND2x1_ASAP7_75t_L g1336 ( 
.A(n_1147),
.B(n_266),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1060),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1052),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1108),
.B(n_52),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1147),
.Y(n_1340)
);

AND3x1_ASAP7_75t_L g1341 ( 
.A(n_1162),
.B(n_54),
.C(n_55),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1177),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1149),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1134),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1078),
.B(n_56),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1072),
.B(n_57),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1130),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1087),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1033),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1286),
.A2(n_268),
.B(n_267),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1258),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1215),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1281),
.B(n_59),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1284),
.A2(n_1338),
.B(n_1336),
.Y(n_1355)
);

CKINVDCx6p67_ASAP7_75t_R g1356 ( 
.A(n_1220),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1230),
.A2(n_1193),
.B(n_1290),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1220),
.B(n_269),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1258),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1202),
.B(n_1225),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1294),
.A2(n_1322),
.B(n_1330),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_L g1362 ( 
.A1(n_1253),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1201),
.B(n_271),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1198),
.B(n_493),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1343),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1281),
.B(n_65),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1198),
.B(n_490),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1290),
.A2(n_273),
.B(n_272),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1337),
.A2(n_68),
.A3(n_66),
.B(n_67),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1293),
.A2(n_275),
.B(n_274),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1191),
.B(n_1317),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1255),
.B(n_67),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1292),
.A2(n_278),
.B(n_277),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1348),
.A2(n_280),
.B(n_279),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1235),
.B(n_69),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1342),
.A2(n_283),
.B(n_281),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1255),
.B(n_69),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1223),
.A2(n_285),
.B(n_284),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1307),
.A2(n_288),
.B(n_286),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1287),
.B(n_70),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1243),
.B(n_1265),
.Y(n_1381)
);

NOR2x1_ASAP7_75t_L g1382 ( 
.A(n_1201),
.B(n_290),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1190),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1315),
.A2(n_292),
.B(n_291),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1350),
.A2(n_488),
.B(n_294),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1257),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1386)
);

AOI211x1_ASAP7_75t_L g1387 ( 
.A1(n_1325),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1340),
.A2(n_295),
.B(n_293),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1241),
.A2(n_297),
.B(n_296),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1226),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1241),
.A2(n_300),
.B(n_299),
.Y(n_1391)
);

INVx5_ASAP7_75t_L g1392 ( 
.A(n_1333),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1257),
.A2(n_303),
.B(n_301),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1329),
.B(n_76),
.C(n_77),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1299),
.A2(n_306),
.B(n_304),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1333),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1220),
.Y(n_1397)
);

OA22x2_ASAP7_75t_L g1398 ( 
.A1(n_1242),
.A2(n_80),
.B1(n_77),
.B2(n_78),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1264),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1214),
.Y(n_1400)
);

AOI21xp33_ASAP7_75t_L g1401 ( 
.A1(n_1332),
.A2(n_81),
.B(n_82),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1301),
.A2(n_309),
.B(n_308),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1223),
.A2(n_312),
.B(n_310),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1318),
.B(n_82),
.Y(n_1404)
);

OAI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1331),
.A2(n_83),
.B(n_84),
.Y(n_1405)
);

OAI22x1_ASAP7_75t_L g1406 ( 
.A1(n_1335),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1295),
.B(n_85),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1334),
.A2(n_314),
.B(n_313),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1228),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1212),
.B(n_86),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1324),
.B(n_1278),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1283),
.A2(n_316),
.B(n_315),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1309),
.B(n_87),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1345),
.A2(n_319),
.B(n_318),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1310),
.A2(n_321),
.B(n_320),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1313),
.A2(n_1321),
.B(n_1300),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1248),
.A2(n_1267),
.B(n_1254),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1222),
.A2(n_324),
.B(n_323),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1231),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1272),
.A2(n_328),
.B(n_325),
.Y(n_1420)
);

AOI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1227),
.A2(n_330),
.B(n_329),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1246),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1316),
.B(n_91),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1213),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1264),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1273),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1200),
.A2(n_333),
.B(n_332),
.Y(n_1427)
);

AO31x2_ASAP7_75t_L g1428 ( 
.A1(n_1320),
.A2(n_93),
.A3(n_91),
.B(n_92),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1261),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1245),
.A2(n_335),
.B(n_334),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1271),
.A2(n_1273),
.B(n_1194),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1234),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1232),
.B(n_94),
.Y(n_1433)
);

INVx6_ASAP7_75t_SL g1434 ( 
.A(n_1261),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1199),
.A2(n_337),
.B(n_336),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1305),
.A2(n_94),
.B(n_95),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1349),
.A2(n_339),
.B(n_338),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1224),
.B(n_96),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1271),
.A2(n_342),
.B(n_341),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1289),
.A2(n_96),
.B(n_98),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1306),
.A2(n_347),
.B(n_343),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1311),
.A2(n_1344),
.B(n_1276),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1216),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1328),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1311),
.A2(n_351),
.B(n_349),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1262),
.B(n_352),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1204),
.A2(n_355),
.B(n_354),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1197),
.A2(n_358),
.B(n_357),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1200),
.B(n_99),
.Y(n_1449)
);

INVx8_ASAP7_75t_L g1450 ( 
.A(n_1213),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1285),
.A2(n_361),
.B(n_360),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1270),
.B(n_362),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1312),
.A2(n_366),
.B(n_365),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1206),
.B(n_101),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1209),
.A2(n_368),
.B(n_367),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1217),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_SL g1457 ( 
.A1(n_1304),
.A2(n_102),
.B(n_103),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1210),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1276),
.A2(n_1314),
.B(n_1298),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1221),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1229),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1275),
.B(n_106),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1277),
.A2(n_373),
.B(n_372),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1208),
.A2(n_375),
.B(n_374),
.Y(n_1464)
);

AOI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1240),
.A2(n_485),
.B(n_376),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1189),
.B(n_106),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1341),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.C(n_110),
.Y(n_1467)
);

OAI22x1_ASAP7_75t_L g1468 ( 
.A1(n_1326),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_1468)
);

AO31x2_ASAP7_75t_L g1469 ( 
.A1(n_1339),
.A2(n_111),
.A3(n_112),
.B(n_113),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1346),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_1470)
);

AND3x4_ASAP7_75t_L g1471 ( 
.A(n_1247),
.B(n_114),
.C(n_115),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1244),
.B(n_116),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1347),
.A2(n_117),
.A3(n_118),
.B(n_119),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1269),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1211),
.A2(n_382),
.B(n_381),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1205),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1239),
.B(n_120),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1268),
.A2(n_121),
.B(n_122),
.C(n_123),
.Y(n_1478)
);

AO21x1_ASAP7_75t_L g1479 ( 
.A1(n_1308),
.A2(n_124),
.B(n_125),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1314),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1237),
.B(n_383),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1319),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1296),
.A2(n_386),
.B(n_385),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1291),
.B(n_129),
.Y(n_1484)
);

INVx6_ASAP7_75t_L g1485 ( 
.A(n_1266),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1217),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_SL g1487 ( 
.A1(n_1280),
.A2(n_388),
.B(n_387),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1296),
.B(n_130),
.Y(n_1488)
);

OAI22x1_ASAP7_75t_L g1489 ( 
.A1(n_1302),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1296),
.B(n_131),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1208),
.B(n_391),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1298),
.B(n_132),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1195),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.C(n_137),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1327),
.A2(n_134),
.A3(n_137),
.B(n_138),
.Y(n_1494)
);

AND2x6_ASAP7_75t_L g1495 ( 
.A(n_1219),
.B(n_395),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1236),
.A2(n_399),
.B(n_396),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1263),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1251),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1355),
.A2(n_1351),
.B(n_1373),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1360),
.A2(n_1196),
.B1(n_1323),
.B2(n_1279),
.C(n_1274),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1357),
.A2(n_1219),
.B(n_1233),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1381),
.B(n_1242),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1353),
.A2(n_1303),
.B(n_1207),
.C(n_1259),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1425),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1491),
.B(n_1207),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_SL g1506 ( 
.A(n_1400),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1491),
.B(n_1333),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1361),
.A2(n_1252),
.B(n_1233),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1416),
.B(n_1282),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1352),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1442),
.A2(n_1256),
.B(n_1252),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1459),
.A2(n_1256),
.B(n_1252),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1463),
.A2(n_1405),
.B(n_1441),
.C(n_1440),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1422),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1430),
.A2(n_1218),
.B(n_1259),
.C(n_1256),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1359),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1375),
.B(n_1303),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1392),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1437),
.A2(n_1263),
.B(n_1288),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1399),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1475),
.A2(n_1263),
.B(n_1288),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1443),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1376),
.A2(n_1288),
.B(n_1260),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1392),
.Y(n_1524)
);

OAI21xp33_ASAP7_75t_L g1525 ( 
.A1(n_1394),
.A2(n_1249),
.B(n_1297),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1427),
.B(n_1203),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1436),
.A2(n_1250),
.B1(n_1238),
.B2(n_1192),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1426),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1432),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1383),
.B(n_1266),
.Y(n_1530)
);

CKINVDCx11_ASAP7_75t_R g1531 ( 
.A(n_1356),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1446),
.A2(n_1266),
.B1(n_1188),
.B2(n_140),
.Y(n_1532)
);

AO21x1_ASAP7_75t_L g1533 ( 
.A1(n_1388),
.A2(n_138),
.B(n_139),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1460),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1417),
.A2(n_139),
.B(n_140),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1429),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1411),
.B(n_141),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1371),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1364),
.B(n_142),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1395),
.A2(n_1415),
.B(n_1445),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1368),
.A2(n_483),
.B(n_417),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1364),
.B(n_143),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1393),
.A2(n_1374),
.B(n_1379),
.Y(n_1543)
);

AO32x2_ASAP7_75t_L g1544 ( 
.A1(n_1386),
.A2(n_145),
.A3(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1454),
.B(n_145),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1384),
.A2(n_482),
.B(n_418),
.Y(n_1546)
);

AO32x2_ASAP7_75t_L g1547 ( 
.A1(n_1444),
.A2(n_147),
.A3(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_L g1548 ( 
.A(n_1467),
.B(n_149),
.C(n_150),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1461),
.B(n_1458),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1402),
.A2(n_420),
.B(n_480),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1404),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1367),
.B(n_154),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1478),
.A2(n_155),
.B(n_157),
.C(n_159),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1419),
.A2(n_155),
.B1(n_159),
.B2(n_161),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1496),
.A2(n_423),
.B(n_479),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1409),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1370),
.A2(n_481),
.B(n_422),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1429),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1389),
.A2(n_476),
.B(n_421),
.Y(n_1559)
);

OAI22x1_ASAP7_75t_L g1560 ( 
.A1(n_1471),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1480),
.A2(n_163),
.B(n_164),
.C(n_165),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1482),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_1562)
);

O2A1O1Ixp5_ASAP7_75t_L g1563 ( 
.A1(n_1479),
.A2(n_169),
.B(n_171),
.C(n_172),
.Y(n_1563)
);

AO31x2_ASAP7_75t_L g1564 ( 
.A1(n_1390),
.A2(n_425),
.A3(n_472),
.B(n_471),
.Y(n_1564)
);

AO31x2_ASAP7_75t_L g1565 ( 
.A1(n_1391),
.A2(n_1406),
.A3(n_1474),
.B(n_1468),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1392),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1449),
.B(n_407),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1435),
.A2(n_169),
.B(n_171),
.C(n_173),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1365),
.A2(n_173),
.B(n_174),
.C(n_175),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1397),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1396),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1397),
.Y(n_1572)
);

BUFx12f_ASAP7_75t_L g1573 ( 
.A(n_1476),
.Y(n_1573)
);

INVx3_ASAP7_75t_SL g1574 ( 
.A(n_1485),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1367),
.B(n_174),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1490),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1462),
.B(n_176),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1396),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1354),
.B(n_177),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1366),
.B(n_178),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_SL g1581 ( 
.A1(n_1372),
.A2(n_179),
.B(n_180),
.C(n_181),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1447),
.A2(n_429),
.B(n_469),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1397),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1498),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1485),
.Y(n_1585)
);

O2A1O1Ixp5_ASAP7_75t_L g1586 ( 
.A1(n_1362),
.A2(n_179),
.B(n_182),
.C(n_183),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_SL g1587 ( 
.A1(n_1377),
.A2(n_1380),
.B(n_1488),
.C(n_1492),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1455),
.A2(n_430),
.B(n_468),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1407),
.B(n_183),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1497),
.B(n_408),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1431),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1453),
.A2(n_184),
.B(n_185),
.C(n_186),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1439),
.A2(n_431),
.B(n_467),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1489),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_1594)
);

BUFx12f_ASAP7_75t_L g1595 ( 
.A(n_1424),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_SL g1596 ( 
.A1(n_1472),
.A2(n_187),
.B(n_188),
.C(n_189),
.Y(n_1596)
);

BUFx4f_ASAP7_75t_L g1597 ( 
.A(n_1495),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1438),
.B(n_188),
.Y(n_1598)
);

AND2x2_ASAP7_75t_SL g1599 ( 
.A(n_1470),
.B(n_189),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1378),
.A2(n_433),
.B(n_466),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1452),
.B(n_432),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1424),
.Y(n_1602)
);

AO31x2_ASAP7_75t_L g1603 ( 
.A1(n_1483),
.A2(n_434),
.A3(n_465),
.B(n_464),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1450),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1477),
.B(n_190),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1396),
.B(n_424),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1423),
.B(n_190),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1369),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1413),
.B(n_191),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1401),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1434),
.Y(n_1611)
);

AO22x2_ASAP7_75t_L g1612 ( 
.A1(n_1387),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1410),
.B(n_1433),
.Y(n_1613)
);

AO31x2_ASAP7_75t_L g1614 ( 
.A1(n_1457),
.A2(n_1448),
.A3(n_1451),
.B(n_1465),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1369),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1412),
.A2(n_196),
.B(n_197),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1424),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1464),
.A2(n_447),
.B(n_410),
.Y(n_1618)
);

AO31x2_ASAP7_75t_L g1619 ( 
.A1(n_1414),
.A2(n_448),
.A3(n_411),
.B(n_413),
.Y(n_1619)
);

AOI21xp33_ASAP7_75t_L g1620 ( 
.A1(n_1493),
.A2(n_198),
.B(n_414),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1484),
.B(n_415),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1452),
.B(n_419),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1487),
.A2(n_475),
.B(n_435),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1403),
.A2(n_1408),
.B(n_1420),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1495),
.B(n_438),
.Y(n_1625)
);

AOI221x1_ASAP7_75t_L g1626 ( 
.A1(n_1487),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.C(n_449),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1513),
.A2(n_1398),
.B1(n_1481),
.B2(n_1466),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1599),
.A2(n_1363),
.B1(n_1382),
.B2(n_1358),
.Y(n_1628)
);

CKINVDCx11_ASAP7_75t_R g1629 ( 
.A(n_1573),
.Y(n_1629)
);

CKINVDCx6p67_ASAP7_75t_R g1630 ( 
.A(n_1574),
.Y(n_1630)
);

CKINVDCx11_ASAP7_75t_R g1631 ( 
.A(n_1531),
.Y(n_1631)
);

INVx6_ASAP7_75t_L g1632 ( 
.A(n_1595),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1597),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1548),
.A2(n_1525),
.B1(n_1533),
.B2(n_1562),
.Y(n_1634)
);

CKINVDCx6p67_ASAP7_75t_R g1635 ( 
.A(n_1514),
.Y(n_1635)
);

BUFx10_ASAP7_75t_L g1636 ( 
.A(n_1530),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1510),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1602),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1516),
.Y(n_1639)
);

INVx4_ASAP7_75t_SL g1640 ( 
.A(n_1526),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1536),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1529),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1520),
.Y(n_1643)
);

CKINVDCx11_ASAP7_75t_R g1644 ( 
.A(n_1526),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1612),
.A2(n_1469),
.B1(n_1450),
.B2(n_1494),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1538),
.A2(n_1486),
.B1(n_1456),
.B2(n_1434),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1609),
.A2(n_1456),
.B1(n_1486),
.B2(n_1469),
.Y(n_1647)
);

BUFx12f_ASAP7_75t_L g1648 ( 
.A(n_1558),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1612),
.A2(n_1494),
.B1(n_1428),
.B2(n_1473),
.Y(n_1649)
);

BUFx2_ASAP7_75t_SL g1650 ( 
.A(n_1549),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1528),
.Y(n_1651)
);

BUFx4f_ASAP7_75t_SL g1652 ( 
.A(n_1585),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1535),
.A2(n_1428),
.B1(n_1473),
.B2(n_1385),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1421),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1570),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1611),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1523),
.A2(n_1418),
.B1(n_451),
.B2(n_452),
.Y(n_1657)
);

CKINVDCx16_ASAP7_75t_R g1658 ( 
.A(n_1506),
.Y(n_1658)
);

BUFx10_ASAP7_75t_L g1659 ( 
.A(n_1570),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1621),
.A2(n_450),
.B1(n_453),
.B2(n_454),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1502),
.B(n_456),
.Y(n_1661)
);

CKINVDCx11_ASAP7_75t_R g1662 ( 
.A(n_1505),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1522),
.Y(n_1663)
);

BUFx12f_ASAP7_75t_L g1664 ( 
.A(n_1529),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1584),
.Y(n_1665)
);

BUFx2_ASAP7_75t_SL g1666 ( 
.A(n_1518),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1576),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1534),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1500),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1602),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1509),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1617),
.Y(n_1672)
);

INVx6_ASAP7_75t_L g1673 ( 
.A(n_1524),
.Y(n_1673)
);

BUFx4f_ASAP7_75t_SL g1674 ( 
.A(n_1572),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1566),
.Y(n_1675)
);

INVx6_ASAP7_75t_L g1676 ( 
.A(n_1507),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1617),
.Y(n_1677)
);

BUFx8_ASAP7_75t_L g1678 ( 
.A(n_1517),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1608),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1620),
.A2(n_1505),
.B1(n_1567),
.B2(n_1560),
.Y(n_1680)
);

INVx8_ASAP7_75t_L g1681 ( 
.A(n_1507),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1615),
.Y(n_1682)
);

CKINVDCx11_ASAP7_75t_R g1683 ( 
.A(n_1606),
.Y(n_1683)
);

INVx6_ASAP7_75t_L g1684 ( 
.A(n_1606),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1504),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1591),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1556),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1551),
.A2(n_1527),
.B1(n_1580),
.B2(n_1579),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1503),
.A2(n_1532),
.B(n_1553),
.Y(n_1689)
);

BUFx8_ASAP7_75t_L g1690 ( 
.A(n_1598),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1605),
.B(n_1545),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1589),
.A2(n_1607),
.B1(n_1577),
.B2(n_1616),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1626),
.A2(n_1552),
.B1(n_1575),
.B2(n_1542),
.Y(n_1693)
);

BUFx12f_ASAP7_75t_L g1694 ( 
.A(n_1604),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1537),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1569),
.A2(n_1515),
.B1(n_1561),
.B2(n_1568),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1587),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1590),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1594),
.A2(n_1554),
.B1(n_1539),
.B2(n_1601),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1544),
.Y(n_1700)
);

CKINVDCx11_ASAP7_75t_R g1701 ( 
.A(n_1583),
.Y(n_1701)
);

CKINVDCx11_ASAP7_75t_R g1702 ( 
.A(n_1571),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1578),
.Y(n_1703)
);

BUFx4f_ASAP7_75t_SL g1704 ( 
.A(n_1622),
.Y(n_1704)
);

CKINVDCx11_ASAP7_75t_R g1705 ( 
.A(n_1581),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1596),
.A2(n_1592),
.B1(n_1540),
.B2(n_1625),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1543),
.A2(n_1501),
.B(n_1521),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1511),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1637),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1639),
.B(n_1508),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1664),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1643),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1651),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1686),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1707),
.A2(n_1499),
.B(n_1624),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.B(n_1564),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1693),
.B(n_1689),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1671),
.B(n_1564),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1681),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1681),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1631),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1642),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1679),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1682),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1668),
.B(n_1565),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1703),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1685),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1649),
.B(n_1700),
.Y(n_1729)
);

INVx5_ASAP7_75t_L g1730 ( 
.A(n_1681),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1629),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1640),
.B(n_1619),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1638),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1676),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1697),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1654),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1676),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1672),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1647),
.B(n_1614),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1695),
.B(n_1692),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1670),
.Y(n_1741)
);

BUFx12f_ASAP7_75t_L g1742 ( 
.A(n_1701),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1677),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1663),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1689),
.A2(n_1623),
.B1(n_1618),
.B2(n_1557),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1708),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1645),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1653),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1709),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1732),
.B(n_1716),
.Y(n_1750)
);

BUFx4f_ASAP7_75t_SL g1751 ( 
.A(n_1742),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1727),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1712),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1741),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1736),
.B(n_1706),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1713),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1734),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1729),
.B(n_1691),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1717),
.A2(n_1696),
.B(n_1627),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1741),
.B(n_1640),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1687),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1717),
.A2(n_1696),
.B(n_1669),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1723),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1724),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1733),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1710),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1718),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1724),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1745),
.B(n_1669),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1729),
.B(n_1565),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1741),
.B(n_1633),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1728),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1715),
.A2(n_1735),
.B(n_1748),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1746),
.A2(n_1680),
.B1(n_1634),
.B2(n_1688),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1740),
.B(n_1699),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1750),
.B(n_1716),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1750),
.B(n_1768),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1750),
.B(n_1719),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1751),
.B(n_1734),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1752),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1750),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1765),
.B(n_1726),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1771),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1760),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1768),
.B(n_1719),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1773),
.B(n_1726),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1771),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1767),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1754),
.B(n_1710),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1761),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1766),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1770),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1787),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1780),
.B(n_1773),
.Y(n_1797)
);

AND4x1_ASAP7_75t_L g1798 ( 
.A(n_1782),
.B(n_1764),
.C(n_1759),
.D(n_1778),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1791),
.A2(n_1772),
.B(n_1777),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1786),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1783),
.A2(n_1772),
.B1(n_1747),
.B2(n_1775),
.C(n_1744),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1790),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1789),
.B(n_1749),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1780),
.B(n_1758),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1800),
.B(n_1789),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1784),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1803),
.Y(n_1808)
);

AND2x4_ASAP7_75t_SL g1809 ( 
.A(n_1797),
.B(n_1762),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1802),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1807),
.B(n_1784),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1809),
.B(n_1779),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1810),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1806),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1805),
.B(n_1779),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1808),
.B(n_1806),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1809),
.B(n_1781),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1805),
.B(n_1799),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1805),
.B(n_1799),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1814),
.B(n_1813),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1818),
.A2(n_1801),
.B1(n_1730),
.B2(n_1755),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1819),
.B(n_1798),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1815),
.B(n_1758),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1816),
.A2(n_1730),
.B1(n_1755),
.B2(n_1757),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1811),
.A2(n_1722),
.B1(n_1763),
.B2(n_1711),
.C(n_1731),
.Y(n_1825)
);

AO221x2_ASAP7_75t_L g1826 ( 
.A1(n_1812),
.A2(n_1742),
.B1(n_1662),
.B2(n_1722),
.C(n_1658),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1811),
.B(n_1788),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1812),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1817),
.A2(n_1705),
.B1(n_1762),
.B2(n_1774),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1818),
.B(n_1731),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1820),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1828),
.B(n_1788),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1830),
.B(n_1822),
.Y(n_1833)
);

OAI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1821),
.A2(n_1699),
.B1(n_1737),
.B2(n_1721),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1826),
.B(n_1781),
.Y(n_1835)
);

O2A1O1Ixp33_ASAP7_75t_SL g1836 ( 
.A1(n_1825),
.A2(n_1737),
.B(n_1641),
.C(n_1656),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1823),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1826),
.B(n_1711),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1833),
.A2(n_1824),
.B(n_1829),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1838),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1835),
.A2(n_1827),
.B(n_1563),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1834),
.A2(n_1831),
.B(n_1836),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1840),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1842),
.B(n_1837),
.Y(n_1844)
);

OAI32xp33_ASAP7_75t_L g1845 ( 
.A1(n_1839),
.A2(n_1832),
.A3(n_1834),
.B1(n_1721),
.B2(n_1720),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1841),
.Y(n_1846)
);

AND4x1_ASAP7_75t_L g1847 ( 
.A(n_1844),
.B(n_1630),
.C(n_1644),
.D(n_1610),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1843),
.B(n_1796),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1846),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1845),
.A2(n_1633),
.B(n_1661),
.Y(n_1850)
);

OAI322xp33_ASAP7_75t_L g1851 ( 
.A1(n_1846),
.A2(n_1763),
.A3(n_1785),
.B1(n_1739),
.B2(n_1754),
.C1(n_1743),
.C2(n_1547),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1849),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1848),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1847),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1850),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1851),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1847),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1849),
.B(n_1635),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1849),
.B(n_1690),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1849),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1849),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1855),
.A2(n_1652),
.B1(n_1650),
.B2(n_1632),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1861),
.B(n_1675),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1860),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1856),
.A2(n_1720),
.B(n_1762),
.C(n_1586),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1859),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1852),
.B(n_1648),
.Y(n_1867)
);

AO22x2_ASAP7_75t_L g1868 ( 
.A1(n_1854),
.A2(n_1857),
.B1(n_1853),
.B2(n_1858),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1857),
.B(n_1702),
.C(n_1690),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1858),
.B(n_1774),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1859),
.B(n_1678),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1868),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1868),
.B(n_1774),
.Y(n_1873)
);

OAI211xp5_ASAP7_75t_L g1874 ( 
.A1(n_1869),
.A2(n_1683),
.B(n_1667),
.C(n_1660),
.Y(n_1874)
);

AOI211x1_ASAP7_75t_SL g1875 ( 
.A1(n_1862),
.A2(n_1655),
.B(n_1559),
.C(n_1541),
.Y(n_1875)
);

NOR3xp33_ASAP7_75t_L g1876 ( 
.A(n_1867),
.B(n_1675),
.C(n_1550),
.Y(n_1876)
);

NOR3x2_ASAP7_75t_L g1877 ( 
.A(n_1863),
.B(n_1632),
.C(n_1694),
.Y(n_1877)
);

NAND4xp25_ASAP7_75t_SL g1878 ( 
.A(n_1865),
.B(n_1646),
.C(n_1628),
.D(n_1678),
.Y(n_1878)
);

NOR2x1p5_ASAP7_75t_L g1879 ( 
.A(n_1864),
.B(n_1655),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1872),
.B(n_1866),
.Y(n_1880)
);

NAND4xp25_ASAP7_75t_SL g1881 ( 
.A(n_1873),
.B(n_1870),
.C(n_1871),
.D(n_1657),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1879),
.B(n_1666),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1878),
.A2(n_1546),
.B1(n_1655),
.B2(n_1795),
.C(n_1794),
.Y(n_1883)
);

NOR2xp67_ASAP7_75t_L g1884 ( 
.A(n_1874),
.B(n_1730),
.Y(n_1884)
);

NOR2x1_ASAP7_75t_L g1885 ( 
.A(n_1877),
.B(n_1674),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1880),
.Y(n_1886)
);

NOR3xp33_ASAP7_75t_L g1887 ( 
.A(n_1885),
.B(n_1876),
.C(n_1875),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1882),
.Y(n_1888)
);

INVx5_ASAP7_75t_L g1889 ( 
.A(n_1884),
.Y(n_1889)
);

AOI32xp33_ASAP7_75t_L g1890 ( 
.A1(n_1881),
.A2(n_1732),
.A3(n_1792),
.B1(n_1738),
.B2(n_1698),
.Y(n_1890)
);

NOR3xp33_ASAP7_75t_SL g1891 ( 
.A(n_1886),
.B(n_1883),
.C(n_1636),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1889),
.B(n_1636),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1888),
.Y(n_1893)
);

AND4x1_ASAP7_75t_L g1894 ( 
.A(n_1891),
.B(n_1887),
.C(n_1890),
.D(n_1659),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1893),
.Y(n_1895)
);

AO22x2_ASAP7_75t_L g1896 ( 
.A1(n_1895),
.A2(n_1892),
.B1(n_1732),
.B2(n_1795),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1894),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1896),
.B1(n_1673),
.B2(n_1704),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1897),
.A2(n_1673),
.B1(n_1730),
.B2(n_1684),
.Y(n_1899)
);

OR3x1_ASAP7_75t_L g1900 ( 
.A(n_1897),
.B(n_1659),
.C(n_1735),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1900),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1898),
.Y(n_1902)
);

XNOR2xp5_ASAP7_75t_L g1903 ( 
.A(n_1902),
.B(n_1899),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1901),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1903),
.A2(n_1519),
.B(n_1512),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1905),
.A2(n_1904),
.B1(n_1792),
.B2(n_1684),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1905),
.A2(n_1792),
.B1(n_1776),
.B2(n_1793),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1906),
.B(n_1603),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1907),
.A2(n_1600),
.B(n_1593),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1908),
.B(n_1603),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1910),
.A2(n_1909),
.B1(n_1753),
.B2(n_1756),
.C(n_1769),
.Y(n_1911)
);

AOI211xp5_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1588),
.B(n_1582),
.C(n_1555),
.Y(n_1912)
);


endmodule