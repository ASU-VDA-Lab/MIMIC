module fake_jpeg_11163_n_432 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_9),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_50),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_57),
.Y(n_95)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_21),
.A2(n_9),
.B1(n_14),
.B2(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_36),
.B1(n_32),
.B2(n_26),
.Y(n_103)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_25),
.B(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_81),
.B(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_93),
.Y(n_141)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_8),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_43),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_57),
.Y(n_98)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_100),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_103),
.A2(n_112),
.B1(n_124),
.B2(n_31),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_106),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_37),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_51),
.A2(n_21),
.B1(n_36),
.B2(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_38),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_126),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_43),
.B1(n_22),
.B2(n_24),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_38),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_26),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_74),
.B1(n_80),
.B2(n_85),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_167),
.B1(n_187),
.B2(n_141),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_156),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_160),
.Y(n_195)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_161),
.Y(n_194)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_162),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_95),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_163),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_169),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_166),
.Y(n_227)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_177),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_100),
.A2(n_63),
.B1(n_90),
.B2(n_50),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_127),
.B1(n_79),
.B2(n_58),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_41),
.Y(n_177)
);

AOI32xp33_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_50),
.A3(n_22),
.B1(n_24),
.B2(n_88),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_183),
.Y(n_192)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_182),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_122),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_87),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_103),
.A2(n_66),
.B1(n_56),
.B2(n_59),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_117),
.A2(n_23),
.B1(n_17),
.B2(n_20),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_119),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_117),
.A2(n_23),
.B1(n_20),
.B2(n_34),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_104),
.A2(n_70),
.B1(n_54),
.B2(n_69),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_193),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_133),
.B1(n_129),
.B2(n_135),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_60),
.B1(n_67),
.B2(n_137),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_137),
.B1(n_104),
.B2(n_107),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_107),
.B1(n_114),
.B2(n_146),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_127),
.B1(n_134),
.B2(n_108),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_114),
.B1(n_183),
.B2(n_134),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_218),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_146),
.B1(n_109),
.B2(n_113),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_164),
.A2(n_180),
.B1(n_155),
.B2(n_109),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_113),
.B1(n_93),
.B2(n_41),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_182),
.B1(n_154),
.B2(n_153),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_158),
.A2(n_75),
.B1(n_131),
.B2(n_120),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_182),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_168),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_150),
.C(n_184),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_244),
.C(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_173),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_218),
.Y(n_266)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_232),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_159),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_241),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_150),
.B(n_149),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_234),
.A2(n_253),
.B(n_254),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_237),
.Y(n_264)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_197),
.B(n_37),
.Y(n_237)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g244 ( 
.A(n_192),
.B(n_152),
.C(n_148),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_246),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_249),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_206),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_175),
.B(n_162),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_219),
.B(n_216),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_252),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_199),
.A2(n_161),
.B(n_191),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_199),
.A2(n_179),
.B(n_171),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_258),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_194),
.B1(n_201),
.B2(n_212),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_215),
.A2(n_218),
.B(n_223),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_210),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_193),
.B1(n_208),
.B2(n_204),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_259),
.A2(n_238),
.B1(n_245),
.B2(n_242),
.Y(n_301)
);

AO22x1_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_198),
.B1(n_211),
.B2(n_202),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_260),
.A2(n_261),
.B(n_276),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_274),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_266),
.B(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_217),
.C(n_205),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_279),
.C(n_251),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_163),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_253),
.B(n_254),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_248),
.A2(n_225),
.B1(n_226),
.B2(n_209),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_277),
.B1(n_250),
.B2(n_249),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_226),
.B1(n_209),
.B2(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_217),
.C(n_227),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_235),
.B(n_216),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_285),
.B(n_263),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_266),
.B(n_261),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_288),
.A2(n_289),
.B(n_276),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_229),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_300),
.C(n_302),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_250),
.A3(n_228),
.B1(n_246),
.B2(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_294),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_293),
.A2(n_295),
.B1(n_309),
.B2(n_273),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_247),
.B1(n_257),
.B2(n_239),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_297),
.B(n_268),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_238),
.B1(n_239),
.B2(n_234),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_301),
.B1(n_277),
.B2(n_275),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_284),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_229),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_230),
.C(n_255),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_304),
.C(n_305),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_258),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_220),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_237),
.Y(n_306)
);

AO22x2_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_240),
.B1(n_232),
.B2(n_236),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_269),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_314),
.B(n_281),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_232),
.B1(n_194),
.B2(n_201),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_219),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_222),
.C(n_196),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_264),
.B(n_232),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_281),
.B(n_280),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_262),
.B(n_224),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_276),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_325),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_321),
.A2(n_327),
.B1(n_335),
.B2(n_323),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_323),
.A2(n_291),
.B(n_292),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_324),
.A2(n_328),
.B1(n_331),
.B2(n_334),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_274),
.Y(n_325)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_262),
.B1(n_280),
.B2(n_265),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_293),
.A2(n_295),
.B1(n_296),
.B2(n_294),
.Y(n_329)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_329),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_265),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_336),
.C(n_339),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_260),
.B1(n_268),
.B2(n_267),
.Y(n_331)
);

XOR2x2_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_337),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_313),
.A2(n_260),
.B1(n_267),
.B2(n_194),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_300),
.B(n_179),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_304),
.B(n_194),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_307),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_222),
.C(n_196),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_SL g341 ( 
.A(n_322),
.B(n_313),
.C(n_288),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_354),
.B1(n_324),
.B2(n_337),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_344),
.A2(n_348),
.B1(n_351),
.B2(n_224),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_319),
.A2(n_291),
.B1(n_311),
.B2(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_308),
.B1(n_307),
.B2(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_339),
.C(n_332),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_315),
.C(n_333),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_326),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_307),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_334),
.Y(n_357)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_360),
.B(n_330),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_369),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_332),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_366),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_325),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_373),
.C(n_358),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_375),
.B1(n_352),
.B2(n_355),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_338),
.C(n_201),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_377),
.Y(n_378)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_347),
.C(n_346),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_382),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_391),
.C(n_361),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_348),
.C(n_347),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_385),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_358),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_343),
.C(n_340),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_388),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_340),
.C(n_350),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_355),
.B1(n_356),
.B2(n_341),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_390),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_351),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_360),
.C(n_40),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_382),
.A2(n_372),
.B(n_367),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_392),
.A2(n_393),
.B(n_394),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_365),
.B(n_374),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_378),
.A2(n_373),
.B(n_368),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_24),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_385),
.A2(n_181),
.B(n_44),
.Y(n_396)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_44),
.B(n_40),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_398),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_34),
.B(n_166),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_379),
.B(n_166),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_401),
.B(n_383),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_413),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_10),
.B1(n_14),
.B2(n_2),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_407),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_24),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_409),
.B(n_413),
.Y(n_418)
);

A2O1A1O1Ixp25_ASAP7_75t_L g411 ( 
.A1(n_403),
.A2(n_8),
.B(n_15),
.C(n_2),
.D(n_3),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_412),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_0),
.C(n_1),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_22),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_403),
.C(n_22),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_415),
.B(n_417),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_22),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_8),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_10),
.C(n_12),
.Y(n_424)
);

OAI321xp33_ASAP7_75t_L g422 ( 
.A1(n_417),
.A2(n_408),
.A3(n_411),
.B1(n_3),
.B2(n_6),
.C(n_7),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_422),
.A2(n_423),
.B(n_7),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_419),
.B(n_416),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_7),
.C(n_11),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_421),
.A2(n_6),
.B(n_7),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_425),
.B(n_426),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_428),
.A2(n_427),
.B(n_12),
.Y(n_429)
);

OAI321xp33_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_0),
.A3(n_1),
.B1(n_12),
.B2(n_13),
.C(n_419),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_430),
.A2(n_13),
.B(n_0),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_1),
.Y(n_432)
);


endmodule