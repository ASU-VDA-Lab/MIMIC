module fake_jpeg_7633_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_17),
.B1(n_26),
.B2(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_52),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_67),
.B1(n_70),
.B2(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_29),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_54),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_22),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_48),
.B1(n_22),
.B2(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_70)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_80),
.B1(n_68),
.B2(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_75),
.Y(n_111)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_48),
.B1(n_37),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_68),
.B1(n_57),
.B2(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_84),
.B(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_99),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_49),
.B(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_53),
.B(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_53),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_103),
.B1(n_25),
.B2(n_30),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_66),
.C(n_61),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_118),
.C(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_54),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_105),
.B1(n_127),
.B2(n_96),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_116),
.B1(n_85),
.B2(n_25),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_54),
.B1(n_69),
.B2(n_37),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_54),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_99),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_60),
.A3(n_38),
.B1(n_42),
.B2(n_47),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_38),
.C(n_55),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_134),
.B1(n_138),
.B2(n_126),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_133),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_122),
.B(n_27),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_88),
.B1(n_93),
.B2(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_99),
.B1(n_74),
.B2(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_78),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_95),
.B(n_21),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_149),
.B(n_155),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_73),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_153),
.B1(n_157),
.B2(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_38),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_154),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_82),
.B1(n_90),
.B2(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_27),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_42),
.C(n_65),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_65),
.C(n_36),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_104),
.A2(n_75),
.B1(n_27),
.B2(n_30),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_171),
.C(n_187),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_164),
.B(n_167),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_151),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_163),
.B(n_166),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_23),
.B(n_110),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_23),
.B(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_168),
.B(n_172),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_38),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_119),
.B1(n_117),
.B2(n_126),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_189),
.B1(n_148),
.B2(n_177),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_32),
.B(n_34),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_185),
.B(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_180),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_182),
.B1(n_130),
.B2(n_136),
.Y(n_197)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_179),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_33),
.A3(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_117),
.B1(n_101),
.B2(n_65),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_140),
.B1(n_157),
.B2(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_176),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_36),
.B(n_34),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_21),
.B(n_47),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_200),
.B1(n_203),
.B2(n_210),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_149),
.B1(n_135),
.B2(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_156),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_165),
.C(n_170),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_208),
.B1(n_211),
.B2(n_177),
.Y(n_240)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_148),
.B1(n_155),
.B2(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_133),
.B1(n_131),
.B2(n_154),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_184),
.B1(n_181),
.B2(n_170),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_13),
.C(n_16),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_15),
.C(n_14),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_218),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_165),
.B(n_133),
.CI(n_131),
.CON(n_218),
.SN(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_168),
.B1(n_163),
.B2(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_220),
.B1(n_21),
.B2(n_47),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_133),
.B1(n_33),
.B2(n_36),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_191),
.B(n_189),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_223),
.Y(n_260)
);

BUFx4f_ASAP7_75t_SL g224 ( 
.A(n_194),
.Y(n_224)
);

INVx11_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_162),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_228),
.C(n_230),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_226),
.A2(n_238),
.B1(n_243),
.B2(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_235),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_187),
.C(n_185),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_175),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_167),
.C(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_164),
.C(n_161),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_179),
.B1(n_177),
.B2(n_36),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_244),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_205),
.B1(n_206),
.B2(n_215),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_47),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_34),
.B1(n_32),
.B2(n_21),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_198),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_195),
.A2(n_34),
.B1(n_21),
.B2(n_2),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_204),
.B1(n_201),
.B2(n_195),
.Y(n_266)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_222),
.B(n_236),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_266),
.B1(n_267),
.B2(n_225),
.Y(n_279)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_264),
.B1(n_265),
.B2(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_199),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_212),
.B1(n_218),
.B2(n_197),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_220),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_232),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_227),
.C(n_230),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_282),
.C(n_287),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_245),
.B(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_246),
.B1(n_198),
.B2(n_241),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_286),
.B1(n_266),
.B2(n_267),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_228),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_13),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_257),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_21),
.C(n_1),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_257),
.B(n_13),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_251),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_0),
.C(n_1),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_256),
.B(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_301),
.B1(n_6),
.B2(n_7),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_297),
.B1(n_288),
.B2(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_254),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_293),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_255),
.C(n_253),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_299),
.C(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_259),
.B1(n_262),
.B2(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_252),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_274),
.B(n_5),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_255),
.C(n_254),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_260),
.B1(n_4),
.B2(n_5),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_309),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_283),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_287),
.C(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_310),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_5),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_301),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_8),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_315),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_8),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_314),
.B(n_295),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_8),
.C(n_9),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_321),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_289),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_324),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_290),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_303),
.B(n_309),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_306),
.B(n_313),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_331),
.B(n_9),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_317),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_305),
.B(n_10),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_330),
.B(n_332),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_9),
.B(n_10),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_323),
.A2(n_317),
.B(n_324),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_327),
.Y(n_337)
);

AO21x2_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_326),
.B(n_11),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_12),
.B(n_10),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_11),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_12),
.Y(n_341)
);


endmodule