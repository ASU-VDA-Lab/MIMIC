module fake_jpeg_3518_n_276 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_10),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_53),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_59),
.Y(n_86)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_36),
.Y(n_84)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_70),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_29),
.B1(n_25),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_75),
.B1(n_21),
.B2(n_27),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_74),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_34),
.B1(n_30),
.B2(n_21),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_18),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_78),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_30),
.C(n_34),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_29),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_52),
.Y(n_114)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_39),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_42),
.A2(n_38),
.B(n_23),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_107),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_45),
.B1(n_62),
.B2(n_50),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_122),
.B1(n_90),
.B2(n_103),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_136),
.Y(n_150)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_127),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_75),
.B1(n_78),
.B2(n_54),
.Y(n_122)
);

OR2x2_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_52),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_114),
.Y(n_147)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_27),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_77),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

BUFx4f_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_76),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_153),
.C(n_154),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_136),
.B1(n_124),
.B2(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_143),
.B(n_157),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_77),
.B(n_98),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_80),
.B(n_133),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_80),
.B(n_81),
.C(n_52),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_136),
.B(n_19),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_152),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_163),
.B(n_105),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_161),
.C(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_54),
.B1(n_82),
.B2(n_25),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_82),
.C(n_33),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_33),
.C(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_13),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_13),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_89),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_126),
.C(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_126),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_179),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_132),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_183),
.C(n_187),
.Y(n_208)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_184),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_181),
.B(n_190),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_188),
.B1(n_163),
.B2(n_137),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_131),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_125),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_162),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_89),
.B(n_115),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_147),
.C(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_113),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_111),
.C(n_38),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_137),
.A2(n_38),
.B(n_1),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_144),
.B(n_152),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_201),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_203),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_178),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_206),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_183),
.B1(n_167),
.B2(n_187),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_154),
.A3(n_12),
.B1(n_14),
.B2(n_16),
.C1(n_4),
.C2(n_3),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_139),
.B(n_159),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_168),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_221),
.C(n_202),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_176),
.B(n_173),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_222),
.B(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_167),
.B1(n_185),
.B2(n_190),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_214),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_12),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_170),
.C(n_151),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_182),
.B(n_170),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_209),
.B(n_192),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_163),
.B(n_164),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_226),
.B(n_195),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_193),
.B(n_204),
.C(n_209),
.D(n_191),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_197),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_212),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_231),
.C(n_237),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_220),
.B(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_196),
.C(n_200),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_235),
.C(n_195),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_239),
.B1(n_241),
.B2(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_196),
.C(n_207),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_213),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_224),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_194),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_230),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_250),
.C(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_3),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_174),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_247),
.B(n_194),
.Y(n_259)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_0),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_263),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_0),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_255),
.C(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_256),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_253),
.C(n_267),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_272),
.B(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_273),
.Y(n_276)
);


endmodule