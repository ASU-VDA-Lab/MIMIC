module fake_netlist_1_3750_n_552 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_552);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_552;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g78 ( .A(n_14), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_72), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_62), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_30), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_64), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_21), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_61), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_20), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_57), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_11), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_31), .Y(n_90) );
NOR2xp67_ASAP7_75t_L g91 ( .A(n_3), .B(n_40), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_48), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_42), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_5), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_8), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_74), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_13), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_43), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_1), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_65), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_70), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_24), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_27), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_46), .B(n_51), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_56), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_16), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_0), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_45), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_93), .B(n_0), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_96), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_113), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_92), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_103), .B(n_2), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_105), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_96), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_92), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_105), .B(n_87), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_112), .B(n_2), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_112), .B(n_3), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_82), .B(n_4), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_79), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_110), .B(n_4), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_80), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_118), .B(n_94), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_117), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_129), .B(n_99), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_118), .B(n_97), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_130), .A2(n_100), .B1(n_78), .B2(n_95), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_116), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
BUFx10_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_122), .B(n_102), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_116), .B(n_85), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_123), .B(n_111), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_122), .A2(n_106), .B1(n_81), .B2(n_102), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_136), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_121), .B(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_115), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_121), .B(n_101), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_115), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_137), .B(n_101), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_129), .B(n_88), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_148), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_164), .A2(n_114), .B1(n_135), .B2(n_119), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_164), .B(n_119), .Y(n_168) );
BUFx4f_ASAP7_75t_SL g169 ( .A(n_145), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_164), .B(n_114), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_160), .B(n_132), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g175 ( .A(n_140), .B(n_128), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_148), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_160), .B(n_132), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_151), .B(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_151), .B(n_88), .Y(n_181) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_160), .B(n_127), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_156), .B(n_126), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_154), .A2(n_124), .B1(n_81), .B2(n_120), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
CKINVDCx14_ASAP7_75t_R g189 ( .A(n_156), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
AOI22xp5_ASAP7_75t_SL g191 ( .A1(n_144), .A2(n_98), .B1(n_90), .B2(n_104), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_154), .A2(n_120), .B1(n_104), .B2(n_108), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_156), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_161), .A2(n_120), .B1(n_108), .B2(n_90), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_141), .B(n_120), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_196), .B(n_158), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_172), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_178), .A2(n_143), .B(n_139), .C(n_141), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_178), .A2(n_139), .B(n_143), .C(n_152), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_180), .Y(n_207) );
INVxp67_ASAP7_75t_SL g208 ( .A(n_165), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_170), .Y(n_210) );
AOI21xp33_ASAP7_75t_L g211 ( .A1(n_181), .A2(n_158), .B(n_152), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_186), .B(n_158), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_167), .A2(n_161), .B1(n_152), .B2(n_150), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_196), .A2(n_144), .B1(n_152), .B2(n_150), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_168), .A2(n_152), .B(n_153), .C(n_155), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_180), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_169), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_186), .B(n_155), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_168), .A2(n_91), .B(n_107), .C(n_159), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_171), .B(n_109), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_174), .A2(n_159), .B(n_157), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_174), .A2(n_157), .B(n_142), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_171), .A2(n_146), .B1(n_125), .B2(n_115), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_184), .B(n_5), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_188), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_183), .A2(n_142), .B(n_147), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_187), .A2(n_125), .B1(n_146), .B2(n_131), .C(n_134), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_188), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_200), .A2(n_189), .B1(n_171), .B2(n_187), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_218), .Y(n_235) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_229), .A2(n_179), .B(n_185), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_222), .A2(n_171), .B1(n_194), .B2(n_177), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_219), .B(n_206), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_206), .B(n_190), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_202), .B(n_190), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_224), .A2(n_179), .B(n_185), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_230), .A2(n_198), .B(n_195), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_222), .A2(n_194), .B1(n_188), .B2(n_173), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_202), .Y(n_245) );
AND2x4_ASAP7_75t_SL g246 ( .A(n_202), .B(n_221), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_202), .B(n_166), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_221), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_199), .A2(n_191), .B1(n_173), .B2(n_183), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_227), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_221), .B(n_182), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_221), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_222), .A2(n_167), .B1(n_182), .B2(n_175), .Y(n_253) );
NOR2xp67_ASAP7_75t_L g254 ( .A(n_209), .B(n_192), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_232), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_209), .B(n_182), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_212), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_205), .B(n_191), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g260 ( .A1(n_249), .A2(n_201), .B1(n_211), .B2(n_215), .C(n_205), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_249), .A2(n_201), .B1(n_213), .B2(n_220), .C(n_226), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
OAI21x1_ASAP7_75t_SL g264 ( .A1(n_248), .A2(n_195), .B(n_223), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_233), .B(n_198), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_244), .A2(n_216), .B1(n_208), .B2(n_232), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_258), .A2(n_182), .B1(n_209), .B2(n_210), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_259), .A2(n_228), .B1(n_175), .B2(n_231), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_236), .A2(n_216), .B(n_220), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_237), .A2(n_197), .B1(n_228), .B2(n_225), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_236), .A2(n_217), .B(n_207), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_259), .A2(n_193), .B1(n_192), .B2(n_204), .C(n_228), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_241), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_241), .A2(n_214), .B(n_210), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_238), .A2(n_193), .B1(n_192), .B2(n_214), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_235), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_242), .A2(n_214), .B(n_210), .C(n_193), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g278 ( .A1(n_253), .A2(n_193), .B1(n_192), .B2(n_176), .C(n_166), .Y(n_278) );
AOI22xp5_ASAP7_75t_SL g279 ( .A1(n_238), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_242), .A2(n_125), .B(n_142), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_242), .A2(n_147), .B(n_134), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_281), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_262), .B(n_238), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_279), .B(n_238), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_273), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_265), .B(n_243), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_273), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_282), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_282), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_277), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_282), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_269), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_280), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_266), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_271), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_274), .Y(n_302) );
NOR2xp67_ASAP7_75t_SL g303 ( .A(n_260), .B(n_248), .Y(n_303) );
NOR2xp33_ASAP7_75t_R g304 ( .A(n_276), .B(n_245), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_261), .B(n_255), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_295), .A2(n_267), .B(n_270), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_289), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_294), .Y(n_308) );
AOI211xp5_ASAP7_75t_L g309 ( .A1(n_286), .A2(n_304), .B(n_303), .C(n_305), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_286), .A2(n_268), .B1(n_272), .B2(n_275), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_288), .B(n_268), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_294), .Y(n_313) );
OAI33xp33_ASAP7_75t_L g314 ( .A1(n_283), .A2(n_6), .A3(n_7), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_298), .B(n_243), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_298), .B(n_243), .Y(n_316) );
CKINVDCx9p33_ASAP7_75t_R g317 ( .A(n_293), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_297), .A2(n_275), .B1(n_239), .B2(n_256), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_295), .B(n_250), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_294), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_297), .A2(n_239), .B1(n_256), .B2(n_250), .Y(n_321) );
NAND2x1_ASAP7_75t_SL g322 ( .A(n_292), .B(n_248), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g323 ( .A1(n_303), .A2(n_245), .B(n_252), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_302), .A2(n_252), .B(n_254), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_290), .B(n_248), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_293), .B(n_250), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_292), .B(n_252), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_287), .B(n_131), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_284), .A2(n_239), .B1(n_240), .B2(n_278), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_291), .B(n_240), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_291), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_288), .B(n_134), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_328), .B(n_301), .Y(n_337) );
NAND4xp25_ASAP7_75t_L g338 ( .A(n_309), .B(n_311), .C(n_318), .D(n_332), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_336), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_324), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_324), .B(n_285), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_313), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_328), .B(n_301), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_312), .B(n_285), .Y(n_344) );
AND2x4_ASAP7_75t_SL g345 ( .A(n_313), .B(n_284), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_334), .B(n_302), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_334), .B(n_300), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_328), .B(n_300), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_336), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_312), .B(n_299), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_336), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_310), .B(n_296), .Y(n_352) );
OAI31xp33_ASAP7_75t_L g353 ( .A1(n_311), .A2(n_257), .A3(n_251), .B(n_246), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_310), .B(n_299), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_310), .B(n_134), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_309), .B(n_246), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_307), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_330), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_335), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_330), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_319), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_330), .B(n_134), .Y(n_365) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_318), .B(n_254), .C(n_239), .D(n_240), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_319), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_308), .B(n_320), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_330), .B(n_134), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_308), .B(n_9), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_330), .B(n_10), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_331), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_314), .B(n_12), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_315), .B(n_13), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_315), .B(n_14), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_322), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_316), .B(n_246), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_308), .B(n_133), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_344), .B(n_316), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_364), .B(n_367), .Y(n_383) );
OR2x2_ASAP7_75t_SL g384 ( .A(n_371), .B(n_317), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_364), .B(n_316), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_379), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_367), .B(n_320), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_359), .B(n_320), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_368), .B(n_335), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_345), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_368), .B(n_306), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_337), .B(n_325), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_340), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_342), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_341), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_337), .B(n_343), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_339), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_343), .B(n_325), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_376), .B(n_306), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_SL g406 ( .A1(n_356), .A2(n_326), .B(n_317), .C(n_323), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_339), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_348), .B(n_325), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_369), .Y(n_410) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_379), .B(n_329), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_345), .Y(n_412) );
NOR2x1p5_ASAP7_75t_L g413 ( .A(n_338), .B(n_314), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_376), .B(n_306), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_348), .B(n_325), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_350), .B(n_347), .Y(n_416) );
NAND4xp25_ASAP7_75t_L g417 ( .A(n_353), .B(n_375), .C(n_366), .D(n_378), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_354), .B(n_306), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_354), .B(n_329), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_372), .A2(n_332), .B1(n_321), .B2(n_329), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_347), .B(n_333), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_373), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_346), .B(n_333), .Y(n_423) );
AND4x1_ASAP7_75t_L g424 ( .A(n_373), .B(n_321), .C(n_331), .D(n_322), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_346), .B(n_333), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_352), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_358), .B(n_329), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_363), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_371), .A2(n_329), .B(n_326), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_349), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_358), .B(n_333), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_361), .B(n_331), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_361), .B(n_323), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_388), .B(n_352), .Y(n_435) );
OAI221xp5_ASAP7_75t_SL g436 ( .A1(n_424), .A2(n_377), .B1(n_380), .B2(n_381), .C(n_374), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_416), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_400), .B(n_374), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_413), .A2(n_370), .B1(n_365), .B2(n_355), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_400), .B(n_351), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_417), .A2(n_351), .B1(n_349), .B2(n_365), .C(n_370), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_384), .A2(n_381), .B1(n_355), .B2(n_247), .Y(n_445) );
AO21x1_ASAP7_75t_L g446 ( .A1(n_411), .A2(n_251), .B(n_257), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_133), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_398), .B(n_399), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_385), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_406), .A2(n_251), .B(n_257), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_387), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_426), .Y(n_452) );
OAI221xp5_ASAP7_75t_SL g453 ( .A1(n_420), .A2(n_247), .B1(n_147), .B2(n_240), .C(n_22), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_406), .A2(n_247), .B(n_133), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_388), .B(n_393), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_418), .B(n_133), .Y(n_458) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_401), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_388), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_420), .A2(n_247), .B1(n_133), .B2(n_162), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_383), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_412), .A2(n_247), .B1(n_176), .B2(n_162), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_429), .A2(n_17), .B(n_18), .C(n_19), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_403), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_410), .B(n_23), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_408), .B(n_25), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_395), .A2(n_162), .B1(n_163), .B2(n_29), .C(n_32), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_418), .B(n_26), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_401), .Y(n_470) );
OAI21xp33_ASAP7_75t_SL g471 ( .A1(n_395), .A2(n_28), .B(n_34), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_402), .B(n_35), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_419), .B(n_36), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_407), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_389), .A2(n_162), .B1(n_163), .B2(n_39), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_389), .A2(n_37), .B(n_38), .C(n_41), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_421), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_404), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_389), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
XNOR2x1_ASAP7_75t_L g482 ( .A(n_445), .B(n_391), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_443), .A2(n_402), .B1(n_422), .B2(n_409), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_462), .B(n_415), .Y(n_484) );
XNOR2x1_ASAP7_75t_L g485 ( .A(n_457), .B(n_423), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_479), .B(n_415), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_448), .A2(n_409), .B1(n_382), .B2(n_427), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_473), .Y(n_489) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_436), .B(n_425), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_471), .A2(n_394), .B(n_405), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_448), .B(n_414), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_436), .A2(n_423), .B1(n_425), .B2(n_392), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_451), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_442), .B(n_386), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_452), .B(n_432), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_455), .B(n_428), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_474), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_456), .B(n_430), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_465), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_478), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_440), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_452), .B(n_434), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_444), .B(n_434), .Y(n_505) );
OAI31xp33_ASAP7_75t_SL g506 ( .A1(n_467), .A2(n_427), .A3(n_431), .B(n_433), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g507 ( .A1(n_441), .A2(n_431), .B(n_433), .Y(n_507) );
XOR2x2_ASAP7_75t_L g508 ( .A(n_435), .B(n_44), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_446), .B(n_430), .Y(n_509) );
AOI221x1_ASAP7_75t_L g510 ( .A1(n_494), .A2(n_458), .B1(n_464), .B2(n_454), .C(n_466), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_494), .A2(n_477), .B1(n_447), .B2(n_461), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_484), .B(n_459), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_507), .A2(n_453), .B1(n_461), .B2(n_459), .C(n_470), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_480), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_506), .A2(n_453), .B1(n_450), .B2(n_460), .C(n_472), .Y(n_515) );
AOI21xp33_ASAP7_75t_SL g516 ( .A1(n_485), .A2(n_460), .B(n_476), .Y(n_516) );
AOI32xp33_ASAP7_75t_L g517 ( .A1(n_482), .A2(n_470), .A3(n_463), .B1(n_468), .B2(n_469), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_491), .B(n_407), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_497), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_506), .A2(n_475), .B1(n_162), .B2(n_163), .C(n_53), .Y(n_520) );
AOI211xp5_ASAP7_75t_L g521 ( .A1(n_509), .A2(n_162), .B(n_50), .C(n_52), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g522 ( .A1(n_483), .A2(n_47), .B1(n_54), .B2(n_55), .C1(n_58), .C2(n_59), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_498), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_498), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_489), .B(n_493), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_490), .A2(n_162), .B1(n_163), .B2(n_66), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_504), .B(n_60), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g528 ( .A1(n_517), .A2(n_488), .B1(n_492), .B2(n_487), .C(n_481), .Y(n_528) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_522), .B(n_502), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_525), .A2(n_486), .B1(n_505), .B2(n_495), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_516), .A2(n_503), .B(n_496), .C(n_501), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g532 ( .A1(n_510), .A2(n_508), .B(n_500), .C(n_499), .Y(n_532) );
NOR4xp25_ASAP7_75t_L g533 ( .A(n_514), .B(n_500), .C(n_163), .D(n_69), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_519), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_523), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_524), .A2(n_63), .B1(n_67), .B2(n_71), .C(n_73), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_520), .A2(n_75), .B(n_76), .C(n_77), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_534), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_531), .A2(n_511), .B1(n_515), .B2(n_526), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_532), .A2(n_513), .B1(n_521), .B2(n_512), .C(n_527), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_530), .B(n_518), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_535), .Y(n_542) );
NOR4xp25_ASAP7_75t_L g543 ( .A(n_539), .B(n_528), .C(n_537), .D(n_536), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_538), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_541), .B(n_529), .Y(n_545) );
OA22x2_ASAP7_75t_L g546 ( .A1(n_545), .A2(n_539), .B1(n_542), .B2(n_540), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_545), .B(n_533), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_546), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_548), .Y(n_549) );
AO22x2_ASAP7_75t_L g550 ( .A1(n_549), .A2(n_544), .B1(n_547), .B2(n_543), .Y(n_550) );
OR2x6_ASAP7_75t_L g551 ( .A(n_550), .B(n_518), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_551), .A2(n_146), .B1(n_546), .B2(n_545), .Y(n_552) );
endmodule