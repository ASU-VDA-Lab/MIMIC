module fake_jpeg_16469_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx24_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_1),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_4),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_5),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_55),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_19),
.A2(n_13),
.B1(n_8),
.B2(n_9),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_32),
.B(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_10),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_58),
.B(n_22),
.C(n_32),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_19),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_36),
.B(n_14),
.Y(n_89)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_6),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_15),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_30),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_18),
.B1(n_31),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_18),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_61),
.B1(n_72),
.B2(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_15),
.C(n_14),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_14),
.C(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_9),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_77),
.B1(n_66),
.B2(n_76),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_114),
.B1(n_90),
.B2(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_46),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_102),
.C(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_50),
.B1(n_52),
.B2(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_66),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_84),
.C(n_73),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_14),
.B1(n_17),
.B2(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_60),
.B(n_17),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_81),
.B1(n_82),
.B2(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_119),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_67),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_88),
.B1(n_67),
.B2(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_60),
.B(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_71),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_71),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_64),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_131),
.B(n_102),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_113),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_87),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_90),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_107),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_107),
.B1(n_104),
.B2(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_97),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_98),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_93),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_151),
.C(n_160),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_154),
.Y(n_166)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_96),
.C(n_100),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_99),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_161),
.C(n_123),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_159),
.B1(n_139),
.B2(n_141),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_129),
.B1(n_136),
.B2(n_131),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_115),
.C(n_132),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_115),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_122),
.B1(n_128),
.B2(n_123),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_149),
.B1(n_162),
.B2(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_168),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_120),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_173),
.C(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_125),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_148),
.B(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_125),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_176),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_160),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_181),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_173),
.B(n_165),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_126),
.B1(n_133),
.B2(n_121),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_126),
.B(n_121),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_151),
.B1(n_149),
.B2(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_176),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_191),
.B1(n_182),
.B2(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_184),
.C(n_180),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_180),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_182),
.B(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_178),
.B1(n_177),
.B2(n_181),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_183),
.B1(n_191),
.B2(n_196),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_198),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_197),
.B(n_201),
.C(n_200),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule