module fake_jpeg_14332_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_68),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_69),
.Y(n_209)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_76),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_77),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_89),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_93),
.Y(n_212)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_98),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_38),
.B(n_9),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_111),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_102),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_105),
.Y(n_201)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_110),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_6),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_113),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

BUFx4f_ASAP7_75t_L g116 ( 
.A(n_20),
.Y(n_116)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_6),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_129),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

BUFx4f_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

CKINVDCx6p67_ASAP7_75t_R g203 ( 
.A(n_126),
.Y(n_203)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_25),
.B(n_18),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_74),
.A2(n_59),
.B1(n_51),
.B2(n_43),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_134),
.A2(n_153),
.B1(n_161),
.B2(n_162),
.Y(n_220)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_85),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_135),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_100),
.B(n_42),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_143),
.B(n_183),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_46),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_145),
.B(n_158),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_71),
.A2(n_55),
.B1(n_46),
.B2(n_43),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_25),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_78),
.B1(n_60),
.B2(n_114),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_62),
.A2(n_59),
.B1(n_51),
.B2(n_27),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_58),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_166),
.B(n_176),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_126),
.B(n_46),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_32),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_32),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_179),
.B(n_191),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g233 ( 
.A(n_180),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_64),
.A2(n_59),
.B1(n_51),
.B2(n_58),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_181),
.A2(n_194),
.B1(n_20),
.B2(n_53),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_92),
.B(n_42),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_182),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_92),
.B(n_12),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_66),
.B(n_48),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_103),
.B(n_36),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_68),
.A2(n_56),
.B1(n_50),
.B2(n_21),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_73),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_199),
.B1(n_153),
.B2(n_161),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_79),
.A2(n_21),
.B1(n_33),
.B2(n_22),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_69),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_27),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_218),
.B(n_227),
.Y(n_330)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_219),
.Y(n_314)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_143),
.A2(n_50),
.B1(n_56),
.B2(n_124),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_221),
.B(n_242),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_131),
.A2(n_33),
.B(n_22),
.C(n_50),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_223),
.A2(n_253),
.B(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_225),
.A2(n_235),
.B1(n_260),
.B2(n_261),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_159),
.A2(n_136),
.B1(n_146),
.B2(n_131),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_226),
.A2(n_230),
.B1(n_256),
.B2(n_270),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_180),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_108),
.B1(n_107),
.B2(n_99),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_98),
.B1(n_93),
.B2(n_89),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_232),
.B(n_277),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_84),
.B1(n_83),
.B2(n_81),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_236),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_237),
.B(n_289),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_182),
.A2(n_77),
.B1(n_36),
.B2(n_29),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_SL g344 ( 
.A(n_238),
.B(n_249),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_239),
.Y(n_323)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_141),
.Y(n_241)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_159),
.B(n_28),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_243),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g245 ( 
.A1(n_135),
.A2(n_56),
.B1(n_20),
.B2(n_2),
.Y(n_245)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_130),
.Y(n_246)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_142),
.Y(n_247)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_133),
.Y(n_248)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_147),
.A2(n_28),
.B1(n_49),
.B2(n_53),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_136),
.B(n_0),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_264),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_145),
.B(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_146),
.A2(n_53),
.B1(n_49),
.B2(n_10),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_160),
.A2(n_49),
.B1(n_53),
.B2(n_10),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_169),
.A2(n_53),
.B1(n_49),
.B2(n_12),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_193),
.A2(n_49),
.B1(n_6),
.B2(n_13),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_150),
.Y(n_263)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_0),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

NAND2x1_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_1),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_283),
.C(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_1),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_177),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_199),
.A2(n_5),
.B1(n_17),
.B2(n_16),
.Y(n_270)
);

HAxp5_ASAP7_75t_SL g271 ( 
.A(n_165),
.B(n_5),
.CON(n_271),
.SN(n_271)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_271),
.Y(n_335)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_132),
.Y(n_273)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_149),
.A2(n_17),
.B1(n_18),
.B2(n_3),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_278),
.B1(n_280),
.B2(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_186),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_139),
.A2(n_17),
.B1(n_18),
.B2(n_4),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_170),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_281),
.B(n_284),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_156),
.A2(n_17),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

AOI32xp33_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_283),
.A3(n_271),
.B1(n_264),
.B2(n_288),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_201),
.A2(n_2),
.B(n_3),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_170),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_202),
.A2(n_2),
.B1(n_4),
.B2(n_175),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_210),
.B1(n_209),
.B2(n_173),
.Y(n_311)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_139),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_287),
.B(n_288),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_165),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_172),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_212),
.A2(n_4),
.B1(n_216),
.B2(n_206),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_212),
.A2(n_4),
.B1(n_216),
.B2(n_206),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_291),
.A2(n_292),
.B1(n_173),
.B2(n_171),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_214),
.A2(n_175),
.B1(n_209),
.B2(n_210),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_144),
.B(n_137),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_311),
.A2(n_287),
.B1(n_257),
.B2(n_276),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_224),
.A2(n_220),
.B1(n_255),
.B2(n_278),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_312),
.A2(n_353),
.B1(n_315),
.B2(n_300),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_279),
.B(n_190),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_327),
.C(n_328),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_318),
.B(n_342),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_204),
.C(n_165),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_338),
.C(n_240),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_293),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_322),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_222),
.B(n_198),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_333),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_242),
.B(n_189),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_229),
.B(n_140),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_222),
.B(n_168),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_240),
.B(n_204),
.C(n_203),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_293),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_339),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_237),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_343),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_252),
.B(n_151),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_267),
.B(n_168),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_254),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_346),
.B(n_259),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_285),
.B(n_187),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_233),
.B1(n_239),
.B2(n_277),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_354),
.B(n_347),
.Y(n_428)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_231),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_335),
.A2(n_262),
.B1(n_253),
.B2(n_230),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_360),
.A2(n_368),
.B(n_372),
.Y(n_426)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_221),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_364),
.B(n_369),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_301),
.A2(n_231),
.B1(n_223),
.B2(n_221),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_365),
.A2(n_366),
.B1(n_370),
.B2(n_373),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_301),
.A2(n_231),
.B1(n_253),
.B2(n_266),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_295),
.A2(n_266),
.B(n_234),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_331),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_303),
.A2(n_294),
.B1(n_298),
.B2(n_296),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_325),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_371),
.A2(n_387),
.B1(n_233),
.B2(n_244),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_297),
.B(n_324),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_303),
.A2(n_248),
.B1(n_251),
.B2(n_243),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_388),
.B1(n_398),
.B2(n_399),
.Y(n_409)
);

BUFx8_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

BUFx24_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_378),
.B(n_386),
.Y(n_418)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_332),
.Y(n_380)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_SL g382 ( 
.A1(n_344),
.A2(n_245),
.B(n_249),
.C(n_238),
.Y(n_382)
);

OA22x2_ASAP7_75t_L g408 ( 
.A1(n_382),
.A2(n_394),
.B1(n_315),
.B2(n_352),
.Y(n_408)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_297),
.A2(n_282),
.B(n_245),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_384),
.A2(n_385),
.B(n_336),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_320),
.A2(n_258),
.B(n_284),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_345),
.Y(n_386)
);

BUFx24_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_294),
.A2(n_291),
.B1(n_290),
.B2(n_274),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_228),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_351),
.Y(n_432)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_353),
.A2(n_265),
.B1(n_272),
.B2(n_236),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_346),
.B1(n_336),
.B2(n_329),
.Y(n_414)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_326),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_300),
.A2(n_280),
.B1(n_152),
.B2(n_192),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_338),
.C(n_305),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_405),
.C(n_407),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_402),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_R g403 ( 
.A(n_356),
.B(n_299),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_403),
.B(n_413),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_340),
.C(n_318),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_339),
.C(n_343),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_408),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_308),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_414),
.A2(n_429),
.B1(n_388),
.B2(n_357),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_374),
.A2(n_344),
.B1(n_305),
.B2(n_307),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_435),
.B(n_382),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_427),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_398),
.A2(n_309),
.B1(n_302),
.B2(n_308),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_421),
.A2(n_363),
.B1(n_380),
.B2(n_392),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_379),
.C(n_397),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_423),
.C(n_428),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_304),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_369),
.B(n_302),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_357),
.Y(n_448)
);

OAI32xp33_ASAP7_75t_L g427 ( 
.A1(n_397),
.A2(n_326),
.A3(n_304),
.B1(n_348),
.B2(n_347),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_366),
.A2(n_350),
.B1(n_307),
.B2(n_337),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_385),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_433),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_381),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_362),
.A2(n_306),
.B(n_316),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_348),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_427),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_442),
.B1(n_449),
.B2(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_409),
.A2(n_362),
.B1(n_365),
.B2(n_393),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_440),
.A2(n_467),
.B1(n_408),
.B2(n_436),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_437),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_457),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_358),
.B1(n_384),
.B2(n_368),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_443),
.B(n_446),
.Y(n_497)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_370),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_446),
.B(n_471),
.C(n_419),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_448),
.B(n_450),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_429),
.A2(n_404),
.B1(n_358),
.B2(n_414),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_386),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_454),
.Y(n_487)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_404),
.A2(n_360),
.B(n_373),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_455),
.A2(n_435),
.B(n_430),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_376),
.Y(n_456)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_433),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_417),
.A2(n_382),
.B1(n_389),
.B2(n_355),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_461),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_359),
.Y(n_463)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_464),
.A2(n_469),
.B1(n_410),
.B2(n_395),
.Y(n_503)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_412),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_468),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_409),
.A2(n_375),
.B1(n_396),
.B2(n_391),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_410),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_438),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_434),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_400),
.B(n_334),
.C(n_306),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_417),
.A2(n_383),
.B1(n_350),
.B2(n_337),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_472),
.A2(n_431),
.B1(n_438),
.B2(n_410),
.Y(n_500)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_415),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_416),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_423),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_475),
.A2(n_498),
.B1(n_463),
.B2(n_455),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_426),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_478),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_405),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_451),
.Y(n_486)
);

INVx11_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_426),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_494),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_490),
.A2(n_501),
.B(n_449),
.Y(n_520)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_495),
.C(n_467),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_407),
.Y(n_493)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_447),
.B(n_418),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_416),
.C(n_436),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_466),
.A2(n_421),
.B1(n_408),
.B2(n_434),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_500),
.B1(n_440),
.B2(n_464),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_505),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_443),
.B(n_408),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_502),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_455),
.A2(n_410),
.B(n_431),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_461),
.B(n_351),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_468),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_411),
.B1(n_383),
.B2(n_371),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_504),
.A2(n_452),
.B1(n_439),
.B2(n_472),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_442),
.B(n_445),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_451),
.Y(n_506)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_506),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_476),
.A2(n_459),
.B(n_481),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_511),
.A2(n_514),
.B1(n_508),
.B2(n_491),
.Y(n_549)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_482),
.Y(n_515)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_515),
.Y(n_540)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_518),
.B(n_519),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_478),
.B(n_494),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_520),
.A2(n_524),
.B(n_537),
.Y(n_555)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_521),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_504),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_522),
.B(n_523),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_485),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_490),
.A2(n_445),
.B(n_452),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_495),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_536),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_527),
.A2(n_528),
.B1(n_535),
.B2(n_496),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_497),
.B(n_492),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_502),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_470),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_531),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_480),
.A2(n_460),
.B(n_455),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_533),
.Y(n_553)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_485),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_481),
.B(n_470),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_534),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_498),
.A2(n_483),
.B1(n_475),
.B2(n_508),
.Y(n_535)
);

OAI21xp33_ASAP7_75t_L g536 ( 
.A1(n_493),
.A2(n_460),
.B(n_473),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_501),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_477),
.C(n_499),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_539),
.B(n_543),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_541),
.A2(n_556),
.B1(n_561),
.B2(n_538),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_480),
.C(n_505),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_554),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_507),
.C(n_483),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_545),
.B(n_529),
.C(n_509),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_549),
.A2(n_527),
.B1(n_523),
.B2(n_513),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_510),
.B(n_488),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_551),
.B(n_560),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_516),
.B(n_487),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_535),
.A2(n_484),
.B1(n_479),
.B2(n_474),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_518),
.B(n_465),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_559),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_526),
.B(n_454),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_526),
.B(n_411),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_453),
.B1(n_444),
.B2(n_469),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_514),
.A2(n_371),
.B1(n_387),
.B2(n_316),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_562),
.A2(n_521),
.B1(n_534),
.B2(n_531),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_512),
.B(n_387),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_512),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_565),
.B(n_579),
.Y(n_590)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_556),
.Y(n_567)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_567),
.Y(n_595)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_540),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_568),
.B(n_569),
.Y(n_594)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_547),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_553),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_570),
.B(n_571),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_532),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_555),
.A2(n_537),
.B(n_524),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_572),
.B(n_581),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_573),
.B(n_577),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_557),
.B(n_530),
.C(n_529),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_575),
.B(n_578),
.C(n_539),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_542),
.B(n_511),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_520),
.C(n_523),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_549),
.B(n_538),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_580),
.A2(n_583),
.B(n_562),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_582),
.A2(n_558),
.B1(n_548),
.B2(n_546),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_555),
.A2(n_361),
.B(n_387),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_241),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_563),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_574),
.B(n_552),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_586),
.B(n_578),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_587),
.B(n_600),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_559),
.C(n_545),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_588),
.B(n_593),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_592),
.A2(n_591),
.B1(n_600),
.B2(n_581),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_575),
.B(n_544),
.C(n_543),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_550),
.C(n_541),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_596),
.B(n_597),
.Y(n_611)
);

CKINVDCx14_ASAP7_75t_R g598 ( 
.A(n_580),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_599),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_579),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_561),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_601),
.B(n_564),
.Y(n_603)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_583),
.A2(n_319),
.B(n_377),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_602),
.A2(n_582),
.B(n_377),
.Y(n_607)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_603),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_604),
.A2(n_608),
.B1(n_609),
.B2(n_610),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_607),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_595),
.A2(n_566),
.B1(n_576),
.B2(n_584),
.Y(n_608)
);

AOI211xp5_ASAP7_75t_L g609 ( 
.A1(n_595),
.A2(n_565),
.B(n_564),
.C(n_566),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_586),
.B(n_377),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_589),
.B(n_314),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_614),
.B(n_616),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_587),
.A2(n_585),
.B(n_591),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_615),
.A2(n_593),
.B(n_590),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_588),
.B(n_314),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_606),
.B(n_594),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_617),
.B(n_610),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_611),
.B(n_596),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_618),
.B(n_621),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_619),
.A2(n_622),
.B(n_624),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_605),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_604),
.A2(n_592),
.B(n_602),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_594),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_623),
.B(n_607),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_613),
.A2(n_590),
.B(n_155),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_627),
.B(n_608),
.Y(n_630)
);

AOI31xp33_ASAP7_75t_L g639 ( 
.A1(n_630),
.A2(n_631),
.A3(n_632),
.B(n_633),
.Y(n_639)
);

XNOR2x2_ASAP7_75t_SL g632 ( 
.A(n_620),
.B(n_626),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_618),
.B(n_609),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_634),
.B(n_268),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_628),
.A2(n_625),
.B(n_627),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_635),
.A2(n_637),
.B(n_638),
.Y(n_641)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_636),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_629),
.A2(n_167),
.B(n_203),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_634),
.A2(n_203),
.B(n_219),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_640),
.B(n_639),
.C(n_152),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_641),
.B(n_205),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_205),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_141),
.Y(n_645)
);


endmodule