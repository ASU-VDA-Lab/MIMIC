module fake_jpeg_7536_n_38 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_28),
.B1(n_13),
.B2(n_27),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_18),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_21),
.B1(n_13),
.B2(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_23),
.B(n_19),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_26),
.B(n_25),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

XNOR2x1_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_14),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_14),
.B1(n_24),
.B2(n_19),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_12),
.C(n_24),
.Y(n_38)
);


endmodule