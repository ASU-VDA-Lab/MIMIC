module fake_jpeg_28404_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_71),
.Y(n_75)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_20),
.B1(n_24),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_33),
.B1(n_42),
.B2(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_28),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_33),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_24),
.B1(n_20),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_50),
.B1(n_46),
.B2(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_23),
.B1(n_16),
.B2(n_29),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_91),
.Y(n_98)
);

OAI22x1_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_44),
.B1(n_30),
.B2(n_34),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_87),
.B1(n_46),
.B2(n_66),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_42),
.B1(n_45),
.B2(n_23),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_41),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_92),
.C(n_23),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_16),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_28),
.B(n_32),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_19),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_100),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_52),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_107),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_52),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_119),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_81),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_75),
.B1(n_96),
.B2(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_51),
.B1(n_65),
.B2(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_115),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_72),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_51),
.B1(n_65),
.B2(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_124),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_74),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_32),
.B1(n_25),
.B2(n_18),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_57),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_80),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_89),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_141),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_72),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_98),
.Y(n_161)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_119),
.Y(n_162)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_106),
.B1(n_108),
.B2(n_105),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_167),
.B1(n_182),
.B2(n_134),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_108),
.C(n_105),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_168),
.C(n_170),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_114),
.B1(n_118),
.B2(n_120),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_173),
.B(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_165),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_47),
.B(n_49),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_138),
.B(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_78),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_78),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_93),
.B1(n_117),
.B2(n_88),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_41),
.C(n_79),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_41),
.C(n_55),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_104),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_104),
.B(n_1),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_123),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_178),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_0),
.B(n_2),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_2),
.B(n_3),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_29),
.B(n_30),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_74),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_128),
.B1(n_127),
.B2(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_127),
.C(n_131),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_192),
.C(n_199),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_184),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_207),
.B(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_133),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_133),
.C(n_70),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_133),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_133),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_59),
.C(n_45),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_136),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

AOI22x1_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_164),
.B1(n_158),
.B2(n_156),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_202),
.B1(n_155),
.B2(n_164),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_147),
.B1(n_88),
.B2(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_155),
.B(n_136),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_145),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_45),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_2),
.B(n_3),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_145),
.Y(n_208)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_220),
.B1(n_232),
.B2(n_186),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_30),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_170),
.B(n_173),
.Y(n_219)
);

AOI221xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_199),
.B1(n_189),
.B2(n_139),
.C(n_132),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_162),
.B1(n_160),
.B2(n_169),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_203),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_132),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_160),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_193),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_235),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_201),
.B(n_190),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_198),
.B(n_209),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_233),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_169),
.B1(n_177),
.B2(n_181),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_176),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_159),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_231),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_159),
.C(n_154),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_88),
.B(n_17),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_215),
.B1(n_232),
.B2(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_187),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_193),
.Y(n_242)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_202),
.B1(n_188),
.B2(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_227),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_207),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_252),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_255),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_132),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_249),
.B(n_250),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_22),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_31),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_256),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_212),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_2),
.B(n_3),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_234),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_17),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_4),
.B(n_5),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_230),
.C(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_265),
.C(n_269),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_271),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_259),
.B1(n_238),
.B2(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_218),
.C(n_233),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_265),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_211),
.C(n_236),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_223),
.B1(n_31),
.B2(n_22),
.Y(n_273)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_22),
.C(n_31),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_252),
.C(n_31),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

BUFx12_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_280),
.B(n_284),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_247),
.B1(n_242),
.B2(n_241),
.C(n_238),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_282),
.B(n_286),
.Y(n_307)
);

OAI211xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_259),
.B(n_246),
.C(n_257),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_283),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_251),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_264),
.B(n_270),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_245),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_259),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_271),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_262),
.C(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_298),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_263),
.B1(n_278),
.B2(n_274),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_290),
.B1(n_287),
.B2(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_304),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_285),
.B(n_293),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_10),
.C(n_5),
.Y(n_315)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_313),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_22),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.C(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_11),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_317)
);

AOI221xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_315),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_298),
.B1(n_305),
.B2(n_296),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_324),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_310),
.Y(n_322)
);

XOR2x2_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_295),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_295),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_311),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_326),
.C(n_322),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_330),
.B(n_329),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_333),
.C(n_327),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_321),
.A3(n_8),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_8),
.B1(n_15),
.B2(n_4),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_15),
.C(n_4),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_4),
.Y(n_339)
);


endmodule