module real_aes_8781_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g421 ( .A(n_0), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_1), .A2(n_137), .B(n_140), .C(n_220), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_2), .A2(n_166), .B(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g470 ( .A(n_3), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_4), .B(n_196), .Y(n_195) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_5), .A2(n_166), .B(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_L g137 ( .A(n_6), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g233 ( .A(n_7), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_8), .B(n_41), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_9), .A2(n_165), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_10), .B(n_149), .Y(n_222) );
INVx1_ASAP7_75t_L g458 ( .A(n_11), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_12), .B(n_190), .Y(n_493) );
INVx1_ASAP7_75t_L g129 ( .A(n_13), .Y(n_129) );
INVx1_ASAP7_75t_L g505 ( .A(n_14), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_15), .A2(n_78), .B1(n_110), .B2(n_111), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_16), .A2(n_174), .B(n_255), .C(n_257), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_17), .B(n_196), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_18), .B(n_436), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_19), .B(n_166), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_20), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_21), .A2(n_190), .B(n_241), .C(n_243), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_22), .B(n_196), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_23), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_24), .A2(n_176), .B(n_257), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_25), .B(n_149), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_26), .Y(n_131) );
INVx1_ASAP7_75t_L g203 ( .A(n_27), .Y(n_203) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_29), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_30), .B(n_149), .Y(n_471) );
INVx1_ASAP7_75t_L g172 ( .A(n_31), .Y(n_172) );
INVx1_ASAP7_75t_L g448 ( .A(n_32), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g106 ( .A1(n_33), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_33), .Y(n_107) );
INVx2_ASAP7_75t_L g135 ( .A(n_34), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_35), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_36), .A2(n_190), .B(n_191), .C(n_193), .Y(n_189) );
INVxp67_ASAP7_75t_L g175 ( .A(n_37), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g188 ( .A(n_38), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_39), .A2(n_140), .B(n_202), .C(n_206), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_40), .A2(n_137), .B(n_140), .C(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g447 ( .A(n_42), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_43), .A2(n_151), .B(n_231), .C(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_44), .B(n_149), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_45), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_46), .Y(n_168) );
INVx1_ASAP7_75t_L g239 ( .A(n_47), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g449 ( .A(n_48), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_49), .A2(n_58), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_49), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_50), .B(n_166), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_51), .A2(n_140), .B1(n_243), .B2(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_52), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_53), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g229 ( .A(n_54), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_55), .A2(n_193), .B(n_231), .C(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_56), .Y(n_517) );
INVx1_ASAP7_75t_L g455 ( .A(n_57), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_58), .Y(n_730) );
INVx1_ASAP7_75t_L g138 ( .A(n_59), .Y(n_138) );
INVx1_ASAP7_75t_L g128 ( .A(n_60), .Y(n_128) );
INVx1_ASAP7_75t_SL g192 ( .A(n_61), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_62), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_63), .A2(n_103), .B1(n_715), .B2(n_724), .C1(n_737), .C2(n_743), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_63), .A2(n_728), .B1(n_731), .B2(n_732), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_63), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_64), .B(n_196), .Y(n_245) );
INVx1_ASAP7_75t_L g144 ( .A(n_65), .Y(n_144) );
AOI222xp33_ASAP7_75t_SL g104 ( .A1(n_66), .A2(n_105), .B1(n_106), .B2(n_112), .C1(n_709), .C2(n_711), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_SL g435 ( .A1(n_67), .A2(n_193), .B(n_436), .C(n_437), .Y(n_435) );
INVxp67_ASAP7_75t_L g438 ( .A(n_68), .Y(n_438) );
INVx1_ASAP7_75t_L g719 ( .A(n_69), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_70), .A2(n_166), .B(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_71), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_72), .A2(n_166), .B(n_252), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_73), .Y(n_451) );
INVx1_ASAP7_75t_L g511 ( .A(n_74), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_75), .A2(n_165), .B(n_167), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_76), .Y(n_200) );
INVx1_ASAP7_75t_L g253 ( .A(n_77), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_78), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_79), .A2(n_137), .B(n_140), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_80), .A2(n_166), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g256 ( .A(n_81), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_82), .B(n_173), .Y(n_482) );
INVx2_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
INVx1_ASAP7_75t_L g221 ( .A(n_84), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_85), .B(n_436), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_86), .A2(n_137), .B(n_140), .C(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g419 ( .A(n_87), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g708 ( .A(n_87), .Y(n_708) );
OR2x2_ASAP7_75t_L g723 ( .A(n_87), .B(n_714), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_88), .A2(n_140), .B(n_143), .C(n_153), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_89), .B(n_158), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_90), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_91), .A2(n_137), .B(n_140), .C(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_92), .Y(n_497) );
INVx1_ASAP7_75t_L g434 ( .A(n_93), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_94), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_95), .B(n_173), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_96), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_97), .B(n_124), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_98), .B(n_124), .Y(n_506) );
INVx2_ASAP7_75t_L g242 ( .A(n_99), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_100), .A2(n_166), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_101), .B(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_419), .B1(n_423), .B2(n_705), .Y(n_112) );
INVx2_ASAP7_75t_L g710 ( .A(n_113), .Y(n_710) );
XOR2xp5_ASAP7_75t_L g726 ( .A(n_113), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_353), .Y(n_113) );
NAND5xp2_ASAP7_75t_L g114 ( .A(n_115), .B(n_282), .C(n_312), .D(n_333), .E(n_339), .Y(n_114) );
AOI221xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_212), .B1(n_246), .B2(n_248), .C(n_259), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_209), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_181), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_SL g333 ( .A1(n_120), .A2(n_197), .B(n_334), .C(n_337), .Y(n_333) );
AND2x2_ASAP7_75t_L g403 ( .A(n_120), .B(n_198), .Y(n_403) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_159), .Y(n_120) );
AND2x2_ASAP7_75t_L g261 ( .A(n_121), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g265 ( .A(n_121), .B(n_262), .Y(n_265) );
OR2x2_ASAP7_75t_L g291 ( .A(n_121), .B(n_198), .Y(n_291) );
AND2x2_ASAP7_75t_L g293 ( .A(n_121), .B(n_184), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_121), .B(n_183), .Y(n_311) );
INVx1_ASAP7_75t_L g344 ( .A(n_121), .Y(n_344) );
INVx2_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g211 ( .A(n_122), .Y(n_211) );
AND2x2_ASAP7_75t_L g247 ( .A(n_122), .B(n_184), .Y(n_247) );
AND2x2_ASAP7_75t_L g400 ( .A(n_122), .B(n_198), .Y(n_400) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_130), .B(n_155), .Y(n_122) );
INVx3_ASAP7_75t_L g196 ( .A(n_123), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_123), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_123), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_SL g484 ( .A(n_123), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_124), .Y(n_185) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_124), .A2(n_432), .B(n_439), .Y(n_431) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_126), .B(n_127), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_139), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_132), .A2(n_158), .B(n_200), .C(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_132), .A2(n_218), .B(n_219), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_132), .A2(n_154), .B1(n_445), .B2(n_449), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_132), .A2(n_467), .B(n_468), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_132), .A2(n_511), .B(n_512), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
AND2x4_ASAP7_75t_L g166 ( .A(n_133), .B(n_137), .Y(n_166) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g244 ( .A(n_135), .Y(n_244) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
INVx1_ASAP7_75t_L g436 ( .A(n_136), .Y(n_436) );
INVx4_ASAP7_75t_SL g154 ( .A(n_137), .Y(n_154) );
BUFx3_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
INVx5_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx3_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_148), .C(n_150), .Y(n_143) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_145), .A2(n_150), .B(n_221), .C(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_146), .A2(n_147), .B1(n_447), .B2(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx4_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx2_ASAP7_75t_L g231 ( .A(n_149), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_150), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_150), .A2(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g257 ( .A(n_152), .Y(n_257) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_154), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_154), .A2(n_169), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_SL g228 ( .A1(n_154), .A2(n_169), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_154), .A2(n_169), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_154), .A2(n_169), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_154), .A2(n_169), .B(n_434), .C(n_435), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_154), .A2(n_169), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_154), .A2(n_169), .B(n_502), .C(n_503), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_157), .A2(n_489), .B(n_496), .Y(n_488) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_158), .A2(n_227), .B(n_234), .Y(n_226) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_158), .A2(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g281 ( .A(n_159), .B(n_182), .Y(n_281) );
OR2x2_ASAP7_75t_L g285 ( .A(n_159), .B(n_198), .Y(n_285) );
AND2x2_ASAP7_75t_L g310 ( .A(n_159), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g357 ( .A(n_159), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_159), .B(n_319), .Y(n_405) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_163), .B(n_178), .Y(n_159) );
INVx1_ASAP7_75t_L g263 ( .A(n_160), .Y(n_263) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_160), .A2(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_SL g478 ( .A1(n_161), .A2(n_479), .B(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_162), .A2(n_444), .B(n_450), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_162), .B(n_451), .Y(n_450) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_162), .A2(n_466), .B(n_473), .Y(n_465) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_164), .A2(n_179), .B(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_171), .B(n_177), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_175), .B2(n_176), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_173), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_173), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_174), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_174), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_174), .B(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_176), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_176), .B(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_176), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g205 ( .A(n_177), .Y(n_205) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI322xp33_ASAP7_75t_L g406 ( .A1(n_181), .A2(n_342), .A3(n_365), .B1(n_386), .B2(n_407), .C1(n_409), .C2(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_182), .B(n_262), .Y(n_409) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_197), .Y(n_182) );
AND2x2_ASAP7_75t_L g210 ( .A(n_183), .B(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g278 ( .A(n_183), .B(n_198), .Y(n_278) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g319 ( .A(n_184), .B(n_198), .Y(n_319) );
AND2x2_ASAP7_75t_L g363 ( .A(n_184), .B(n_197), .Y(n_363) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_195), .Y(n_184) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_185), .A2(n_237), .B(n_245), .Y(n_236) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_185), .A2(n_251), .B(n_258), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_190), .B(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_194), .Y(n_494) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_196), .A2(n_453), .B(n_459), .Y(n_452) );
AND2x2_ASAP7_75t_L g246 ( .A(n_197), .B(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g264 ( .A(n_197), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_197), .B(n_293), .Y(n_417) );
INVx3_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g209 ( .A(n_198), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_198), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g331 ( .A(n_198), .B(n_262), .Y(n_331) );
AND2x2_ASAP7_75t_L g358 ( .A(n_198), .B(n_293), .Y(n_358) );
OR2x2_ASAP7_75t_L g414 ( .A(n_198), .B(n_265), .Y(n_414) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_207), .Y(n_198) );
INVx1_ASAP7_75t_SL g300 ( .A(n_209), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_210), .B(n_331), .Y(n_332) );
AND2x2_ASAP7_75t_L g366 ( .A(n_210), .B(n_356), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_210), .B(n_289), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_210), .B(n_411), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g384 ( .A1(n_212), .A2(n_246), .A3(n_385), .B(n_387), .Y(n_384) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_225), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_213), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g367 ( .A(n_213), .B(n_302), .Y(n_367) );
OR2x2_ASAP7_75t_L g374 ( .A(n_213), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g386 ( .A(n_213), .B(n_275), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g320 ( .A(n_214), .B(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g248 ( .A(n_215), .B(n_249), .Y(n_248) );
INVx4_ASAP7_75t_L g269 ( .A(n_215), .Y(n_269) );
AND2x2_ASAP7_75t_L g306 ( .A(n_215), .B(n_250), .Y(n_306) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_223), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_216), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_216), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_216), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g305 ( .A(n_225), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g375 ( .A(n_225), .Y(n_375) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_235), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_226), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g275 ( .A(n_226), .B(n_236), .Y(n_275) );
INVx2_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_226), .B(n_236), .Y(n_309) );
AND2x2_ASAP7_75t_L g316 ( .A(n_226), .B(n_272), .Y(n_316) );
BUFx3_ASAP7_75t_L g326 ( .A(n_226), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_226), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
AND2x2_ASAP7_75t_L g279 ( .A(n_235), .B(n_269), .Y(n_279) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g249 ( .A(n_236), .B(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_236), .Y(n_303) );
INVx2_ASAP7_75t_L g472 ( .A(n_243), .Y(n_472) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_SL g286 ( .A(n_247), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_247), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_247), .B(n_356), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_248), .B(n_326), .Y(n_379) );
INVx1_ASAP7_75t_SL g413 ( .A(n_248), .Y(n_413) );
INVx1_ASAP7_75t_SL g321 ( .A(n_249), .Y(n_321) );
INVx1_ASAP7_75t_SL g272 ( .A(n_250), .Y(n_272) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_250), .Y(n_283) );
OR2x2_ASAP7_75t_L g294 ( .A(n_250), .B(n_269), .Y(n_294) );
AND2x2_ASAP7_75t_L g308 ( .A(n_250), .B(n_269), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_250), .B(n_298), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_264), .B(n_266), .C(n_277), .Y(n_259) );
AOI31xp33_ASAP7_75t_L g376 ( .A1(n_260), .A2(n_377), .A3(n_378), .B(n_379), .Y(n_376) );
AND2x2_ASAP7_75t_L g349 ( .A(n_261), .B(n_278), .Y(n_349) );
BUFx3_ASAP7_75t_L g289 ( .A(n_262), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_262), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g325 ( .A(n_262), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_262), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g280 ( .A(n_265), .Y(n_280) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_265), .A2(n_390), .B1(n_393), .B2(n_394), .C1(n_395), .C2(n_396), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_267), .B(n_273), .Y(n_266) );
INVx1_ASAP7_75t_L g395 ( .A(n_267), .Y(n_395) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_269), .B(n_272), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_269), .B(n_295), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_269), .B(n_270), .Y(n_365) );
INVx1_ASAP7_75t_L g416 ( .A(n_269), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_270), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g418 ( .A(n_270), .Y(n_418) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_272), .Y(n_341) );
AOI32xp33_ASAP7_75t_L g277 ( .A1(n_273), .A2(n_278), .A3(n_279), .B1(n_280), .B2(n_281), .Y(n_277) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_275), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g352 ( .A(n_275), .Y(n_352) );
OR2x2_ASAP7_75t_L g393 ( .A(n_275), .B(n_294), .Y(n_393) );
INVx1_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_278), .B(n_289), .Y(n_314) );
INVx3_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_278), .A2(n_323), .A3(n_340), .B1(n_342), .B2(n_345), .C1(n_349), .C2(n_350), .Y(n_339) );
AND2x2_ASAP7_75t_L g315 ( .A(n_279), .B(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_L g392 ( .A(n_279), .Y(n_392) );
A2O1A1O1Ixp25_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_287), .C(n_295), .D(n_296), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_283), .B(n_326), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_285), .A2(n_297), .B1(n_300), .B2(n_301), .C(n_304), .Y(n_296) );
INVx1_ASAP7_75t_SL g411 ( .A(n_285), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B(n_294), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_289), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI221xp5_ASAP7_75t_SL g381 ( .A1(n_291), .A2(n_375), .B1(n_382), .B2(n_383), .C(n_384), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g412 ( .A1(n_292), .A2(n_413), .B1(n_414), .B2(n_415), .C1(n_417), .C2(n_418), .Y(n_412) );
AND2x2_ASAP7_75t_L g370 ( .A(n_293), .B(n_356), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_293), .A2(n_308), .B(n_355), .Y(n_382) );
INVx1_ASAP7_75t_L g396 ( .A(n_293), .Y(n_396) );
INVx2_ASAP7_75t_SL g299 ( .A(n_294), .Y(n_299) );
AND2x2_ASAP7_75t_L g302 ( .A(n_295), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_SL g336 ( .A(n_298), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_298), .B(n_308), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_299), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_299), .B(n_309), .Y(n_338) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI21xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_307), .B(n_310), .Y(n_304) );
INVx1_ASAP7_75t_SL g322 ( .A(n_306), .Y(n_322) );
AND2x2_ASAP7_75t_L g369 ( .A(n_306), .B(n_352), .Y(n_369) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g408 ( .A(n_308), .B(n_326), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_309), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g394 ( .A(n_310), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B1(n_317), .B2(n_324), .C(n_327), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B1(n_322), .B2(n_323), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_321), .A2(n_328), .B1(n_330), .B2(n_332), .Y(n_327) );
OR2x2_ASAP7_75t_L g398 ( .A(n_322), .B(n_326), .Y(n_398) );
OR2x2_ASAP7_75t_L g401 ( .A(n_322), .B(n_336), .Y(n_401) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_343), .A2(n_398), .B1(n_399), .B2(n_401), .C(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND3xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_368), .C(n_380), .Y(n_353) );
AOI222xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_359), .B1(n_361), .B2(n_364), .C1(n_366), .C2(n_367), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_356), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g378 ( .A(n_358), .Y(n_378) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_373), .C(n_376), .Y(n_368) );
INVx1_ASAP7_75t_L g383 ( .A(n_369), .Y(n_383) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g402 ( .A1(n_373), .A2(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NOR5xp2_ASAP7_75t_L g380 ( .A(n_381), .B(n_389), .C(n_397), .D(n_406), .E(n_412), .Y(n_380) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_SL g709 ( .A1(n_419), .A2(n_424), .B1(n_705), .B2(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g707 ( .A(n_420), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g714 ( .A(n_420), .Y(n_714) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_642), .Y(n_424) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_572), .C(n_603), .D(n_622), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g426 ( .A(n_427), .B(n_530), .C(n_545), .D(n_563), .Y(n_426) );
AOI222xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_475), .B1(n_507), .B2(n_518), .C1(n_523), .C2(n_525), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_460), .Y(n_428) );
INVx1_ASAP7_75t_L g586 ( .A(n_429), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_440), .Y(n_429) );
AND2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_452), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_430), .B(n_464), .Y(n_615) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g522 ( .A(n_431), .B(n_442), .Y(n_522) );
AND2x2_ASAP7_75t_L g531 ( .A(n_431), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g557 ( .A(n_431), .Y(n_557) );
AND2x2_ASAP7_75t_L g578 ( .A(n_431), .B(n_442), .Y(n_578) );
BUFx2_ASAP7_75t_L g601 ( .A(n_431), .Y(n_601) );
AND2x2_ASAP7_75t_L g625 ( .A(n_431), .B(n_443), .Y(n_625) );
AND2x2_ASAP7_75t_L g689 ( .A(n_431), .B(n_452), .Y(n_689) );
AND2x2_ASAP7_75t_L g590 ( .A(n_440), .B(n_521), .Y(n_590) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_441), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_452), .Y(n_441) );
OR2x2_ASAP7_75t_L g550 ( .A(n_442), .B(n_465), .Y(n_550) );
AND2x2_ASAP7_75t_L g562 ( .A(n_442), .B(n_521), .Y(n_562) );
BUFx2_ASAP7_75t_L g694 ( .A(n_442), .Y(n_694) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g463 ( .A(n_443), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g544 ( .A(n_443), .B(n_465), .Y(n_544) );
AND2x2_ASAP7_75t_L g597 ( .A(n_443), .B(n_452), .Y(n_597) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_443), .Y(n_633) );
AND2x2_ASAP7_75t_L g520 ( .A(n_452), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_SL g532 ( .A(n_452), .Y(n_532) );
INVx2_ASAP7_75t_L g543 ( .A(n_452), .Y(n_543) );
BUFx2_ASAP7_75t_L g567 ( .A(n_452), .Y(n_567) );
AND2x2_ASAP7_75t_SL g624 ( .A(n_452), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AOI332xp33_ASAP7_75t_L g545 ( .A1(n_461), .A2(n_546), .A3(n_550), .B1(n_551), .B2(n_555), .B3(n_558), .C1(n_559), .C2(n_561), .Y(n_545) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_461), .B(n_521), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_461), .B(n_535), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_SL g563 ( .A1(n_462), .A2(n_564), .B(n_567), .C(n_568), .Y(n_563) );
AND2x2_ASAP7_75t_L g702 ( .A(n_462), .B(n_543), .Y(n_702) );
INVx3_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g599 ( .A(n_463), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g604 ( .A(n_463), .B(n_601), .Y(n_604) );
INVx1_ASAP7_75t_L g535 ( .A(n_464), .Y(n_535) );
AND2x2_ASAP7_75t_L g638 ( .A(n_464), .B(n_597), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_464), .B(n_578), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_464), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_464), .B(n_556), .Y(n_664) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g521 ( .A(n_465), .Y(n_521) );
OAI31xp33_ASAP7_75t_L g703 ( .A1(n_475), .A2(n_624), .A3(n_631), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AND2x2_ASAP7_75t_L g507 ( .A(n_476), .B(n_508), .Y(n_507) );
NAND2x1_ASAP7_75t_SL g526 ( .A(n_476), .B(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_476), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_476), .B(n_529), .Y(n_618) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_477), .A2(n_531), .B(n_533), .C(n_536), .Y(n_530) );
OR2x2_ASAP7_75t_L g547 ( .A(n_477), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
AND2x2_ASAP7_75t_L g566 ( .A(n_477), .B(n_509), .Y(n_566) );
INVx2_ASAP7_75t_L g584 ( .A(n_477), .Y(n_584) );
AND2x2_ASAP7_75t_L g595 ( .A(n_477), .B(n_549), .Y(n_595) );
AND2x2_ASAP7_75t_L g627 ( .A(n_477), .B(n_585), .Y(n_627) );
AND2x2_ASAP7_75t_L g631 ( .A(n_477), .B(n_554), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_477), .B(n_486), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_477), .B(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_477), .B(n_573), .Y(n_704) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_484), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_486), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g612 ( .A(n_486), .Y(n_612) );
AND2x2_ASAP7_75t_L g674 ( .A(n_486), .B(n_595), .Y(n_674) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
OR2x2_ASAP7_75t_L g528 ( .A(n_487), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g538 ( .A(n_487), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_487), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g646 ( .A(n_487), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_487), .B(n_509), .Y(n_663) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g554 ( .A(n_488), .B(n_498), .Y(n_554) );
AND2x2_ASAP7_75t_L g583 ( .A(n_488), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g594 ( .A(n_488), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_488), .B(n_549), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g508 ( .A(n_499), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g529 ( .A(n_499), .Y(n_529) );
AND2x2_ASAP7_75t_L g585 ( .A(n_499), .B(n_549), .Y(n_585) );
INVx1_ASAP7_75t_L g687 ( .A(n_507), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_508), .Y(n_691) );
INVx2_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_520), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_520), .B(n_625), .Y(n_683) );
OR2x2_ASAP7_75t_L g524 ( .A(n_521), .B(n_522), .Y(n_524) );
INVx1_ASAP7_75t_SL g576 ( .A(n_521), .Y(n_576) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_527), .A2(n_580), .B1(n_582), .B2(n_586), .C(n_587), .Y(n_579) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g607 ( .A(n_528), .B(n_571), .Y(n_607) );
INVx2_ASAP7_75t_L g539 ( .A(n_529), .Y(n_539) );
INVx1_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_529), .B(n_549), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_529), .B(n_552), .Y(n_659) );
INVx1_ASAP7_75t_L g667 ( .A(n_529), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_531), .B(n_535), .Y(n_581) );
AND2x4_ASAP7_75t_L g556 ( .A(n_532), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g669 ( .A(n_535), .B(n_625), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_538), .B(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g677 ( .A(n_539), .Y(n_677) );
INVxp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g577 ( .A(n_543), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g649 ( .A(n_543), .B(n_625), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_543), .B(n_562), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g609 ( .A1(n_544), .A2(n_578), .A3(n_585), .B1(n_610), .B2(n_613), .C1(n_614), .C2(n_616), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_544), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g675 ( .A(n_547), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g621 ( .A(n_548), .Y(n_621) );
INVx2_ASAP7_75t_L g552 ( .A(n_549), .Y(n_552) );
INVx1_ASAP7_75t_L g611 ( .A(n_549), .Y(n_611) );
CKINVDCx16_ASAP7_75t_R g558 ( .A(n_550), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g647 ( .A(n_552), .B(n_560), .Y(n_647) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g559 ( .A(n_554), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g602 ( .A(n_554), .B(n_595), .Y(n_602) );
AND2x2_ASAP7_75t_L g606 ( .A(n_554), .B(n_566), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_555), .A2(n_617), .B(n_619), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_555), .A2(n_687), .B1(n_688), .B2(n_690), .Y(n_686) );
INVx3_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g561 ( .A(n_556), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_556), .B(n_576), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_558), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g698 ( .A(n_565), .Y(n_698) );
INVx4_ASAP7_75t_L g571 ( .A(n_566), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_566), .B(n_593), .Y(n_641) );
INVx1_ASAP7_75t_SL g653 ( .A(n_567), .Y(n_653) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_571), .B(n_667), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B(n_579), .C(n_596), .Y(n_572) );
OAI221xp5_ASAP7_75t_SL g692 ( .A1(n_574), .A2(n_612), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_692) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_576), .B(n_689), .Y(n_688) );
OAI31xp33_ASAP7_75t_L g668 ( .A1(n_577), .A2(n_654), .A3(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g608 ( .A(n_578), .Y(n_608) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g658 ( .A(n_583), .Y(n_658) );
AND2x2_ASAP7_75t_L g671 ( .A(n_585), .B(n_594), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_595), .B(n_698), .Y(n_697) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI221xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B1(n_607), .B2(n_608), .C(n_609), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_604), .A2(n_673), .B(n_675), .C(n_678), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_607), .B(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g634 ( .A(n_615), .Y(n_634) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g620 ( .A(n_618), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g662 ( .A(n_618), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_628), .C(n_637), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_626), .A2(n_636), .B1(n_700), .B2(n_701), .C(n_703), .Y(n_699) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_632), .B2(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_SL g700 ( .A(n_639), .Y(n_700) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR4xp25_ASAP7_75t_L g642 ( .A(n_643), .B(n_672), .C(n_692), .D(n_699), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B(n_650), .C(n_668), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B(n_656), .C(n_660), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g679 ( .A(n_657), .Y(n_679) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OR2x2_ASAP7_75t_L g690 ( .A(n_658), .B(n_691), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_684), .C(n_686), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_689), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NOR2x2_ASAP7_75t_L g713 ( .A(n_708), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .Y(n_716) );
NOR2xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_SL g742 ( .A(n_718), .Y(n_742) );
INVx1_ASAP7_75t_L g741 ( .A(n_720), .Y(n_741) );
OA21x2_ASAP7_75t_L g744 ( .A1(n_720), .A2(n_742), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_723), .Y(n_733) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_723), .Y(n_735) );
BUFx2_ASAP7_75t_L g745 ( .A(n_723), .Y(n_745) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_733), .B(n_734), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_728), .Y(n_732) );
NOR2xp33_ASAP7_75t_SL g734 ( .A(n_735), .B(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
CKINVDCx6p67_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
endmodule