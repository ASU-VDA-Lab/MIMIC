module fake_jpeg_25403_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_23),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_16),
.B1(n_10),
.B2(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_5),
.CI(n_6),
.CON(n_23),
.SN(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_10),
.C(n_18),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_22),
.B(n_1),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_41),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_16),
.B1(n_10),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_40),
.B1(n_34),
.B2(n_32),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_0),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_36),
.B1(n_40),
.B2(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_48),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_23),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_53),
.C(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_9),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_35),
.C(n_17),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_51),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_47),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.C(n_9),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_7),
.B1(n_32),
.B2(n_44),
.Y(n_61)
);


endmodule