module fake_jpeg_16415_n_358 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_36),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_37),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_46),
.B(n_30),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_22),
.B1(n_37),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_73),
.B1(n_41),
.B2(n_29),
.Y(n_92)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_0),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_27),
.B1(n_33),
.B2(n_26),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_26),
.B1(n_35),
.B2(n_27),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_52),
.B1(n_42),
.B2(n_14),
.Y(n_87)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_50),
.Y(n_91)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx2_ASAP7_75t_SL g125 ( 
.A(n_85),
.Y(n_125)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_86),
.B(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_32),
.B1(n_34),
.B2(n_30),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_62),
.B(n_11),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_103),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_45),
.B1(n_53),
.B2(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_107),
.B1(n_99),
.B2(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_20),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_45),
.B1(n_51),
.B2(n_34),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_73),
.B(n_65),
.C(n_62),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_135),
.B(n_32),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_123),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_34),
.B(n_28),
.C(n_30),
.Y(n_147)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_69),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_40),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_72),
.Y(n_162)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_55),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_66),
.B1(n_63),
.B2(n_59),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_109),
.B1(n_100),
.B2(n_88),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_161)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_88),
.A2(n_83),
.B1(n_112),
.B2(n_81),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_83),
.B1(n_80),
.B2(n_59),
.Y(n_150)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_150),
.B1(n_159),
.B2(n_161),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_162),
.B(n_163),
.Y(n_186)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_118),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_111),
.B1(n_94),
.B2(n_93),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_164),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_137),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_111),
.B1(n_76),
.B2(n_108),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_134),
.B1(n_141),
.B2(n_115),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_55),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_135),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_80),
.B1(n_85),
.B2(n_29),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_168),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_55),
.B(n_1),
.Y(n_163)
);

AOI22x1_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_104),
.B1(n_89),
.B2(n_21),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_166),
.B(n_167),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_36),
.B(n_29),
.C(n_32),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_38),
.Y(n_168)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_171),
.A2(n_181),
.B(n_132),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_128),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_117),
.C(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_139),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_136),
.B1(n_137),
.B2(n_115),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_163),
.B1(n_147),
.B2(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

XNOR2x2_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_144),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_152),
.B(n_132),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_143),
.C(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_192),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_120),
.B1(n_129),
.B2(n_121),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_167),
.B(n_147),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_211),
.B1(n_180),
.B2(n_184),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_195),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_214),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_147),
.B1(n_155),
.B2(n_153),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_208),
.B1(n_216),
.B2(n_28),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_148),
.B(n_145),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_210),
.A2(n_219),
.B1(n_172),
.B2(n_192),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_161),
.B1(n_146),
.B2(n_130),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_122),
.B1(n_120),
.B2(n_130),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_208),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_20),
.B(n_38),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_20),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_222),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_177),
.C(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_184),
.C(n_188),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_195),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_181),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_243),
.C(n_203),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_193),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_241),
.B1(n_244),
.B2(n_216),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_182),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_239),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_206),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_218),
.C(n_200),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_196),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_207),
.B(n_222),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_252),
.A2(n_258),
.B(n_259),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_219),
.C(n_196),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_232),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_264),
.B1(n_212),
.B2(n_4),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_197),
.B(n_215),
.Y(n_259)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_263),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_214),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_199),
.C(n_213),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_237),
.C(n_225),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_241),
.B(n_236),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_213),
.B1(n_199),
.B2(n_201),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_258),
.B1(n_265),
.B2(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_252),
.B(n_270),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_275),
.B(n_281),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_287),
.C(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_247),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_221),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_288),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_259),
.A2(n_246),
.B(n_201),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_28),
.B1(n_19),
.B2(n_3),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_268),
.B1(n_269),
.B2(n_248),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_38),
.C(n_19),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_38),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_19),
.C(n_4),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_253),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_275),
.C(n_288),
.Y(n_315)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_272),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_279),
.B(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_287),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_274),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_312),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_280),
.B1(n_249),
.B2(n_283),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_311),
.A2(n_310),
.B1(n_317),
.B2(n_256),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_301),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_282),
.B(n_285),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_294),
.B(n_295),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_306),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_281),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_302),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_320),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_327),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_329),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_314),
.A2(n_294),
.B1(n_293),
.B2(n_249),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_8),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_326),
.C(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_286),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_330),
.B(n_331),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_253),
.B1(n_6),
.B2(n_7),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_5),
.C(n_7),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_318),
.B1(n_315),
.B2(n_312),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_337),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_338),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_5),
.C(n_7),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_8),
.B(n_9),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_10),
.B(n_11),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_9),
.Y(n_342)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_342),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_343),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_324),
.C(n_321),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_345),
.A2(n_346),
.B(n_340),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_349),
.B(n_340),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_352),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_347),
.B(n_327),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_341),
.B(n_13),
.C(n_14),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_355),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_10),
.B(n_13),
.Y(n_357)
);

AO22x1_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_16),
.B1(n_17),
.B2(n_350),
.Y(n_358)
);


endmodule