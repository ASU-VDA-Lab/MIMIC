module fake_jpeg_20237_n_24 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_24;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

AOI22xp33_ASAP7_75t_L g11 ( 
.A1(n_8),
.A2(n_3),
.B1(n_2),
.B2(n_9),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NAND3xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_3),
.C(n_6),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_10),
.C(n_1),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_17),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_0),
.B(n_2),
.Y(n_16)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_4),
.C(n_5),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_4),
.B(n_5),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_18),
.A2(n_20),
.B(n_6),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_12),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_21),
.Y(n_24)
);


endmodule