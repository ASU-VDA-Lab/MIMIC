module fake_jpeg_2665_n_173 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_0),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_43),
.B1(n_58),
.B2(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_72),
.B1(n_73),
.B2(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_58),
.B1(n_44),
.B2(n_53),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_47),
.B1(n_45),
.B2(n_51),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_56),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_3),
.B(n_4),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_48),
.B1(n_56),
.B2(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_55),
.B1(n_52),
.B2(n_5),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_89),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_0),
.C(n_2),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_3),
.Y(n_105)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_106),
.B1(n_109),
.B2(n_13),
.Y(n_128)
);

OAI21x1_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_105),
.B(n_78),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_23),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_110),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_7),
.Y(n_110)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_90),
.Y(n_118)
);

NOR2x1_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_9),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_10),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_11),
.B(n_12),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_112),
.B(n_15),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_29),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_12),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_13),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_20),
.C1(n_22),
.C2(n_26),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_31),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_124),
.C(n_116),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_137),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_138),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_112),
.B(n_14),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_144),
.B(n_147),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_41),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_27),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_122),
.B1(n_117),
.B2(n_125),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g154 ( 
.A(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_146),
.C(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_158),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_133),
.C(n_139),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_144),
.C(n_136),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_149),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_154),
.B1(n_149),
.B2(n_137),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_162),
.B1(n_158),
.B2(n_160),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_135),
.A3(n_147),
.B1(n_164),
.B2(n_151),
.C1(n_35),
.C2(n_30),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_32),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_167),
.B1(n_147),
.B2(n_37),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_33),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_147),
.Y(n_173)
);


endmodule