module fake_netlist_6_1801_n_107 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_0, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_107);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_0;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_107;

wire n_52;
wire n_91;
wire n_46;
wire n_88;
wire n_98;
wire n_63;
wire n_39;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_100;
wire n_47;
wire n_62;
wire n_75;
wire n_45;
wire n_70;
wire n_67;
wire n_82;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_69;
wire n_79;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_8),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_L g49 ( 
.A(n_3),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_0),
.B(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_R g57 ( 
.A(n_2),
.B(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_R g59 ( 
.A(n_2),
.B(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_23),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_R g70 ( 
.A(n_53),
.B(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_15),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_42),
.B(n_43),
.C(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_48),
.B(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_65),
.B1(n_64),
.B2(n_63),
.Y(n_84)
);

OA21x2_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_58),
.B(n_47),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_87)
);

OAI221xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_70),
.B1(n_73),
.B2(n_55),
.C(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_78),
.A3(n_60),
.B1(n_44),
.B2(n_54),
.C(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_74),
.Y(n_92)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_49),
.B(n_39),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_69),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_83),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_86),
.C(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_83),
.Y(n_100)
);

NAND4xp25_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_91),
.C(n_81),
.D(n_93),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_93),
.B1(n_83),
.B2(n_56),
.C(n_38),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_96),
.B1(n_98),
.B2(n_51),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI222xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_61),
.B1(n_81),
.B2(n_85),
.C1(n_103),
.C2(n_88),
.Y(n_107)
);


endmodule