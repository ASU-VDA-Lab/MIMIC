module real_jpeg_11403_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_238;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_202;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_27),
.B(n_33),
.C(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_3),
.B(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_28),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_3),
.A2(n_28),
.B(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_62),
.C(n_67),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_38),
.B1(n_47),
.B2(n_51),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_83),
.B1(n_84),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_3),
.B(n_111),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_47),
.B1(n_51),
.B2(n_54),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_5),
.A2(n_54),
.B1(n_66),
.B2(n_67),
.Y(n_170)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_7),
.A2(n_47),
.B1(n_51),
.B2(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_87),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_87),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_8),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_8),
.A2(n_47),
.B1(n_51),
.B2(n_89),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_89),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_47),
.B1(n_51),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_72),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_13),
.A2(n_47),
.B1(n_51),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_13),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_75),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_75),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_75),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_14),
.A2(n_41),
.B1(n_47),
.B2(n_51),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_41),
.B1(n_66),
.B2(n_67),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_15),
.A2(n_47),
.B1(n_51),
.B2(n_56),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_15),
.A2(n_56),
.B1(n_66),
.B2(n_67),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_277),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_255),
.B(n_276),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_228),
.B(n_254),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_123),
.B(n_204),
.C(n_227),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_21),
.B(n_102),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_93),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_57),
.C(n_77),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_24),
.B(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_25),
.A2(n_26),
.B1(n_106),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_25),
.A2(n_221),
.B(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_25),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_26),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_28),
.A2(n_31),
.B(n_38),
.Y(n_92)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g141 ( 
.A(n_29),
.B(n_49),
.C(n_51),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_38),
.B(n_84),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_38),
.B(n_65),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_42),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_42),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_45),
.A2(n_55),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_45),
.A2(n_46),
.B1(n_101),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_45),
.A2(n_110),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_45),
.A2(n_223),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_46),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_47),
.A2(n_50),
.B(n_139),
.C(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_47),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_70),
.B(n_73),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_59),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_59),
.A2(n_65),
.B(n_70),
.Y(n_288)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_74),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_60),
.A2(n_76),
.B1(n_134),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_60),
.A2(n_76),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_60),
.A2(n_76),
.B1(n_157),
.B2(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_60),
.A2(n_76),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_60),
.A2(n_214),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_66),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_84),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_76),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_73),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_79),
.B1(n_93),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_90),
.B2(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_90),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_82),
.A2(n_121),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_82),
.A2(n_85),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_83),
.A2(n_84),
.B1(n_170),
.B2(n_178),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_83),
.A2(n_172),
.B(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_83),
.A2(n_84),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_86),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_85),
.B(n_144),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_96),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_103),
.B(n_114),
.C(n_122),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_105),
.B(n_107),
.C(n_112),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_111),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_111),
.A2(n_247),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_115),
.B(n_118),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_116),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_117),
.B(n_135),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_202),
.B(n_203),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_145),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_126),
.B(n_129),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_136),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_142),
.B1(n_143),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_158),
.B(n_201),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_195),
.B(n_200),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_184),
.B(n_194),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_173),
.B(n_183),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_168),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_165),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_179),
.B(n_182),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_190),
.C(n_193),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_226),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_226),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.C(n_216),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_215),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_219),
.C(n_225),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_225),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_253),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_239),
.B1(n_251),
.B2(n_252),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_252),
.C(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_233),
.A2(n_234),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_236),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_234),
.A2(n_267),
.B(n_269),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_244),
.C(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_245),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_275),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_275),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_274),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_260),
.C(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_264),
.B(n_265),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_281),
.CI(n_282),
.CON(n_280),
.SN(n_280)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_294),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_280),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_280),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_290),
.B2(n_293),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);


endmodule