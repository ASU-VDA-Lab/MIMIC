module fake_jpeg_1869_n_223 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_223);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_49),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_0),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_67),
.Y(n_88)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_63),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_73),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_68),
.B1(n_58),
.B2(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_77),
.B1(n_68),
.B2(n_55),
.Y(n_114)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_80),
.B1(n_51),
.B2(n_58),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_83),
.B1(n_78),
.B2(n_84),
.Y(n_112)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_76),
.B1(n_50),
.B2(n_66),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_116),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_77),
.C(n_54),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_113),
.Y(n_124)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_97),
.CON(n_111),
.SN(n_111)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_112),
.Y(n_132)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_76),
.B1(n_91),
.B2(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_118),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_99),
.B1(n_85),
.B2(n_77),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_139),
.B1(n_119),
.B2(n_133),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_125),
.B1(n_133),
.B2(n_3),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_66),
.B1(n_73),
.B2(n_59),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_57),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_135),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_72),
.B1(n_59),
.B2(n_60),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_74),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_84),
.B(n_86),
.C(n_60),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_144),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_117),
.C(n_62),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_142),
.C(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_103),
.C(n_53),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_75),
.B(n_71),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_153),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_138),
.B(n_121),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_152),
.B(n_156),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_118),
.C(n_65),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_31),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_102),
.B(n_65),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_61),
.B1(n_57),
.B2(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_158),
.B1(n_164),
.B2(n_12),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_61),
.B(n_40),
.C(n_35),
.D(n_32),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_1),
.B(n_2),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_8),
.C(n_9),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_3),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_154),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_7),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_30),
.A3(n_29),
.B1(n_28),
.B2(n_26),
.C1(n_25),
.C2(n_18),
.Y(n_178)
);

OAI321xp33_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_156),
.A3(n_17),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_160),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_24),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_16),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_151),
.C(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_188),
.C(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_149),
.C(n_152),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_16),
.CI(n_17),
.CON(n_196),
.SN(n_196)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_197),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_21),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_176),
.B(n_181),
.Y(n_202)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_179),
.C(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_201),
.B(n_207),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_172),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_168),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_170),
.C(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_168),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_203),
.C(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_210),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_192),
.C(n_190),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_202),
.Y(n_216)
);

OAI21x1_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_216),
.B(n_208),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_218),
.B1(n_206),
.B2(n_194),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_211),
.A3(n_200),
.B1(n_206),
.B2(n_196),
.C1(n_212),
.C2(n_177),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_181),
.B(n_175),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_181),
.C(n_22),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_22),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_23),
.Y(n_223)
);


endmodule