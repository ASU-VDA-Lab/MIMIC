module fake_jpeg_2467_n_230 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_24),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_73),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_85),
.Y(n_105)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_63),
.B1(n_72),
.B2(n_58),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_86),
.B1(n_95),
.B2(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_108),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_0),
.C(n_1),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_81),
.B(n_86),
.C(n_53),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_59),
.B(n_62),
.C(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_66),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_55),
.B1(n_65),
.B2(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_64),
.B1(n_56),
.B2(n_57),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx4f_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_54),
.B1(n_60),
.B2(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_91),
.B1(n_56),
.B2(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_96),
.B1(n_92),
.B2(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_130),
.B1(n_107),
.B2(n_67),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_128),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_132),
.B1(n_3),
.B2(n_5),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_138),
.B1(n_92),
.B2(n_78),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_75),
.B1(n_69),
.B2(n_61),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_117),
.B1(n_106),
.B2(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_139),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_75),
.B1(n_69),
.B2(n_79),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_76),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_96),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_151),
.B1(n_157),
.B2(n_158),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_67),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_78),
.B1(n_92),
.B2(n_81),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_11),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_51),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_136),
.B(n_141),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_153),
.B(n_155),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_0),
.B(n_2),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_26),
.B1(n_49),
.B2(n_48),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_28),
.C(n_45),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_6),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_8),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_167),
.B1(n_13),
.B2(n_14),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_44),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_160),
.C(n_163),
.Y(n_191)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_183),
.B1(n_157),
.B2(n_155),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_153),
.B(n_160),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_196),
.C(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_194),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_145),
.C(n_34),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_15),
.B(n_17),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_168),
.B(n_173),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_35),
.C(n_23),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_199),
.B(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_178),
.C(n_186),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_204),
.C(n_209),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_185),
.C(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_207),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_197),
.B1(n_189),
.B2(n_193),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_174),
.C(n_172),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_213),
.B(n_216),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_188),
.B1(n_171),
.B2(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_193),
.B1(n_179),
.B2(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_201),
.A3(n_175),
.B1(n_200),
.B2(n_32),
.C1(n_33),
.C2(n_37),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_217),
.C(n_211),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_211),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_221),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_43),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_25),
.B(n_30),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_40),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_41),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_42),
.Y(n_230)
);


endmodule