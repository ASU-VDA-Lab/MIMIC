module fake_netlist_1_8446_n_1042 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1042);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1042;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_947;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_189), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_197), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_20), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_235), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_34), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_32), .B(n_65), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_49), .Y(n_251) );
BUFx8_ASAP7_75t_SL g252 ( .A(n_209), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_224), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_13), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_225), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_78), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_79), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_236), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_202), .Y(n_259) );
BUFx10_ASAP7_75t_L g260 ( .A(n_13), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_126), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_219), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_38), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_74), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_93), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_124), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_186), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_106), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_214), .Y(n_270) );
BUFx8_ASAP7_75t_SL g271 ( .A(n_73), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_200), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_159), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_192), .Y(n_275) );
BUFx5_ASAP7_75t_L g276 ( .A(n_227), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_154), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_162), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_96), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_195), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_134), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_49), .Y(n_282) );
CKINVDCx16_ASAP7_75t_R g283 ( .A(n_122), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_72), .Y(n_284) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_125), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_145), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_201), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_131), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_66), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_156), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_92), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_217), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_164), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_62), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_36), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_215), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_54), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_198), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_136), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_23), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_223), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_66), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_38), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_50), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_158), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_205), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_161), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_85), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_119), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_127), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_233), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_8), .Y(n_312) );
CKINVDCx14_ASAP7_75t_R g313 ( .A(n_221), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_163), .Y(n_314) );
INVxp67_ASAP7_75t_SL g315 ( .A(n_204), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_226), .Y(n_316) );
INVxp33_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_41), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_203), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_76), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_7), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_187), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_18), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_199), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_15), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_210), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_167), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_52), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_123), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_95), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_138), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_180), .Y(n_333) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_139), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_181), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_178), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_116), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_168), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_92), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_98), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_185), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_95), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_100), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_108), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_232), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_182), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_207), .Y(n_347) );
NOR2xp67_ASAP7_75t_L g348 ( .A(n_9), .B(n_141), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_40), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_193), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_160), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_144), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_35), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_64), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_71), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_58), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_220), .Y(n_357) );
CKINVDCx14_ASAP7_75t_R g358 ( .A(n_129), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_133), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_179), .Y(n_360) );
BUFx8_ASAP7_75t_SL g361 ( .A(n_137), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_194), .Y(n_362) );
BUFx10_ASAP7_75t_L g363 ( .A(n_212), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_240), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_103), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_213), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_102), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_7), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_18), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_31), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_25), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_211), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_140), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_155), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_208), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_27), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_135), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_23), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_278), .A2(n_110), .B(n_109), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_278), .A2(n_112), .B(n_111), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
INVx4_ASAP7_75t_L g382 ( .A(n_272), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_269), .B(n_0), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_276), .Y(n_384) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_363), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_269), .B(n_0), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_243), .A2(n_114), .B(n_113), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_318), .B(n_1), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_251), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_341), .Y(n_392) );
INVx4_ASAP7_75t_L g393 ( .A(n_293), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_276), .B(n_1), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_276), .Y(n_397) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_318), .B(n_2), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_251), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_252), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_254), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_276), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_254), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_247), .A2(n_117), .B(n_115), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_344), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_276), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_249), .A2(n_120), .B(n_118), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_258), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_339), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_341), .Y(n_410) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_345), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_345), .Y(n_412) );
INVx5_ASAP7_75t_L g413 ( .A(n_345), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_291), .B(n_5), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_276), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_317), .B(n_6), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_352), .Y(n_418) );
AND2x6_ASAP7_75t_L g419 ( .A(n_275), .B(n_121), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_352), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_346), .B(n_6), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_382), .B(n_317), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_384), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_386), .B(n_283), .Y(n_430) );
BUFx10_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
AND2x6_ASAP7_75t_L g434 ( .A(n_383), .B(n_275), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_386), .Y(n_435) );
NAND2xp33_ASAP7_75t_L g436 ( .A(n_419), .B(n_244), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
AND3x1_ASAP7_75t_L g438 ( .A(n_405), .B(n_246), .C(n_257), .Y(n_438) );
NAND2xp33_ASAP7_75t_SL g439 ( .A(n_400), .B(n_258), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_402), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_396), .B(n_285), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_414), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_406), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_396), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_406), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_417), .A2(n_306), .B1(n_311), .B2(n_262), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
BUFx6f_ASAP7_75t_SL g450 ( .A(n_383), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_382), .B(n_334), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_396), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_382), .B(n_313), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_381), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_408), .B(n_264), .C(n_308), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_381), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_393), .B(n_255), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
AND3x2_ASAP7_75t_L g459 ( .A(n_417), .B(n_274), .C(n_271), .Y(n_459) );
NAND2xp33_ASAP7_75t_L g460 ( .A(n_419), .B(n_245), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_388), .Y(n_461) );
BUFx6f_ASAP7_75t_SL g462 ( .A(n_383), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_448), .A2(n_405), .B1(n_408), .B2(n_393), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_443), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_453), .B(n_393), .Y(n_465) );
INVx8_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_431), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_434), .A2(n_390), .B1(n_387), .B2(n_414), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_430), .B(n_393), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_443), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_423), .B(n_387), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_443), .B(n_387), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_443), .B(n_387), .Y(n_473) );
BUFx6f_ASAP7_75t_SL g474 ( .A(n_434), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_431), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_441), .A2(n_385), .B1(n_390), .B2(n_421), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_438), .A2(n_306), .B1(n_311), .B2(n_262), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_431), .B(n_385), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_457), .B(n_390), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_455), .A2(n_390), .B1(n_414), .B2(n_351), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_442), .B(n_414), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_451), .B(n_253), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_434), .B(n_415), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_436), .A2(n_380), .B(n_379), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_434), .B(n_398), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_434), .B(n_398), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_422), .A2(n_404), .B(n_407), .C(n_389), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_435), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_446), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_460), .B(n_395), .C(n_256), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_422), .B(n_259), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_424), .A2(n_380), .B(n_379), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_429), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_424), .B(n_425), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_428), .B(n_419), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_462), .B(n_313), .Y(n_498) );
OR2x6_ASAP7_75t_L g499 ( .A(n_459), .B(n_389), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_438), .A2(n_351), .B1(n_267), .B2(n_280), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_448), .B(n_370), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_447), .A2(n_380), .B(n_379), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_437), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_449), .B(n_358), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_449), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_458), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_440), .B(n_391), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_444), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_444), .A2(n_419), .B1(n_266), .B2(n_279), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_445), .B(n_315), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_445), .B(n_391), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_439), .B(n_268), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_427), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_426), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_432), .A2(n_373), .B1(n_319), .B2(n_265), .Y(n_516) );
INVx8_ASAP7_75t_L g517 ( .A(n_426), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_426), .B(n_270), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_433), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_433), .B(n_327), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_461), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_454), .B(n_399), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_454), .A2(n_380), .B(n_379), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_454), .B(n_260), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_456), .B(n_399), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_466), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_465), .B(n_248), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_495), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_465), .B(n_284), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_495), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_466), .B(n_273), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_484), .A2(n_473), .B(n_472), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_481), .B(n_289), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_472), .A2(n_404), .B(n_389), .Y(n_534) );
INVx3_ASAP7_75t_SL g535 ( .A(n_466), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_473), .A2(n_407), .B(n_404), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_493), .A2(n_502), .B(n_471), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_479), .B(n_294), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_469), .B(n_300), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_468), .A2(n_295), .B(n_297), .C(n_282), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_464), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_480), .A2(n_344), .B1(n_303), .B2(n_321), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_470), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_506), .A2(n_325), .B(n_329), .C(n_312), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_501), .B(n_260), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_463), .A2(n_343), .B1(n_355), .B2(n_340), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_503), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_497), .A2(n_263), .B(n_261), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_474), .A2(n_368), .B1(n_378), .B2(n_369), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_509), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_482), .B(n_302), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_513), .B(n_323), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_467), .B(n_277), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_483), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_524), .B(n_331), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_508), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_496), .B(n_367), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_509), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_505), .A2(n_288), .B(n_286), .Y(n_560) );
NOR2x1_ASAP7_75t_R g561 ( .A(n_477), .B(n_342), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_507), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_475), .B(n_281), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_474), .A2(n_250), .B1(n_376), .B2(n_356), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_511), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_485), .B(n_354), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_509), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_486), .B(n_365), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_500), .A2(n_371), .B1(n_304), .B2(n_320), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_511), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_488), .A2(n_299), .B(n_298), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_486), .B(n_309), .C(n_305), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_478), .B(n_401), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_516), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_491), .B(n_328), .C(n_324), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_489), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_492), .B(n_361), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_520), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_490), .A2(n_521), .B(n_504), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_494), .A2(n_336), .B(n_332), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_499), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_499), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_498), .B(n_403), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_522), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_525), .A2(n_348), .B(n_337), .C(n_347), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_510), .B(n_287), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_518), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_514), .A2(n_360), .B(n_364), .C(n_357), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_519), .B(n_339), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_517), .B(n_301), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_515), .B(n_339), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_515), .A2(n_338), .B(n_330), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_469), .B(n_339), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_466), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_476), .B(n_290), .Y(n_597) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_523), .A2(n_409), .B(n_420), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_463), .A2(n_353), .B1(n_409), .B2(n_296), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_465), .B(n_292), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_466), .Y(n_601) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_523), .A2(n_409), .B(n_413), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_463), .A2(n_409), .B(n_353), .C(n_10), .Y(n_603) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_468), .A2(n_310), .B(n_307), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_SL g605 ( .A1(n_487), .A2(n_130), .B(n_132), .C(n_128), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_463), .A2(n_316), .B1(n_322), .B2(n_314), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_463), .A2(n_333), .B1(n_335), .B2(n_326), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_495), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_495), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_468), .A2(n_353), .B1(n_374), .B2(n_352), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_501), .B(n_8), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_465), .B(n_350), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_484), .A2(n_362), .B(n_359), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_465), .B(n_366), .Y(n_614) );
O2A1O1Ixp5_ASAP7_75t_L g615 ( .A1(n_484), .A2(n_375), .B(n_377), .C(n_372), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_495), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_466), .B(n_374), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_484), .A2(n_392), .B(n_388), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_484), .A2(n_392), .B(n_388), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_493), .A2(n_392), .B(n_388), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_503), .Y(n_621) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_598), .A2(n_411), .B(n_410), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_538), .B(n_9), .Y(n_623) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_537), .A2(n_411), .B(n_410), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_528), .B(n_10), .Y(n_625) );
NAND3xp33_ASAP7_75t_SL g626 ( .A(n_599), .B(n_11), .C(n_12), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_532), .A2(n_411), .B(n_410), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_530), .B(n_11), .Y(n_628) );
AO21x2_ASAP7_75t_L g629 ( .A1(n_620), .A2(n_411), .B(n_410), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_608), .B(n_12), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_609), .B(n_14), .Y(n_631) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_602), .A2(n_416), .B(n_412), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_616), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_535), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_570), .A2(n_416), .B1(n_418), .B2(n_412), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_603), .A2(n_416), .B(n_418), .C(n_412), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_573), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_526), .B(n_418), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_601), .B(n_14), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_562), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_560), .A2(n_418), .B(n_19), .C(n_16), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_565), .A2(n_20), .B(n_16), .C(n_17), .Y(n_642) );
INVx5_ASAP7_75t_L g643 ( .A(n_596), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_591), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_561), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_557), .B(n_21), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_534), .A2(n_143), .B(n_142), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_548), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_546), .B(n_21), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_595), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_596), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_585), .A2(n_22), .B(n_24), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_576), .A2(n_25), .B(n_22), .C(n_24), .Y(n_653) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_550), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_536), .A2(n_147), .B(n_146), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_613), .A2(n_149), .B(n_148), .Y(n_656) );
O2A1O1Ixp5_ASAP7_75t_L g657 ( .A1(n_615), .A2(n_151), .B(n_152), .C(n_150), .Y(n_657) );
BUFx12f_ASAP7_75t_L g658 ( .A(n_583), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_543), .B(n_26), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_549), .A2(n_157), .B(n_153), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_542), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_543), .B(n_27), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_611), .B(n_28), .Y(n_663) );
OR2x6_ASAP7_75t_L g664 ( .A(n_584), .B(n_29), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_547), .B(n_29), .Y(n_665) );
INVx4_ASAP7_75t_L g666 ( .A(n_548), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_580), .A2(n_30), .B1(n_32), .B2(n_33), .Y(n_667) );
OAI21x1_ASAP7_75t_L g668 ( .A1(n_594), .A2(n_166), .B(n_165), .Y(n_668) );
BUFx2_ASAP7_75t_R g669 ( .A(n_531), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_547), .B(n_33), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_581), .A2(n_171), .B(n_170), .Y(n_671) );
NOR2xp33_ASAP7_75t_SL g672 ( .A(n_548), .B(n_172), .Y(n_672) );
AO31x2_ASAP7_75t_L g673 ( .A1(n_610), .A2(n_34), .A3(n_36), .B(n_37), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_555), .Y(n_674) );
AO31x2_ASAP7_75t_L g675 ( .A1(n_610), .A2(n_37), .A3(n_39), .B(n_40), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g676 ( .A1(n_590), .A2(n_41), .B(n_42), .C(n_43), .Y(n_676) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_567), .A2(n_174), .B(n_173), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_578), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_574), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_541), .B(n_44), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_575), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_681) );
OAI21x1_ASAP7_75t_L g682 ( .A1(n_567), .A2(n_177), .B(n_176), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_606), .B(n_47), .C(n_48), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_539), .B(n_48), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_527), .B(n_529), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_555), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_558), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_544), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_558), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_584), .B(n_51), .Y(n_690) );
O2A1O1Ixp5_ASAP7_75t_L g691 ( .A1(n_617), .A2(n_191), .B(n_242), .C(n_241), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_600), .A2(n_190), .B(n_238), .Y(n_692) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_545), .A2(n_53), .B(n_55), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_551), .B(n_55), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_533), .B(n_56), .Y(n_695) );
AO32x2_ASAP7_75t_L g696 ( .A1(n_564), .A2(n_56), .A3(n_57), .B1(n_58), .B2(n_59), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_559), .Y(n_697) );
AO31x2_ASAP7_75t_L g698 ( .A1(n_587), .A2(n_57), .A3(n_59), .B(n_60), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_586), .Y(n_699) );
INVx4_ASAP7_75t_L g700 ( .A(n_621), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_572), .A2(n_188), .B(n_234), .Y(n_701) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_593), .Y(n_702) );
AOI211x1_ASAP7_75t_L g703 ( .A1(n_582), .A2(n_60), .B(n_61), .C(n_62), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_589), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_607), .B(n_61), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_556), .B(n_63), .Y(n_706) );
INVx8_ASAP7_75t_L g707 ( .A(n_569), .Y(n_707) );
INVx6_ASAP7_75t_SL g708 ( .A(n_579), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_612), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_566), .B(n_67), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_568), .A2(n_206), .B(n_231), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_614), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_592), .B(n_70), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g714 ( .A(n_604), .B(n_183), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_540), .B(n_71), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_597), .B(n_73), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_554), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_563), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_577), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g720 ( .A(n_571), .B(n_184), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_552), .B(n_75), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_553), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_588), .A2(n_77), .B1(n_78), .B2(n_79), .Y(n_723) );
AOI211x1_ASAP7_75t_L g724 ( .A1(n_605), .A2(n_77), .B(n_80), .C(n_81), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_528), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_725) );
OAI21x1_ASAP7_75t_SL g726 ( .A1(n_528), .A2(n_82), .B(n_83), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_528), .B(n_83), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_535), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_528), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_528), .B(n_84), .Y(n_730) );
INVx4_ASAP7_75t_L g731 ( .A(n_535), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_528), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_528), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_528), .B(n_86), .Y(n_734) );
OAI21x1_ASAP7_75t_SL g735 ( .A1(n_528), .A2(n_86), .B(n_87), .Y(n_735) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_537), .A2(n_218), .B(n_230), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_537), .A2(n_216), .B(n_229), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g738 ( .A1(n_528), .A2(n_87), .B(n_88), .C(n_89), .Y(n_738) );
CKINVDCx11_ASAP7_75t_R g739 ( .A(n_535), .Y(n_739) );
NOR4xp25_ASAP7_75t_L g740 ( .A(n_603), .B(n_88), .C(n_89), .D(n_90), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_707), .A2(n_90), .B1(n_91), .B2(n_93), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_699), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_640), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_633), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_654), .B(n_94), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_664), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_728), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_732), .B(n_97), .Y(n_748) );
OR2x6_ASAP7_75t_L g749 ( .A(n_731), .B(n_99), .Y(n_749) );
INVx2_ASAP7_75t_SL g750 ( .A(n_634), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_707), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_733), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_645), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_753) );
NOR4xp25_ASAP7_75t_L g754 ( .A(n_693), .B(n_104), .C(n_105), .D(n_107), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_661), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_688), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_674), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_722), .B(n_222), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_678), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_687), .B(n_689), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_724), .B(n_636), .C(n_703), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_659), .A2(n_662), .B1(n_665), .B2(n_670), .Y(n_762) );
INVx1_ASAP7_75t_SL g763 ( .A(n_674), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_SL g764 ( .A1(n_721), .A2(n_647), .B(n_655), .C(n_736), .Y(n_764) );
INVx8_ASAP7_75t_L g765 ( .A(n_643), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_646), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_724), .B(n_703), .C(n_676), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_625), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g769 ( .A1(n_657), .A2(n_730), .B(n_734), .Y(n_769) );
INVx4_ASAP7_75t_L g770 ( .A(n_643), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_629), .A2(n_656), .B(n_710), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_679), .A2(n_686), .B1(n_639), .B2(n_652), .Y(n_772) );
AO21x2_ASAP7_75t_L g773 ( .A1(n_629), .A2(n_737), .B(n_711), .Y(n_773) );
AO21x2_ASAP7_75t_L g774 ( .A1(n_701), .A2(n_660), .B(n_652), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_693), .B(n_641), .C(n_642), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_L g776 ( .A1(n_716), .A2(n_683), .B(n_649), .C(n_705), .Y(n_776) );
OAI21x1_ASAP7_75t_L g777 ( .A1(n_677), .A2(n_682), .B(n_668), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_628), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_L g779 ( .A1(n_706), .A2(n_684), .B(n_715), .C(n_713), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_623), .A2(n_679), .B1(n_695), .B2(n_626), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_630), .Y(n_781) );
AOI21x1_ASAP7_75t_L g782 ( .A1(n_635), .A2(n_690), .B(n_694), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_637), .B(n_631), .Y(n_783) );
AO21x2_ASAP7_75t_L g784 ( .A1(n_726), .A2(n_735), .B(n_740), .Y(n_784) );
AO31x2_ASAP7_75t_L g785 ( .A1(n_671), .A2(n_653), .A3(n_738), .B(n_692), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_727), .Y(n_786) );
OA21x2_ASAP7_75t_L g787 ( .A1(n_691), .A2(n_720), .B(n_663), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_704), .B(n_719), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_666), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_704), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_680), .A2(n_709), .B1(n_712), .B2(n_667), .Y(n_791) );
OR2x6_ASAP7_75t_L g792 ( .A(n_658), .B(n_651), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_740), .A2(n_720), .B(n_644), .Y(n_793) );
OAI21xp5_ASAP7_75t_L g794 ( .A1(n_723), .A2(n_650), .B(n_725), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_717), .B(n_666), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_697), .A2(n_638), .B(n_681), .Y(n_796) );
NAND3xp33_ASAP7_75t_SL g797 ( .A(n_718), .B(n_714), .C(n_672), .Y(n_797) );
NAND2x1p5_ASAP7_75t_L g798 ( .A(n_648), .B(n_700), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_669), .A2(n_702), .B1(n_696), .B2(n_708), .Y(n_799) );
AO21x2_ASAP7_75t_L g800 ( .A1(n_698), .A2(n_673), .B(n_675), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_698), .B(n_696), .Y(n_801) );
BUFx3_ASAP7_75t_L g802 ( .A(n_739), .Y(n_802) );
NOR4xp25_ASAP7_75t_L g803 ( .A(n_693), .B(n_652), .C(n_683), .D(n_603), .Y(n_803) );
AO22x2_ASAP7_75t_L g804 ( .A1(n_703), .A2(n_477), .B1(n_724), .B2(n_543), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_729), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_739), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_729), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_729), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_739), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_729), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_674), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_685), .A2(n_532), .B(n_537), .Y(n_812) );
OA21x2_ASAP7_75t_L g813 ( .A1(n_622), .A2(n_627), .B(n_619), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_731), .B(n_729), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_728), .B(n_550), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_729), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_699), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_699), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_664), .A2(n_530), .B1(n_608), .B2(n_528), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_622), .A2(n_624), .B(n_632), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_699), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_699), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_664), .A2(n_530), .B1(n_608), .B2(n_528), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_627), .A2(n_619), .B(n_618), .Y(n_824) );
AND2x4_ASAP7_75t_L g825 ( .A(n_731), .B(n_729), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_731), .B(n_729), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_729), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_731), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_664), .A2(n_530), .B1(n_608), .B2(n_528), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_724), .B(n_636), .C(n_703), .Y(n_830) );
AND2x4_ASAP7_75t_L g831 ( .A(n_731), .B(n_729), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_699), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_744), .Y(n_833) );
BUFx3_ASAP7_75t_L g834 ( .A(n_765), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_743), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_757), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_742), .Y(n_837) );
BUFx3_ASAP7_75t_L g838 ( .A(n_765), .Y(n_838) );
INVx3_ASAP7_75t_L g839 ( .A(n_798), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_805), .B(n_807), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_817), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_755), .B(n_756), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_818), .Y(n_843) );
BUFx2_ASAP7_75t_L g844 ( .A(n_828), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_821), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_822), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_814), .B(n_825), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_763), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_832), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g850 ( .A1(n_780), .A2(n_776), .B(n_803), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_780), .A2(n_803), .B(n_775), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_759), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_752), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_825), .B(n_826), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_813), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_808), .Y(n_856) );
INVxp67_ASAP7_75t_L g857 ( .A(n_747), .Y(n_857) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_811), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_804), .A2(n_745), .B1(n_819), .B2(n_829), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_810), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_816), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_827), .Y(n_862) );
OR2x6_ASAP7_75t_L g863 ( .A(n_823), .B(n_829), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_748), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_748), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_820), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_831), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_788), .Y(n_868) );
BUFx2_ASAP7_75t_L g869 ( .A(n_792), .Y(n_869) );
OR2x6_ASAP7_75t_L g870 ( .A(n_749), .B(n_746), .Y(n_870) );
INVx4_ASAP7_75t_L g871 ( .A(n_770), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_746), .Y(n_872) );
BUFx2_ASAP7_75t_L g873 ( .A(n_792), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_777), .Y(n_874) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_772), .A2(n_783), .B1(n_766), .B2(n_768), .C1(n_781), .C2(n_806), .Y(n_875) );
INVx3_ASAP7_75t_L g876 ( .A(n_770), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_772), .A2(n_749), .B1(n_799), .B2(n_762), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_815), .B(n_760), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_800), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_783), .Y(n_880) );
NOR2x1_ASAP7_75t_SL g881 ( .A(n_795), .B(n_797), .Y(n_881) );
AOI211x1_ASAP7_75t_L g882 ( .A1(n_794), .A2(n_767), .B(n_793), .C(n_830), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_809), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_801), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_789), .Y(n_885) );
AND2x4_ASAP7_75t_L g886 ( .A(n_790), .B(n_812), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_758), .B(n_750), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_762), .A2(n_786), .B1(n_778), .B2(n_791), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_753), .B(n_751), .Y(n_889) );
OR2x6_ASAP7_75t_L g890 ( .A(n_795), .B(n_802), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_779), .B(n_794), .Y(n_891) );
OA21x2_ASAP7_75t_L g892 ( .A1(n_793), .A2(n_771), .B(n_824), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_784), .Y(n_893) );
INVx3_ASAP7_75t_L g894 ( .A(n_789), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_784), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_796), .Y(n_896) );
INVx2_ASAP7_75t_SL g897 ( .A(n_871), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_848), .B(n_754), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_884), .B(n_761), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_848), .B(n_830), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_880), .B(n_741), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_851), .B(n_774), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_886), .B(n_774), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_886), .B(n_773), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_886), .B(n_773), .Y(n_905) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_858), .Y(n_906) );
BUFx2_ASAP7_75t_L g907 ( .A(n_863), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_863), .B(n_785), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_855), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_858), .B(n_785), .Y(n_910) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_844), .Y(n_911) );
OR2x2_ASAP7_75t_L g912 ( .A(n_863), .B(n_785), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_878), .B(n_769), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_850), .B(n_769), .Y(n_914) );
BUFx3_ASAP7_75t_L g915 ( .A(n_876), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_879), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_836), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_840), .B(n_787), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_893), .B(n_782), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_895), .B(n_764), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_871), .Y(n_921) );
OR2x2_ASAP7_75t_L g922 ( .A(n_872), .B(n_870), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_868), .B(n_888), .Y(n_923) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_847), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_888), .B(n_833), .Y(n_925) );
BUFx2_ASAP7_75t_L g926 ( .A(n_870), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_891), .B(n_837), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_882), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_877), .B(n_842), .Y(n_929) );
NAND2x1p5_ASAP7_75t_L g930 ( .A(n_876), .B(n_885), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_841), .B(n_843), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_854), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_845), .B(n_846), .Y(n_933) );
OR2x2_ASAP7_75t_L g934 ( .A(n_864), .B(n_865), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_849), .B(n_852), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_856), .B(n_860), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_909), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_916), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_927), .B(n_875), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_931), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_931), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_908), .B(n_892), .Y(n_942) );
INVxp67_ASAP7_75t_SL g943 ( .A(n_917), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_922), .B(n_892), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_908), .B(n_892), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_933), .B(n_835), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_899), .B(n_859), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_935), .B(n_925), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_899), .B(n_859), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_934), .Y(n_950) );
BUFx6f_ASAP7_75t_L g951 ( .A(n_919), .Y(n_951) );
NAND2x1p5_ASAP7_75t_L g952 ( .A(n_897), .B(n_834), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_900), .B(n_857), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_920), .B(n_896), .Y(n_954) );
BUFx2_ASAP7_75t_L g955 ( .A(n_915), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_920), .B(n_896), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_936), .B(n_853), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_912), .B(n_874), .Y(n_958) );
INVx4_ASAP7_75t_L g959 ( .A(n_915), .Y(n_959) );
BUFx2_ASAP7_75t_L g960 ( .A(n_915), .Y(n_960) );
NAND2x1p5_ASAP7_75t_SL g961 ( .A(n_897), .B(n_889), .Y(n_961) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_911), .Y(n_962) );
AND2x4_ASAP7_75t_L g963 ( .A(n_926), .B(n_881), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_918), .B(n_866), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_923), .B(n_862), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_921), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_921), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_938), .Y(n_968) );
INVx3_ASAP7_75t_L g969 ( .A(n_951), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_940), .B(n_928), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_941), .B(n_928), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_938), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_942), .B(n_904), .Y(n_973) );
INVx2_ASAP7_75t_SL g974 ( .A(n_966), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_945), .B(n_905), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_945), .B(n_905), .Y(n_976) );
AND2x4_ASAP7_75t_L g977 ( .A(n_954), .B(n_903), .Y(n_977) );
OR2x2_ASAP7_75t_L g978 ( .A(n_948), .B(n_910), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_937), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_964), .B(n_902), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_954), .B(n_902), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_953), .B(n_898), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_956), .B(n_907), .Y(n_983) );
INVxp67_ASAP7_75t_L g984 ( .A(n_967), .Y(n_984) );
AND2x4_ASAP7_75t_L g985 ( .A(n_951), .B(n_919), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_950), .B(n_906), .Y(n_986) );
INVx3_ASAP7_75t_L g987 ( .A(n_951), .Y(n_987) );
INVxp33_ASAP7_75t_L g988 ( .A(n_952), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_958), .B(n_914), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_943), .Y(n_990) );
AOI21xp33_ASAP7_75t_SL g991 ( .A1(n_988), .A2(n_961), .B(n_952), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_979), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_989), .B(n_947), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_973), .B(n_944), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_973), .B(n_944), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_968), .Y(n_996) );
AND2x4_ASAP7_75t_L g997 ( .A(n_985), .B(n_951), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_975), .B(n_949), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_972), .Y(n_999) );
NAND2xp5_ASAP7_75t_SL g1000 ( .A(n_974), .B(n_959), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_975), .B(n_951), .Y(n_1001) );
INVxp67_ASAP7_75t_L g1002 ( .A(n_990), .Y(n_1002) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_982), .B(n_962), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_982), .B(n_965), .Y(n_1004) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_985), .B(n_955), .Y(n_1005) );
NAND2x1p5_ASAP7_75t_L g1006 ( .A(n_986), .B(n_959), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_976), .B(n_919), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_984), .Y(n_1008) );
INVx2_ASAP7_75t_L g1009 ( .A(n_992), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_1006), .A2(n_939), .B1(n_978), .B2(n_963), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_1002), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1003), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1003), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_994), .B(n_980), .Y(n_1014) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_1000), .B(n_983), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1016 ( .A(n_1006), .Y(n_1016) );
NAND3xp33_ASAP7_75t_L g1017 ( .A(n_1008), .B(n_971), .C(n_970), .Y(n_1017) );
NAND3x2_ASAP7_75t_L g1018 ( .A(n_1004), .B(n_873), .C(n_869), .Y(n_1018) );
INVx1_ASAP7_75t_SL g1019 ( .A(n_1015), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_1016), .A2(n_991), .B1(n_1004), .B2(n_993), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_1010), .A2(n_1007), .B1(n_1001), .B2(n_1005), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_1018), .A2(n_1005), .B1(n_998), .B2(n_995), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1011), .B(n_981), .Y(n_1023) );
XNOR2x1_ASAP7_75t_L g1024 ( .A(n_1019), .B(n_883), .Y(n_1024) );
AOI211x1_ASAP7_75t_L g1025 ( .A1(n_1020), .A2(n_1013), .B(n_1012), .C(n_1017), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1021), .B(n_1014), .Y(n_1026) );
OAI322xp33_ASAP7_75t_L g1027 ( .A1(n_1022), .A2(n_946), .A3(n_957), .B1(n_986), .B2(n_929), .C1(n_934), .C2(n_913), .Y(n_1027) );
NAND2xp5_ASAP7_75t_SL g1028 ( .A(n_1023), .B(n_1009), .Y(n_1028) );
NAND3xp33_ASAP7_75t_L g1029 ( .A(n_1025), .B(n_883), .C(n_887), .Y(n_1029) );
NOR3x1_ASAP7_75t_SL g1030 ( .A(n_1024), .B(n_890), .C(n_924), .Y(n_1030) );
NOR4xp75_ASAP7_75t_L g1031 ( .A(n_1030), .B(n_1027), .C(n_1028), .D(n_1026), .Y(n_1031) );
NOR2x1_ASAP7_75t_L g1032 ( .A(n_1029), .B(n_838), .Y(n_1032) );
INVx1_ASAP7_75t_SL g1033 ( .A(n_1032), .Y(n_1033) );
NAND2xp5_ASAP7_75t_SL g1034 ( .A(n_1033), .B(n_1031), .Y(n_1034) );
OAI22x1_ASAP7_75t_SL g1035 ( .A1(n_1034), .A2(n_867), .B1(n_839), .B2(n_885), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_1035), .B(n_932), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_1036), .A2(n_997), .B1(n_987), .B2(n_969), .Y(n_1037) );
OAI21xp33_ASAP7_75t_L g1038 ( .A1(n_1037), .A2(n_901), .B(n_997), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_1038), .A2(n_861), .B1(n_894), .B2(n_999), .C(n_996), .Y(n_1039) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_1039), .A2(n_930), .B1(n_960), .B2(n_987), .C(n_969), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1040), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_1041), .A2(n_985), .B1(n_977), .B2(n_987), .Y(n_1042) );
endmodule