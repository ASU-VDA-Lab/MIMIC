module real_aes_6825_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_0), .Y(n_161) );
INVx1_ASAP7_75t_L g276 ( .A(n_1), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g124 ( .A1(n_2), .A2(n_19), .B1(n_125), .B2(n_133), .Y(n_124) );
AOI21xp33_ASAP7_75t_L g245 ( .A1(n_3), .A2(n_220), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g203 ( .A(n_4), .Y(n_203) );
AND2x6_ASAP7_75t_L g225 ( .A(n_4), .B(n_201), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_4), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_5), .A2(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g252 ( .A(n_6), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_7), .B(n_318), .Y(n_317) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_8), .A2(n_28), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g218 ( .A(n_9), .Y(n_218) );
INVx1_ASAP7_75t_L g332 ( .A(n_10), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g115 ( .A1(n_11), .A2(n_51), .B1(n_116), .B2(n_120), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_12), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_13), .A2(n_81), .B1(n_82), .B2(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_13), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_14), .A2(n_34), .B1(n_178), .B2(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g179 ( .A(n_14), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_14), .B(n_233), .Y(n_305) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_15), .A2(n_29), .B1(n_89), .B2(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_16), .B(n_220), .Y(n_288) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_17), .A2(n_58), .B1(n_182), .B2(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_17), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_18), .B(n_241), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_20), .A2(n_330), .B(n_331), .C(n_333), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g139 ( .A1(n_21), .A2(n_24), .B1(n_140), .B2(n_142), .Y(n_139) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_22), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_23), .B(n_250), .Y(n_278) );
INVx1_ASAP7_75t_L g265 ( .A(n_25), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g147 ( .A1(n_26), .A2(n_32), .B1(n_148), .B2(n_151), .Y(n_147) );
INVx2_ASAP7_75t_L g223 ( .A(n_27), .Y(n_223) );
OAI221xp5_ASAP7_75t_L g194 ( .A1(n_29), .A2(n_43), .B1(n_52), .B2(n_195), .C(n_196), .Y(n_194) );
INVxp67_ASAP7_75t_L g197 ( .A(n_29), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_30), .A2(n_81), .B1(n_82), .B2(n_173), .Y(n_80) );
INVx1_ASAP7_75t_L g173 ( .A(n_30), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_31), .A2(n_225), .B(n_228), .C(n_290), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_33), .Y(n_168) );
INVx1_ASAP7_75t_L g178 ( .A(n_34), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_35), .B(n_250), .Y(n_304) );
AOI211xp5_ASAP7_75t_L g155 ( .A1(n_36), .A2(n_156), .B(n_158), .C(n_167), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_37), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_38), .B(n_220), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_39), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_40), .A2(n_228), .B1(n_260), .B2(n_262), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_41), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g273 ( .A(n_42), .Y(n_273) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_43), .A2(n_60), .B1(n_89), .B2(n_93), .Y(n_96) );
INVxp67_ASAP7_75t_L g198 ( .A(n_43), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_44), .A2(n_237), .B(n_249), .C(n_251), .Y(n_248) );
AOI22xp5_ASAP7_75t_SL g536 ( .A1(n_44), .A2(n_81), .B1(n_82), .B2(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_44), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_45), .Y(n_308) );
INVx1_ASAP7_75t_L g247 ( .A(n_46), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_47), .Y(n_108) );
INVx1_ASAP7_75t_L g201 ( .A(n_48), .Y(n_201) );
INVx1_ASAP7_75t_L g217 ( .A(n_49), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_50), .Y(n_195) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_52), .A2(n_66), .B1(n_89), .B2(n_90), .Y(n_98) );
A2O1A1Ixp33_ASAP7_75t_SL g232 ( .A1(n_53), .A2(n_233), .B(n_234), .C(n_237), .Y(n_232) );
INVxp67_ASAP7_75t_L g235 ( .A(n_54), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_55), .Y(n_269) );
INVx1_ASAP7_75t_L g301 ( .A(n_56), .Y(n_301) );
INVx1_ASAP7_75t_L g190 ( .A(n_57), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_58), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_59), .A2(n_225), .B(n_228), .C(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_61), .B(n_277), .Y(n_291) );
INVx2_ASAP7_75t_L g215 ( .A(n_62), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_63), .B(n_233), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_64), .A2(n_225), .B(n_228), .C(n_275), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_65), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_65), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_67), .B(n_254), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_68), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_69), .A2(n_225), .B(n_228), .C(n_315), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_70), .Y(n_322) );
INVx1_ASAP7_75t_L g231 ( .A(n_71), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_72), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_73), .B(n_277), .Y(n_316) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_75), .B(n_213), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_76), .A2(n_220), .B(n_226), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_77), .Y(n_113) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_191), .B1(n_204), .B2(n_527), .C(n_535), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_174), .Y(n_79) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND3x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_138), .C(n_155), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_114), .Y(n_83) );
OAI222xp33_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_99), .B1(n_100), .B2(n_108), .C1(n_109), .C2(n_113), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x6_ASAP7_75t_L g86 ( .A(n_87), .B(n_94), .Y(n_86) );
AND2x4_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
AND2x2_ASAP7_75t_L g107 ( .A(n_88), .B(n_96), .Y(n_107) );
INVx2_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
INVx2_ASAP7_75t_L g106 ( .A(n_92), .Y(n_106) );
INVx1_ASAP7_75t_L g119 ( .A(n_92), .Y(n_119) );
OR2x2_ASAP7_75t_L g131 ( .A(n_92), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g137 ( .A(n_92), .B(n_132), .Y(n_137) );
AND2x4_ASAP7_75t_L g141 ( .A(n_94), .B(n_137), .Y(n_141) );
AND2x2_ASAP7_75t_L g157 ( .A(n_94), .B(n_146), .Y(n_157) );
AND2x6_ASAP7_75t_L g172 ( .A(n_94), .B(n_130), .Y(n_172) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_97), .Y(n_94) );
AND2x2_ASAP7_75t_L g129 ( .A(n_95), .B(n_98), .Y(n_129) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g145 ( .A(n_96), .B(n_123), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_96), .B(n_98), .Y(n_154) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx1_ASAP7_75t_L g105 ( .A(n_98), .Y(n_105) );
INVx1_ASAP7_75t_L g123 ( .A(n_98), .Y(n_123) );
INVx2_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g112 ( .A(n_105), .Y(n_112) );
AND2x2_ASAP7_75t_L g146 ( .A(n_106), .B(n_132), .Y(n_146) );
AND2x4_ASAP7_75t_L g111 ( .A(n_107), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g117 ( .A(n_107), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_124), .Y(n_114) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OR2x6_ASAP7_75t_L g165 ( .A(n_119), .B(n_154), .Y(n_165) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x6_ASAP7_75t_L g136 ( .A(n_129), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g150 ( .A(n_129), .B(n_146), .Y(n_150) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx4f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_137), .B(n_145), .Y(n_160) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_147), .Y(n_138) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g152 ( .A(n_146), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_159), .A2(n_161), .B1(n_162), .B2(n_166), .Y(n_158) );
BUFx2_ASAP7_75t_R g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx6_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx11_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B1(n_185), .B2(n_186), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B1(n_181), .B2(n_184), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_177), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g262 ( .A1(n_178), .A2(n_263), .B1(n_264), .B2(n_265), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
AND3x1_ASAP7_75t_SL g193 ( .A(n_194), .B(n_199), .C(n_202), .Y(n_193) );
INVxp67_ASAP7_75t_L g541 ( .A(n_194), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx1_ASAP7_75t_SL g543 ( .A(n_199), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_199), .A2(n_546), .B(n_548), .Y(n_545) );
INVx1_ASAP7_75t_L g554 ( .A(n_199), .Y(n_554) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_200), .B(n_203), .Y(n_548) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_SL g553 ( .A(n_202), .B(n_554), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND4x1_ASAP7_75t_L g205 ( .A(n_206), .B(n_445), .C(n_492), .D(n_512), .Y(n_205) );
NOR3xp33_ASAP7_75t_SL g206 ( .A(n_207), .B(n_375), .C(n_400), .Y(n_206) );
OAI211xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_283), .B(n_335), .C(n_365), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_255), .Y(n_209) );
INVx3_ASAP7_75t_SL g417 ( .A(n_210), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_210), .B(n_348), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_210), .B(n_270), .Y(n_498) );
AND2x2_ASAP7_75t_L g521 ( .A(n_210), .B(n_387), .Y(n_521) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_243), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g339 ( .A(n_212), .B(n_244), .Y(n_339) );
INVx3_ASAP7_75t_L g352 ( .A(n_212), .Y(n_352) );
AND2x2_ASAP7_75t_L g357 ( .A(n_212), .B(n_243), .Y(n_357) );
OR2x2_ASAP7_75t_L g408 ( .A(n_212), .B(n_349), .Y(n_408) );
BUFx2_ASAP7_75t_L g428 ( .A(n_212), .Y(n_428) );
AND2x2_ASAP7_75t_L g438 ( .A(n_212), .B(n_349), .Y(n_438) );
AND2x2_ASAP7_75t_L g444 ( .A(n_212), .B(n_256), .Y(n_444) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_240), .Y(n_212) );
INVx4_ASAP7_75t_L g242 ( .A(n_213), .Y(n_242) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g257 ( .A(n_214), .Y(n_257) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_215), .B(n_216), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
BUFx2_ASAP7_75t_L g326 ( .A(n_220), .Y(n_326) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g267 ( .A(n_221), .B(n_225), .Y(n_267) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g534 ( .A(n_222), .Y(n_534) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g229 ( .A(n_223), .Y(n_229) );
INVx1_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
INVx1_ASAP7_75t_L g230 ( .A(n_224), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_224), .Y(n_233) );
INVx3_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_224), .Y(n_250) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_224), .Y(n_263) );
INVx4_ASAP7_75t_SL g239 ( .A(n_225), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_231), .B(n_232), .C(n_239), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_227), .A2(n_239), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_227), .A2(n_239), .B(n_328), .C(n_329), .Y(n_327) );
INVx5_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_229), .Y(n_238) );
BUFx3_ASAP7_75t_L g295 ( .A(n_229), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_236), .B(n_252), .Y(n_251) );
INVx5_ASAP7_75t_L g277 ( .A(n_236), .Y(n_277) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_238), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g258 ( .A1(n_239), .A2(n_259), .B1(n_266), .B2(n_267), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_239), .B(n_533), .Y(n_532) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_241), .A2(n_245), .B(n_253), .Y(n_244) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_242), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_244), .B(n_349), .Y(n_363) );
INVx2_ASAP7_75t_L g373 ( .A(n_244), .Y(n_373) );
AND2x2_ASAP7_75t_L g386 ( .A(n_244), .B(n_352), .Y(n_386) );
OR2x2_ASAP7_75t_L g397 ( .A(n_244), .B(n_349), .Y(n_397) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_244), .B(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g455 ( .A(n_244), .Y(n_455) );
AND2x2_ASAP7_75t_L g501 ( .A(n_244), .B(n_256), .Y(n_501) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g318 ( .A(n_250), .Y(n_318) );
OAI322xp33_ASAP7_75t_L g535 ( .A1(n_252), .A2(n_536), .A3(n_538), .B1(n_542), .B2(n_544), .C1(n_549), .C2(n_551), .Y(n_535) );
INVx1_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
INVx2_ASAP7_75t_L g312 ( .A(n_254), .Y(n_312) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_254), .A2(n_325), .B(n_334), .Y(n_324) );
INVx3_ASAP7_75t_SL g374 ( .A(n_255), .Y(n_374) );
OR2x2_ASAP7_75t_L g427 ( .A(n_255), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_270), .Y(n_255) );
INVx3_ASAP7_75t_L g349 ( .A(n_256), .Y(n_349) );
AND2x2_ASAP7_75t_L g416 ( .A(n_256), .B(n_271), .Y(n_416) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_256), .Y(n_484) );
AOI33xp33_ASAP7_75t_L g488 ( .A1(n_256), .A2(n_417), .A3(n_424), .B1(n_433), .B2(n_489), .B3(n_490), .Y(n_488) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_268), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_257), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_257), .A2(n_272), .B(n_280), .Y(n_271) );
INVx2_ASAP7_75t_L g296 ( .A(n_257), .Y(n_296) );
INVx2_ASAP7_75t_L g279 ( .A(n_260), .Y(n_279) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g264 ( .A(n_263), .Y(n_264) );
INVx4_ASAP7_75t_L g330 ( .A(n_263), .Y(n_330) );
INVx2_ASAP7_75t_L g531 ( .A(n_264), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_267), .A2(n_273), .B(n_274), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_270), .B(n_352), .Y(n_351) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_270), .B(n_412), .C(n_414), .Y(n_411) );
AND2x2_ASAP7_75t_L g437 ( .A(n_270), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_270), .B(n_444), .Y(n_447) );
AND2x2_ASAP7_75t_L g500 ( .A(n_270), .B(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g356 ( .A(n_271), .Y(n_356) );
OR2x2_ASAP7_75t_L g450 ( .A(n_271), .B(n_349), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .B(n_278), .C(n_279), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_282), .B(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_282), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_309), .Y(n_283) );
AOI32xp33_ASAP7_75t_L g401 ( .A1(n_284), .A2(n_402), .A3(n_404), .B1(n_406), .B2(n_409), .Y(n_401) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_284), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g504 ( .A(n_284), .Y(n_504) );
INVx4_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g436 ( .A(n_285), .B(n_420), .Y(n_436) );
AND2x2_ASAP7_75t_L g456 ( .A(n_285), .B(n_382), .Y(n_456) );
AND2x2_ASAP7_75t_L g524 ( .A(n_285), .B(n_442), .Y(n_524) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_299), .Y(n_285) );
INVx3_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
AND2x2_ASAP7_75t_L g359 ( .A(n_286), .B(n_343), .Y(n_359) );
OR2x2_ASAP7_75t_L g364 ( .A(n_286), .B(n_342), .Y(n_364) );
INVx1_ASAP7_75t_L g371 ( .A(n_286), .Y(n_371) );
AND2x2_ASAP7_75t_L g379 ( .A(n_286), .B(n_353), .Y(n_379) );
AND2x2_ASAP7_75t_L g381 ( .A(n_286), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_286), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g434 ( .A(n_286), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_286), .B(n_519), .Y(n_518) );
OR2x6_ASAP7_75t_L g286 ( .A(n_287), .B(n_297), .Y(n_286) );
AOI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_289), .B(n_296), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_293), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_293), .A2(n_304), .B(n_305), .Y(n_303) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx1_ASAP7_75t_L g306 ( .A(n_296), .Y(n_306) );
INVx2_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
AND2x2_ASAP7_75t_L g389 ( .A(n_299), .B(n_310), .Y(n_389) );
AND2x2_ASAP7_75t_L g399 ( .A(n_299), .B(n_324), .Y(n_399) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B(n_307), .Y(n_299) );
INVx2_ASAP7_75t_L g519 ( .A(n_309), .Y(n_519) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_323), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_310), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g360 ( .A(n_310), .Y(n_360) );
AND2x2_ASAP7_75t_L g404 ( .A(n_310), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g420 ( .A(n_310), .B(n_383), .Y(n_420) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
AND2x2_ASAP7_75t_L g382 ( .A(n_311), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g433 ( .A(n_311), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_311), .B(n_343), .Y(n_465) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B(n_321), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_320), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_319), .Y(n_315) );
AND2x2_ASAP7_75t_L g344 ( .A(n_323), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g405 ( .A(n_323), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_323), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g442 ( .A(n_323), .Y(n_442) );
INVx1_ASAP7_75t_L g475 ( .A(n_323), .Y(n_475) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g353 ( .A(n_324), .B(n_343), .Y(n_353) );
INVx1_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_330), .B(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B1(n_346), .B2(n_353), .C(n_354), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_337), .B(n_357), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_337), .B(n_420), .Y(n_497) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_339), .B(n_387), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_339), .B(n_348), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_339), .B(n_362), .Y(n_491) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g413 ( .A(n_343), .Y(n_413) );
AND2x2_ASAP7_75t_L g388 ( .A(n_344), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g466 ( .A(n_344), .Y(n_466) );
AND2x2_ASAP7_75t_L g398 ( .A(n_345), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_345), .B(n_368), .Y(n_414) );
AND2x2_ASAP7_75t_L g478 ( .A(n_345), .B(n_404), .Y(n_478) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g387 ( .A(n_349), .B(n_356), .Y(n_387) );
AND2x2_ASAP7_75t_L g483 ( .A(n_350), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_352), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_353), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_353), .B(n_360), .Y(n_448) );
AND2x2_ASAP7_75t_L g468 ( .A(n_353), .B(n_368), .Y(n_468) );
AND2x2_ASAP7_75t_L g489 ( .A(n_353), .B(n_433), .Y(n_489) );
OAI32xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .A3(n_360), .B1(n_361), .B2(n_364), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_SL g362 ( .A(n_356), .Y(n_362) );
NAND2x1_ASAP7_75t_L g403 ( .A(n_356), .B(n_386), .Y(n_403) );
OR2x2_ASAP7_75t_L g407 ( .A(n_356), .B(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_356), .B(n_455), .Y(n_508) );
INVx1_ASAP7_75t_L g376 ( .A(n_357), .Y(n_376) );
OAI221xp5_ASAP7_75t_SL g494 ( .A1(n_358), .A2(n_449), .B1(n_495), .B2(n_498), .C(n_499), .Y(n_494) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g366 ( .A(n_359), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g409 ( .A(n_359), .B(n_382), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_359), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g487 ( .A(n_359), .B(n_420), .Y(n_487) );
INVxp67_ASAP7_75t_L g423 ( .A(n_360), .Y(n_423) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g493 ( .A(n_362), .B(n_480), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_362), .B(n_443), .Y(n_516) );
INVx1_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_364), .B(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g509 ( .A(n_364), .B(n_510), .Y(n_509) );
OAI21xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_369), .B(n_372), .Y(n_365) );
AND2x2_ASAP7_75t_L g378 ( .A(n_367), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g462 ( .A(n_371), .B(n_382), .Y(n_462) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g480 ( .A(n_373), .B(n_438), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_373), .B(n_437), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_374), .B(n_386), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_380), .C(n_390), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_376), .A2(n_411), .B1(n_415), .B2(n_418), .C(n_421), .Y(n_410) );
AOI31xp33_ASAP7_75t_L g505 ( .A1(n_376), .A2(n_506), .A3(n_507), .B(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B1(n_386), .B2(n_388), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g506 ( .A(n_386), .Y(n_506) );
INVx1_ASAP7_75t_L g469 ( .A(n_387), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_389), .A2(n_513), .B(n_515), .C(n_517), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_394), .B2(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_395), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_SL g485 ( .A1(n_397), .A2(n_431), .B1(n_450), .B2(n_486), .C(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g481 ( .A(n_398), .Y(n_481) );
INVx1_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_410), .C(n_425), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g451 ( .A1(n_402), .A2(n_452), .B(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_404), .B(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_L g511 ( .A(n_405), .Y(n_511) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g449 ( .A(n_412), .B(n_432), .Y(n_449) );
INVx1_ASAP7_75t_L g424 ( .A(n_413), .Y(n_424) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_416), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_416), .B(n_454), .Y(n_453) );
NOR4xp25_ASAP7_75t_L g421 ( .A(n_417), .B(n_422), .C(n_423), .D(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B1(n_436), .B2(n_437), .C1(n_439), .C2(n_443), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g523 ( .A(n_427), .Y(n_523) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_439), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g499 ( .A1(n_444), .A2(n_500), .B(n_502), .Y(n_499) );
NOR4xp25_ASAP7_75t_L g445 ( .A(n_446), .B(n_457), .C(n_470), .D(n_485), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_448), .B1(n_449), .B2(n_450), .C(n_451), .Y(n_446) );
INVx1_ASAP7_75t_L g526 ( .A(n_447), .Y(n_526) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_454), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OAI222xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B1(n_463), .B2(n_464), .C1(n_467), .C2(n_469), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g492 ( .A1(n_462), .A2(n_493), .B(n_494), .C(n_505), .Y(n_492) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
OAI222xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_476), .B1(n_477), .B2(n_479), .C1(n_481), .C2(n_482), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_487), .A2(n_490), .B1(n_523), .B2(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI211xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_520), .B(n_522), .C(n_525), .Y(n_517) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g547 ( .A(n_530), .Y(n_547) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_533), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
endmodule