module fake_jpeg_26655_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_6),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_22),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_62),
.B1(n_21),
.B2(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_22),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_29),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_19),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_36),
.C(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_62),
.B1(n_23),
.B2(n_16),
.Y(n_102)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_75),
.Y(n_99)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_41),
.B1(n_45),
.B2(n_64),
.Y(n_90)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_65),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_41),
.B(n_33),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_40),
.B(n_31),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_50),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_48),
.B1(n_60),
.B2(n_81),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_94),
.C(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_100),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_57),
.C(n_44),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_63),
.B(n_54),
.C(n_49),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_42),
.B(n_66),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_57),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_40),
.B1(n_33),
.B2(n_27),
.C(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_81),
.B1(n_48),
.B2(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_47),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_42),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_47),
.B1(n_53),
.B2(n_49),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_116),
.B1(n_103),
.B2(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_119),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_122),
.B1(n_20),
.B2(n_26),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_85),
.C(n_75),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_69),
.B1(n_68),
.B2(n_42),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_89),
.B1(n_86),
.B2(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_100),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_91),
.B(n_87),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_145),
.B1(n_146),
.B2(n_111),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_148),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_94),
.B1(n_101),
.B2(n_98),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_42),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_122),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_106),
.B(n_16),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_74),
.B1(n_95),
.B2(n_16),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_116),
.B(n_106),
.C(n_108),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_95),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_145),
.B1(n_138),
.B2(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_114),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_172),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_165),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_131),
.B(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_126),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_124),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_109),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_128),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_115),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_24),
.B(n_23),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_119),
.C(n_121),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_142),
.C(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_3),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_138),
.B1(n_149),
.B2(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_171),
.B1(n_21),
.B2(n_42),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_140),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_189),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_164),
.B1(n_163),
.B2(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_180),
.C(n_178),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_187),
.B(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_136),
.B(n_143),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_136),
.B(n_144),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_130),
.Y(n_189)
);

OAI321xp33_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_155),
.A3(n_156),
.B1(n_24),
.B2(n_21),
.C(n_171),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_1),
.B(n_2),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_24),
.B(n_23),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_163),
.B(n_25),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_194),
.B(n_25),
.CI(n_36),
.CON(n_203),
.SN(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_199),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_184),
.B1(n_188),
.B2(n_179),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_154),
.A3(n_157),
.B1(n_155),
.B2(n_156),
.C1(n_175),
.C2(n_164),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_3),
.C(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_192),
.B1(n_182),
.B2(n_188),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_207),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_36),
.C(n_25),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_193),
.C(n_4),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_2),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_209),
.B(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_224)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_217),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_189),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_219),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_194),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_222),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_221),
.B(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_224),
.A2(n_204),
.B1(n_203),
.B2(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_204),
.B(n_203),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_230),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_219),
.A2(n_212),
.B(n_217),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_5),
.B(n_6),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

OAI21x1_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_211),
.B(n_220),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_239),
.B1(n_5),
.B2(n_10),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_235),
.B(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_237),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_245),
.A3(n_242),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_237),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_234),
.C(n_226),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_5),
.Y(n_250)
);

AOI321xp33_ASAP7_75t_SL g252 ( 
.A1(n_250),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_251),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_14),
.Y(n_254)
);


endmodule