module fake_jpeg_2768_n_652 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_652);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_652;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_60),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_62),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_82),
.Y(n_138)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_19),
.B(n_2),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_67),
.B(n_90),
.Y(n_225)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_70),
.B(n_122),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_78),
.Y(n_189)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_83),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_86),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_34),
.Y(n_87)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_29),
.B(n_0),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_22),
.B(n_0),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_96),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_112),
.Y(n_146)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_98),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_49),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_49),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_119),
.Y(n_152)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

BUFx16f_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_51),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_39),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_127),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_0),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_130),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_117),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_27),
.B(n_2),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_133),
.B(n_136),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_41),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_27),
.B1(n_32),
.B2(n_53),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_137),
.A2(n_180),
.B1(n_187),
.B2(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_64),
.B(n_42),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_143),
.B(n_145),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_42),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_48),
.B1(n_32),
.B2(n_53),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_153),
.A2(n_163),
.B1(n_166),
.B2(n_172),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_61),
.A2(n_48),
.B1(n_38),
.B2(n_52),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_155),
.A2(n_170),
.B1(n_194),
.B2(n_198),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_111),
.A2(n_52),
.B1(n_47),
.B2(n_40),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_81),
.A2(n_47),
.B1(n_40),
.B2(n_38),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_66),
.A2(n_57),
.B1(n_44),
.B2(n_56),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_87),
.A2(n_57),
.B1(n_44),
.B2(n_5),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_2),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_177),
.B(n_190),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_73),
.B(n_2),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_179),
.B(n_181),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_120),
.A2(n_57),
.B1(n_5),
.B2(n_6),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_70),
.B(n_3),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_78),
.A2(n_57),
.B1(n_6),
.B2(n_7),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_182),
.A2(n_188),
.B(n_224),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_71),
.A2(n_57),
.B1(n_7),
.B2(n_8),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_101),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_62),
.B(n_8),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_84),
.B(n_10),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_192),
.B(n_193),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_10),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_72),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_74),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_75),
.B(n_11),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g280 ( 
.A(n_199),
.B(n_213),
.C(n_221),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_83),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_201),
.A2(n_188),
.B(n_224),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_101),
.B(n_11),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_208),
.B(n_227),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_85),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_215),
.A2(n_220),
.B1(n_201),
.B2(n_170),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_89),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_91),
.A2(n_110),
.B1(n_93),
.B2(n_95),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_99),
.A2(n_123),
.B1(n_122),
.B2(n_127),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_222),
.A2(n_195),
.B1(n_200),
.B2(n_211),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_122),
.A2(n_45),
.B1(n_114),
.B2(n_82),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_129),
.B(n_80),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_94),
.B(n_65),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_228),
.B(n_223),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_140),
.B(n_139),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_230),
.B(n_250),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_231),
.Y(n_331)
);

AO22x1_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_226),
.B1(n_178),
.B2(n_174),
.Y(n_232)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

FAx1_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_138),
.CI(n_186),
.CON(n_235),
.SN(n_235)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_236),
.Y(n_333)
);

OR2x4_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_226),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_238),
.A2(n_262),
.B(n_272),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_144),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_144),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_160),
.A2(n_167),
.B(n_206),
.C(n_162),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_247),
.B(n_260),
.Y(n_326)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_134),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_147),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_176),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_252),
.A2(n_308),
.B1(n_311),
.B2(n_241),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_173),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_255),
.B(n_256),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_146),
.B(n_152),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_258),
.Y(n_332)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_142),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_259),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_261),
.B(n_270),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_166),
.A2(n_153),
.B(n_163),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_175),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_263),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_148),
.B(n_132),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_276),
.Y(n_321)
);

AO22x2_ASAP7_75t_L g265 ( 
.A1(n_172),
.A2(n_182),
.B1(n_210),
.B2(n_159),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_265),
.B(n_289),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_205),
.A2(n_203),
.B(n_212),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_267),
.B(n_273),
.Y(n_334)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_196),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

NAND2xp67_ASAP7_75t_SL g272 ( 
.A(n_203),
.B(n_212),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_197),
.B(n_171),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_275),
.B(n_278),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_155),
.B(n_215),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_142),
.B(n_171),
.C(n_184),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_280),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_197),
.B(n_184),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_213),
.B(n_218),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_149),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_159),
.B(n_214),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_279),
.C(n_260),
.Y(n_325)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_183),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_285),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_219),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_161),
.B(n_204),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_302),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_294),
.Y(n_348)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_135),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_210),
.Y(n_291)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_157),
.Y(n_294)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_175),
.Y(n_295)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_189),
.A2(n_169),
.B(n_154),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_279),
.B(n_264),
.Y(n_354)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_134),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_299),
.B(n_301),
.Y(n_360)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_154),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_303),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_169),
.B(n_189),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_185),
.B(n_202),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_191),
.B(n_204),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_304),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_195),
.B(n_200),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_305),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_135),
.B(n_191),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_306),
.Y(n_365)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_202),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_309),
.B1(n_303),
.B2(n_257),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_221),
.B(n_211),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_223),
.A2(n_225),
.B(n_138),
.C(n_143),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_220),
.A2(n_177),
.B1(n_170),
.B2(n_199),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_138),
.B(n_181),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_323),
.A2(n_328),
.B1(n_367),
.B2(n_303),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_325),
.B(n_269),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_363),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_276),
.A2(n_268),
.B1(n_262),
.B2(n_287),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_251),
.A2(n_238),
.B1(n_241),
.B2(n_252),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_362),
.B1(n_265),
.B2(n_293),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_255),
.C(n_235),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_355),
.C(n_247),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_237),
.A2(n_303),
.B1(n_235),
.B2(n_311),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_353),
.A2(n_363),
.B1(n_307),
.B2(n_286),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_354),
.A2(n_272),
.B(n_243),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_237),
.B(n_244),
.C(n_274),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_268),
.A2(n_232),
.B1(n_308),
.B2(n_287),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_232),
.A2(n_288),
.B1(n_302),
.B2(n_265),
.Y(n_367)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_368),
.B(n_346),
.Y(n_429)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_364),
.Y(n_370)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_266),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_373),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_372),
.A2(n_381),
.B1(n_394),
.B2(n_406),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_229),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_282),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_374),
.B(n_385),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_376),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_312),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_297),
.B(n_265),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_378),
.A2(n_395),
.B(n_403),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_354),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_397),
.Y(n_427)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_380),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_382),
.A2(n_384),
.B(n_389),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_337),
.C(n_317),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_387),
.C(n_401),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_282),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_358),
.B(n_256),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_388),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_233),
.C(n_234),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_275),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_292),
.B(n_261),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_240),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_390),
.B(n_393),
.Y(n_445)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_391),
.Y(n_417)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_355),
.C(n_334),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_392),
.B(n_413),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_298),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_323),
.A2(n_296),
.B1(n_281),
.B2(n_283),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_357),
.A2(n_300),
.B(n_245),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_291),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_407),
.Y(n_446)
);

AO21x1_ASAP7_75t_L g400 ( 
.A1(n_313),
.A2(n_334),
.B(n_362),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_345),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_320),
.B(n_271),
.C(n_239),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_412),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_249),
.B(n_259),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_290),
.B(n_248),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g454 ( 
.A1(n_405),
.A2(n_319),
.B(n_349),
.C(n_315),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_328),
.A2(n_254),
.B1(n_295),
.B2(n_231),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_242),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_367),
.A2(n_246),
.B(n_257),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_315),
.B(n_322),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_246),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_410),
.B(n_411),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_236),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_313),
.B(n_253),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_329),
.B(n_258),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_345),
.A2(n_263),
.B1(n_342),
.B2(n_325),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_402),
.B1(n_397),
.B2(n_379),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_360),
.B(n_345),
.C(n_351),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_352),
.C(n_351),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_393),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_424),
.B(n_386),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_428),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_444),
.C(n_455),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_372),
.A2(n_346),
.B1(n_318),
.B2(n_338),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_430),
.A2(n_431),
.B1(n_432),
.B2(n_447),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_381),
.A2(n_338),
.B1(n_359),
.B2(n_341),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_378),
.A2(n_359),
.B1(n_341),
.B2(n_333),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_405),
.B1(n_374),
.B2(n_385),
.Y(n_467)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_441),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_412),
.A2(n_349),
.B1(n_333),
.B2(n_331),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_427),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_405),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_352),
.C(n_339),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_409),
.A2(n_331),
.B1(n_347),
.B2(n_332),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_456),
.A2(n_395),
.B1(n_406),
.B2(n_414),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_427),
.A2(n_382),
.B1(n_388),
.B2(n_375),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_457),
.A2(n_458),
.B(n_459),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_449),
.A2(n_403),
.B(n_400),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_400),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_478),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_417),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_461),
.B(n_473),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_399),
.Y(n_462)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_462),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_469),
.B1(n_489),
.B2(n_450),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_449),
.A2(n_427),
.B(n_428),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_464),
.A2(n_477),
.B(n_485),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_440),
.Y(n_465)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_466),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_467),
.A2(n_456),
.B1(n_422),
.B2(n_423),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_430),
.A2(n_394),
.B1(n_371),
.B2(n_373),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_435),
.B(n_368),
.CI(n_434),
.CON(n_470),
.SN(n_470)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_474),
.Y(n_500)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_472),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_420),
.B(n_410),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_418),
.B(n_387),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_418),
.B(n_401),
.C(n_415),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_486),
.C(n_487),
.Y(n_501)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_416),
.Y(n_483)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_483),
.Y(n_513)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_428),
.A2(n_453),
.B(n_433),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_390),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_384),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_431),
.A2(n_407),
.B1(n_389),
.B2(n_376),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_426),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_426),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_444),
.B(n_436),
.C(n_439),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_433),
.C(n_442),
.Y(n_506)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_493),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_495),
.A2(n_518),
.B1(n_530),
.B2(n_516),
.Y(n_547)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_502),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_506),
.B(n_512),
.C(n_516),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_462),
.B(n_446),
.Y(n_508)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_446),
.Y(n_509)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_509),
.Y(n_535)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_445),
.C(n_434),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_487),
.B(n_437),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_514),
.B(n_527),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_443),
.C(n_432),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_336),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_517),
.B(n_500),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_454),
.Y(n_518)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_518),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_468),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_523),
.Y(n_537)
);

XOR2x2_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_405),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_SL g552 ( 
.A(n_520),
.B(n_377),
.C(n_369),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_530),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_419),
.C(n_421),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_485),
.C(n_457),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_477),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_438),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_470),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_467),
.A2(n_454),
.B1(n_451),
.B2(n_448),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_526),
.A2(n_458),
.B1(n_494),
.B2(n_463),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_492),
.B(n_421),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_475),
.Y(n_528)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_528),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_489),
.B(n_454),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_495),
.A2(n_459),
.B1(n_494),
.B2(n_488),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_534),
.A2(n_496),
.B1(n_497),
.B2(n_505),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_507),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_536),
.A2(n_539),
.B1(n_560),
.B2(n_505),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_538),
.B(n_546),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_521),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_540),
.B(n_514),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_542),
.A2(n_543),
.B1(n_547),
.B2(n_555),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_526),
.A2(n_491),
.B1(n_477),
.B2(n_464),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_470),
.C(n_482),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_544),
.B(n_549),
.C(n_553),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_509),
.B(n_465),
.Y(n_545)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_545),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_525),
.B(n_481),
.C(n_479),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_529),
.A2(n_438),
.B(n_452),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_550),
.A2(n_524),
.B(n_529),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_510),
.B(n_441),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_557),
.Y(n_571)
);

AO21x1_ASAP7_75t_L g570 ( 
.A1(n_552),
.A2(n_496),
.B(n_504),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_501),
.B(n_322),
.C(n_391),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_499),
.B(n_465),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_501),
.B(n_380),
.C(n_370),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_556),
.B(n_520),
.C(n_512),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_510),
.B(n_336),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_508),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_555),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_562),
.A2(n_566),
.B1(n_581),
.B2(n_583),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_563),
.A2(n_568),
.B(n_570),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_545),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_567),
.B(n_533),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_550),
.A2(n_524),
.B(n_504),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_537),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_549),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_572),
.B(n_575),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_559),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_573),
.B(n_582),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_556),
.C(n_533),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_541),
.Y(n_576)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_576),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_527),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_551),
.Y(n_594)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_541),
.Y(n_578)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_578),
.Y(n_600)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_559),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_579),
.A2(n_515),
.B1(n_574),
.B2(n_558),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_580),
.A2(n_542),
.B1(n_558),
.B2(n_531),
.Y(n_599)
);

BUFx24_ASAP7_75t_SL g582 ( 
.A(n_554),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_531),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_586),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_544),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_587),
.B(n_589),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_543),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_599),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_564),
.B(n_546),
.C(n_538),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_591),
.A2(n_596),
.B1(n_535),
.B2(n_579),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_572),
.B(n_506),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_601),
.Y(n_612)
);

MAJx2_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_598),
.C(n_561),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_583),
.A2(n_566),
.B1(n_565),
.B2(n_562),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_571),
.B(n_548),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_548),
.C(n_534),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_567),
.B(n_532),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_602),
.B(n_571),
.Y(n_615)
);

OAI321xp33_ASAP7_75t_L g603 ( 
.A1(n_588),
.A2(n_532),
.A3(n_565),
.B1(n_535),
.B2(n_576),
.C(n_578),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_603),
.B(n_607),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_590),
.B(n_498),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_605),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_595),
.B(n_580),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_561),
.C(n_577),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_SL g623 ( 
.A(n_606),
.B(n_611),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_592),
.A2(n_570),
.B(n_563),
.Y(n_607)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_609),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_613),
.B(n_598),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_596),
.A2(n_592),
.B1(n_600),
.B2(n_584),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_615),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_511),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_616),
.A2(n_528),
.B(n_503),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_513),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_617),
.B(n_618),
.C(n_552),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_599),
.B(n_601),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_607),
.A2(n_589),
.B(n_597),
.Y(n_619)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_619),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_343),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_623),
.B(n_613),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_624),
.A2(n_627),
.B(n_629),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_626),
.B(n_628),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_612),
.A2(n_594),
.B(n_515),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_610),
.B(n_503),
.C(n_344),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_608),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_630),
.B(n_332),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_629),
.B(n_606),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_632),
.B(n_634),
.Y(n_643)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_633),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_622),
.B(n_608),
.C(n_609),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_621),
.B(n_616),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_635),
.B(n_631),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_637),
.A2(n_638),
.B(n_622),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_639),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_641),
.B(n_642),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_643),
.A2(n_636),
.B(n_625),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_645),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_640),
.A2(n_637),
.B(n_639),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_646),
.A2(n_644),
.B1(n_647),
.B2(n_620),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_347),
.B1(n_324),
.B2(n_344),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_650),
.B(n_648),
.Y(n_651)
);

BUFx24_ASAP7_75t_SL g652 ( 
.A(n_651),
.Y(n_652)
);


endmodule