module fake_jpeg_909_n_136 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_56),
.Y(n_65)
);

BUFx12f_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_54),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_36),
.B1(n_43),
.B2(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_66),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_47),
.C(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_69),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_36),
.CI(n_37),
.CON(n_69),
.SN(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_0),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_52),
.B1(n_34),
.B2(n_33),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_38),
.B1(n_60),
.B2(n_37),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_79),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_86),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_86),
.B1(n_74),
.B2(n_68),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_60),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_0),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_13),
.B1(n_29),
.B2(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_1),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_7),
.B(n_8),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_103),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_3),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_107),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_11),
.C(n_25),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_108),
.C(n_9),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_88),
.B1(n_82),
.B2(n_92),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_7),
.B(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_3),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_4),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_21),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_116),
.C(n_101),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_118),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_99),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_113),
.B(n_96),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_119),
.C(n_114),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_121),
.B(n_115),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_110),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_123),
.B(n_117),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_111),
.Y(n_136)
);


endmodule