module fake_jpeg_24804_n_308 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_26),
.Y(n_66)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_27),
.B1(n_38),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_61),
.B1(n_28),
.B2(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_38),
.B1(n_27),
.B2(n_29),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_68),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_69),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_27),
.B1(n_38),
.B2(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_71),
.B1(n_76),
.B2(n_28),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_39),
.B1(n_49),
.B2(n_40),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_35),
.B1(n_31),
.B2(n_19),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_69),
.B1(n_73),
.B2(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_31),
.B1(n_19),
.B2(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_31),
.B1(n_36),
.B2(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_28),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_33),
.B1(n_24),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_32),
.B1(n_26),
.B2(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_79),
.B1(n_47),
.B2(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_10),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_36),
.B1(n_23),
.B2(n_18),
.Y(n_79)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_98),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_86),
.B(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_100),
.B1(n_58),
.B2(n_80),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_22),
.B1(n_23),
.B2(n_37),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_91),
.B1(n_95),
.B2(n_107),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_99),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_76),
.B1(n_65),
.B2(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_92),
.B(n_0),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_114),
.B(n_105),
.C(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_39),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_39),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_23),
.B1(n_37),
.B2(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_112),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_108),
.B1(n_70),
.B2(n_48),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_60),
.B1(n_62),
.B2(n_54),
.Y(n_107)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_49),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_39),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_39),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_117),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_49),
.B1(n_48),
.B2(n_40),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_1),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_125),
.B1(n_81),
.B2(n_83),
.Y(n_163)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_121),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_127),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_104),
.B1(n_103),
.B2(n_109),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_48),
.C(n_40),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_5),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_0),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_139),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_80),
.B(n_56),
.C(n_1),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_85),
.B(n_3),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_82),
.B(n_1),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_144),
.Y(n_181)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_82),
.B(n_2),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_92),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_151),
.A2(n_161),
.B(n_165),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_84),
.B1(n_95),
.B2(n_107),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_163),
.B1(n_174),
.B2(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_172),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_154),
.B(n_171),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_84),
.B(n_99),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_130),
.B(n_133),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_158),
.A2(n_160),
.B1(n_162),
.B2(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_115),
.B1(n_116),
.B2(n_112),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_86),
.C(n_106),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_86),
.B1(n_81),
.B2(n_90),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_85),
.B1(n_3),
.B2(n_5),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_179),
.B1(n_122),
.B2(n_134),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_137),
.C(n_124),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_6),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_119),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_150),
.Y(n_183)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_182),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_195),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_123),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_199),
.C(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_154),
.B(n_166),
.C(n_142),
.D(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_160),
.B1(n_158),
.B2(n_179),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_143),
.Y(n_195)
);

NAND2x1_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_131),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_203),
.B(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_152),
.B(n_151),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_134),
.B(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_210),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_208),
.B1(n_174),
.B2(n_166),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_142),
.B1(n_146),
.B2(n_138),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_127),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_189),
.A3(n_192),
.B1(n_194),
.B2(n_188),
.C1(n_200),
.C2(n_198),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_184),
.B1(n_206),
.B2(n_208),
.Y(n_236)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_219),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_197),
.B1(n_172),
.B2(n_155),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_169),
.C(n_149),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_231),
.C(n_128),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_201),
.Y(n_238)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_164),
.B1(n_168),
.B2(n_167),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_168),
.B1(n_193),
.B2(n_186),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_155),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_233),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_149),
.C(n_121),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_196),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_201),
.B(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_247),
.B1(n_248),
.B2(n_220),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_221),
.C(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_239),
.C(n_243),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_244),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_199),
.C(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_205),
.C(n_185),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_205),
.C(n_195),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_252),
.C(n_222),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_246),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_186),
.B1(n_203),
.B2(n_202),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_190),
.B1(n_209),
.B2(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_228),
.B1(n_227),
.B2(n_222),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_183),
.Y(n_251)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

AO21x2_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_223),
.B(n_220),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_268),
.B1(n_223),
.B2(n_218),
.Y(n_272)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_259),
.B(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_237),
.C(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_265),
.B(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_224),
.B1(n_219),
.B2(n_232),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_239),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_261),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_271),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_279),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_253),
.C(n_261),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_243),
.C(n_245),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_277),
.C(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_252),
.C(n_255),
.Y(n_277)
);

AOI31xp67_ASAP7_75t_SL g279 ( 
.A1(n_255),
.A2(n_238),
.A3(n_214),
.B(n_187),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_256),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_269),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_257),
.B1(n_178),
.B2(n_153),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_293),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_278),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_295),
.B1(n_270),
.B2(n_280),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_299),
.B1(n_300),
.B2(n_147),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_283),
.B1(n_276),
.B2(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_276),
.B1(n_277),
.B2(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_281),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_302),
.A3(n_303),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_264),
.A3(n_275),
.B1(n_274),
.B2(n_272),
.C1(n_147),
.C2(n_141),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_300),
.C(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.C(n_12),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_12),
.B(n_14),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_14),
.Y(n_308)
);


endmodule