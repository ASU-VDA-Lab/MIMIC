module fake_aes_1002_n_678 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_678);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_678;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_195;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_41), .Y(n_77) );
OR2x2_ASAP7_75t_L g78 ( .A(n_45), .B(n_50), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_48), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_26), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_1), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_73), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_44), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_49), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_6), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_10), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_15), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_54), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_14), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_75), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_11), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_37), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_31), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_66), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_57), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_19), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_23), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_70), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_69), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_52), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_59), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_65), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_34), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_20), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_27), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_56), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_61), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_68), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_64), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_39), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_8), .Y(n_123) );
CKINVDCx6p67_ASAP7_75t_R g124 ( .A(n_97), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_79), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_97), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_86), .B(n_0), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_121), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_120), .B(n_2), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_112), .B(n_2), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_92), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_77), .B(n_3), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_96), .B(n_3), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_98), .B(n_4), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_110), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_99), .B(n_4), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_87), .B(n_5), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_87), .B(n_5), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_114), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_131), .B(n_116), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_159), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_159), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_160), .B(n_101), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_125), .B(n_118), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_126), .B(n_119), .Y(n_175) );
BUFx10_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_160), .Y(n_178) );
INVx5_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_129), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_124), .B(n_102), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_124), .B(n_85), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_127), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_127), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_129), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
INVxp33_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
OR2x6_ASAP7_75t_L g189 ( .A(n_130), .B(n_95), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_126), .B(n_85), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_128), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_130), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
OR2x6_ASAP7_75t_L g196 ( .A(n_134), .B(n_95), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_128), .Y(n_197) );
AO22x2_ASAP7_75t_L g198 ( .A1(n_135), .A2(n_93), .B1(n_116), .B2(n_109), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_140), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
CKINVDCx14_ASAP7_75t_R g201 ( .A(n_162), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
BUFx4_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
AND2x6_ASAP7_75t_L g206 ( .A(n_135), .B(n_105), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_138), .B(n_109), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_138), .B(n_117), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_139), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_139), .A2(n_123), .B1(n_94), .B2(n_107), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_141), .B(n_89), .Y(n_215) );
INVx4_ASAP7_75t_SL g216 ( .A(n_141), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_144), .Y(n_218) );
AND2x6_ASAP7_75t_L g219 ( .A(n_142), .B(n_106), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_151), .B(n_78), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_142), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_145), .A2(n_123), .B1(n_94), .B2(n_88), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_145), .B(n_113), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_147), .B(n_78), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_157), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_201), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_193), .B(n_192), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_177), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_211), .B(n_165), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_193), .A2(n_165), .B1(n_164), .B2(n_163), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_173), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_177), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_193), .B(n_164), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_190), .B(n_163), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_201), .Y(n_238) );
NAND3xp33_ASAP7_75t_SL g239 ( .A(n_214), .B(n_158), .C(n_152), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_192), .B(n_161), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_200), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_198), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_198), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_188), .B(n_161), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_176), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_173), .A2(n_156), .B1(n_155), .B2(n_147), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_173), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_174), .B(n_156), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_189), .A2(n_155), .B1(n_153), .B2(n_150), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_176), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_168), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_192), .B(n_153), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_167), .Y(n_258) );
OR2x6_ASAP7_75t_L g259 ( .A(n_189), .B(n_150), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_167), .Y(n_260) );
BUFx12f_ASAP7_75t_L g261 ( .A(n_189), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_196), .B(n_157), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_181), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_224), .B(n_111), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_196), .B(n_133), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_196), .B(n_133), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_172), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_188), .B(n_88), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_171), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_176), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_171), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_221), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_221), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_196), .B(n_82), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_172), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_173), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_173), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_180), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_203), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_224), .B(n_103), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_186), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_222), .B(n_115), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_166), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_173), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_221), .B(n_82), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_222), .B(n_88), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_221), .B(n_88), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_259), .B(n_208), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_228), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_259), .A2(n_178), .B1(n_170), .B2(n_169), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_230), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_228), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_241), .B(n_166), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_230), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_259), .B(n_166), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_244), .A2(n_206), .B1(n_219), .B2(n_225), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_254), .B(n_216), .Y(n_301) );
INVx3_ASAP7_75t_SL g302 ( .A(n_274), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_244), .A2(n_206), .B1(n_219), .B2(n_225), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_237), .A2(n_210), .B(n_175), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_238), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_231), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_245), .A2(n_219), .B1(n_206), .B2(n_208), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_245), .A2(n_219), .B1(n_206), .B2(n_208), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_251), .A2(n_206), .B1(n_219), .B2(n_215), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_238), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_235), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_241), .B(n_223), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_SL g315 ( .A1(n_289), .A2(n_175), .B(n_210), .C(n_217), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_229), .B(n_205), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_235), .Y(n_317) );
BUFx12f_ASAP7_75t_L g318 ( .A(n_261), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_261), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_229), .B(n_216), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_251), .A2(n_219), .B1(n_206), .B2(n_205), .Y(n_323) );
OAI22x1_ASAP7_75t_L g324 ( .A1(n_254), .A2(n_204), .B1(n_184), .B2(n_191), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_277), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_281), .Y(n_328) );
AOI33xp33_ASAP7_75t_L g329 ( .A1(n_268), .A2(n_226), .A3(n_213), .B1(n_209), .B2(n_186), .B3(n_212), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_229), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_236), .A2(n_183), .B(n_182), .Y(n_331) );
CKINVDCx8_ASAP7_75t_R g332 ( .A(n_274), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_241), .B(n_207), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_229), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_262), .B(n_207), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_282), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_240), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_282), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_227), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_234), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_321), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_326), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_314), .A2(n_239), .B(n_283), .C(n_264), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_291), .B(n_243), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_306), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_321), .A2(n_253), .B1(n_290), .B2(n_288), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_291), .A2(n_232), .B1(n_262), .B2(n_233), .Y(n_348) );
AO221x2_ASAP7_75t_L g349 ( .A1(n_324), .A2(n_253), .B1(n_252), .B2(n_257), .C(n_273), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_295), .Y(n_350) );
INVx8_ASAP7_75t_L g351 ( .A(n_291), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_327), .A2(n_290), .B1(n_288), .B2(n_262), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_305), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_291), .A2(n_273), .B1(n_266), .B2(n_265), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_327), .A2(n_290), .B1(n_288), .B2(n_265), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_298), .A2(n_286), .B1(n_275), .B2(n_265), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_298), .B(n_247), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_299), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_302), .B(n_266), .Y(n_363) );
INVx6_ASAP7_75t_L g364 ( .A(n_299), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_299), .B(n_250), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_299), .A2(n_275), .B1(n_266), .B2(n_279), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_318), .Y(n_369) );
INVx6_ASAP7_75t_L g370 ( .A(n_299), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_296), .B(n_258), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_332), .A2(n_249), .B1(n_285), .B2(n_276), .C(n_260), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
INVx4_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_342), .A2(n_332), .B(n_331), .C(n_338), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_361), .A2(n_302), .B1(n_334), .B2(n_330), .C(n_328), .Y(n_376) );
AO21x1_ASAP7_75t_SL g377 ( .A1(n_354), .A2(n_338), .B(n_336), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_350), .B(n_324), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_355), .B(n_302), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_275), .B1(n_334), .B2(n_336), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_346), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_360), .B(n_316), .Y(n_382) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_351), .A2(n_369), .B(n_363), .Y(n_383) );
AO21x1_ASAP7_75t_L g384 ( .A1(n_341), .A2(n_293), .B(n_301), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_349), .A2(n_310), .B1(n_268), .B2(n_316), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_354), .A2(n_308), .B1(n_307), .B2(n_309), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_366), .B(n_311), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_352), .B(n_311), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_343), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_344), .A2(n_303), .B(n_300), .C(n_304), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_349), .A2(n_318), .B1(n_292), .B2(n_337), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_353), .B(n_294), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_345), .A2(n_319), .B1(n_333), .B2(n_335), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_348), .A2(n_339), .B(n_294), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_365), .A2(n_297), .B(n_317), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_345), .A2(n_317), .B1(n_312), .B2(n_311), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_359), .A2(n_329), .B(n_184), .C(n_197), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_397), .A2(n_297), .B(n_317), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_396), .A2(n_361), .B1(n_371), .B2(n_372), .C(n_356), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_376), .A2(n_358), .B(n_371), .C(n_347), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_382), .B(n_351), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_358), .B(n_347), .C(n_368), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_373), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_382), .B(n_351), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_392), .B(n_357), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_375), .A2(n_276), .A3(n_258), .B(n_260), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_394), .A2(n_88), .B1(n_100), .B2(n_104), .C1(n_185), .C2(n_197), .Y(n_413) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_375), .A2(n_154), .B(n_185), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_389), .A2(n_357), .B1(n_364), .B2(n_370), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_386), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_357), .B1(n_364), .B2(n_370), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_390), .B(n_362), .Y(n_420) );
BUFx12f_ASAP7_75t_L g421 ( .A(n_374), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_400), .A2(n_364), .B1(n_370), .B2(n_362), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_399), .A2(n_323), .B1(n_362), .B2(n_312), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_399), .A2(n_312), .B1(n_278), .B2(n_279), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_391), .B(n_386), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_378), .B(n_146), .C(n_154), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_385), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_388), .A2(n_287), .B1(n_278), .B2(n_340), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_380), .A2(n_287), .B1(n_340), .B2(n_367), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_374), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_400), .A2(n_313), .B1(n_337), .B2(n_185), .C(n_184), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_385), .B(n_339), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_387), .A3(n_393), .B(n_379), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_416), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_425), .B(n_385), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_421), .A2(n_387), .B1(n_374), .B2(n_395), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_425), .B(n_395), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_403), .B(n_398), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_426), .B(n_395), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_430), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_402), .A2(n_383), .B1(n_393), .B2(n_374), .C(n_397), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_428), .B(n_398), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g448 ( .A(n_433), .B(n_383), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_412), .B(n_398), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_417), .B(n_384), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_407), .A2(n_367), .B(n_322), .C(n_197), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_428), .B(n_384), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_413), .A2(n_377), .B1(n_367), .B2(n_191), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_429), .B(n_377), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_404), .A2(n_191), .B1(n_337), .B2(n_313), .C(n_154), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_420), .B(n_7), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_420), .B(n_7), .Y(n_458) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_401), .B(n_339), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_404), .A2(n_337), .B1(n_313), .B2(n_322), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_435), .B(n_8), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_435), .B(n_9), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_408), .B(n_46), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_427), .B(n_146), .C(n_154), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_408), .B(n_9), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_408), .B(n_10), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
OAI31xp33_ASAP7_75t_SL g468 ( .A1(n_410), .A2(n_322), .A3(n_12), .B(n_13), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_421), .A2(n_313), .B1(n_320), .B2(n_322), .Y(n_469) );
INVx4_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_406), .B(n_11), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_408), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_401), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_401), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_418), .B(n_53), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_418), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_418), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
OAI211xp5_ASAP7_75t_SL g479 ( .A1(n_415), .A2(n_315), .B(n_212), .C(n_195), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_418), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_419), .Y(n_481) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_414), .A2(n_220), .B(n_195), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_434), .A2(n_146), .B1(n_240), .B2(n_267), .C(n_272), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_433), .B(n_13), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_411), .B(n_146), .C(n_179), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_439), .B(n_442), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_455), .B(n_470), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_465), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
OAI21x1_ASAP7_75t_L g490 ( .A1(n_459), .A2(n_423), .B(n_422), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_437), .B(n_433), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_440), .B(n_409), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_455), .B(n_433), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_465), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_449), .B(n_14), .Y(n_495) );
AOI22x1_ASAP7_75t_L g496 ( .A1(n_470), .A2(n_146), .B1(n_16), .B2(n_17), .Y(n_496) );
AOI33xp33_ASAP7_75t_L g497 ( .A1(n_457), .A2(n_15), .A3(n_16), .B1(n_17), .B2(n_18), .B3(n_220), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_461), .B(n_18), .Y(n_498) );
AND4x1_ASAP7_75t_L g499 ( .A(n_468), .B(n_24), .C(n_28), .D(n_29), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_437), .B(n_432), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_445), .Y(n_501) );
AND3x2_ASAP7_75t_L g502 ( .A(n_484), .B(n_438), .C(n_462), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_459), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_461), .B(n_146), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
NAND2x1_ASAP7_75t_L g506 ( .A(n_470), .B(n_424), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_450), .B(n_431), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_484), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
AND4x1_ASAP7_75t_L g510 ( .A(n_485), .B(n_30), .C(n_32), .D(n_35), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_462), .B(n_179), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_444), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_446), .B(n_179), .C(n_187), .Y(n_513) );
NOR2x1p5_ASAP7_75t_L g514 ( .A(n_485), .B(n_340), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_457), .B(n_38), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_458), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_458), .B(n_40), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_436), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_436), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_456), .A2(n_270), .A3(n_248), .B(n_255), .Y(n_521) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_448), .B(n_320), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_443), .B(n_179), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_443), .B(n_179), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_447), .B(n_42), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_447), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_466), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_481), .B(n_43), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_455), .B(n_47), .Y(n_529) );
OAI33xp33_ASAP7_75t_L g530 ( .A1(n_471), .A2(n_194), .A3(n_269), .B1(n_256), .B2(n_271), .B3(n_284), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_481), .B(n_51), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_455), .B(n_55), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_451), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_473), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_473), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_474), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_441), .B(n_58), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_448), .B(n_60), .Y(n_538) );
NAND4xp25_ASAP7_75t_L g539 ( .A(n_454), .B(n_194), .C(n_267), .D(n_272), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_453), .B(n_62), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_453), .B(n_63), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_452), .B(n_272), .C(n_267), .D(n_280), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_512), .B(n_474), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_489), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_517), .B(n_460), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_534), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_497), .B(n_479), .C(n_483), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_526), .B(n_486), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_529), .B(n_475), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_487), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_499), .B(n_469), .C(n_476), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_498), .B(n_480), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_513), .B(n_464), .C(n_475), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_509), .B(n_480), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_526), .B(n_472), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_495), .B(n_463), .C(n_475), .D(n_477), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_491), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_491), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_493), .B(n_463), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_535), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_519), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_478), .Y(n_564) );
AND3x2_ASAP7_75t_L g565 ( .A(n_493), .B(n_475), .C(n_463), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_536), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_533), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_488), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_494), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_527), .B(n_478), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_529), .B(n_477), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_531), .B(n_467), .C(n_256), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_514), .B(n_467), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_520), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_508), .B(n_482), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_504), .B(n_482), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_487), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_523), .B(n_67), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_500), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_496), .B(n_187), .C(n_218), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_507), .B(n_76), .Y(n_582) );
AOI211xp5_ASAP7_75t_SL g583 ( .A1(n_532), .A2(n_271), .B(n_269), .C(n_284), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_522), .B(n_320), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_507), .B(n_187), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_525), .B(n_187), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_540), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_541), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_578), .B(n_502), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_573), .A2(n_516), .B1(n_518), .B2(n_506), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_551), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_577), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_580), .B(n_502), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_567), .B(n_568), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_558), .A2(n_542), .B(n_537), .C(n_521), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_581), .A2(n_530), .B(n_503), .Y(n_598) );
OAI211xp5_ASAP7_75t_L g599 ( .A1(n_558), .A2(n_539), .B(n_515), .C(n_503), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_549), .B(n_515), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_559), .Y(n_601) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_584), .A2(n_511), .B1(n_525), .B2(n_530), .C1(n_538), .C2(n_490), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_553), .A2(n_528), .B(n_510), .C(n_218), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_547), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_583), .A2(n_320), .B1(n_250), .B2(n_255), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_564), .Y(n_606) );
XNOR2x2_ASAP7_75t_L g607 ( .A(n_552), .B(n_320), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_560), .B(n_218), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_544), .Y(n_609) );
XOR2x2_ASAP7_75t_L g610 ( .A(n_550), .B(n_270), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_563), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_590), .B(n_218), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_562), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_581), .A2(n_250), .B(n_320), .C(n_248), .Y(n_614) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_573), .A2(n_571), .B(n_550), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_545), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_588), .B(n_227), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_556), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_554), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_543), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_589), .B(n_246), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
OAI31xp33_ASAP7_75t_L g625 ( .A1(n_552), .A2(n_280), .A3(n_250), .B(n_216), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_570), .Y(n_626) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_571), .B(n_250), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_546), .B(n_586), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_572), .A2(n_250), .B(n_216), .Y(n_629) );
AO21x1_ASAP7_75t_L g630 ( .A1(n_561), .A2(n_555), .B(n_585), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_585), .B(n_246), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_575), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_548), .A2(n_246), .B(n_263), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_565), .B(n_246), .Y(n_635) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_579), .B(n_263), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_582), .B(n_263), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_551), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_547), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_568), .B(n_263), .C(n_569), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_578), .B(n_263), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_558), .A2(n_468), .B(n_441), .C(n_583), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_639), .Y(n_644) );
NAND2xp33_ASAP7_75t_SL g645 ( .A(n_639), .B(n_592), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_596), .A2(n_624), .B1(n_621), .B2(n_633), .C(n_626), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_591), .A2(n_595), .B1(n_630), .B2(n_597), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g648 ( .A1(n_593), .A2(n_594), .A3(n_603), .B1(n_619), .B2(n_600), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_632), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_615), .A2(n_641), .B1(n_598), .B2(n_628), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_606), .B(n_611), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_599), .A2(n_643), .B1(n_614), .B2(n_601), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_625), .B(n_602), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_610), .A2(n_614), .B(n_605), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_634), .B(n_623), .C(n_637), .Y(n_655) );
OAI32xp33_ASAP7_75t_L g656 ( .A1(n_607), .A2(n_596), .A3(n_620), .B1(n_613), .B2(n_617), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_645), .A2(n_616), .B1(n_609), .B2(n_622), .C(n_638), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_649), .Y(n_658) );
AO22x2_ASAP7_75t_L g659 ( .A1(n_652), .A2(n_607), .B1(n_611), .B2(n_604), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_646), .B(n_604), .Y(n_660) );
OAI321xp33_ASAP7_75t_L g661 ( .A1(n_648), .A2(n_635), .A3(n_623), .B1(n_605), .B2(n_637), .C(n_642), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_651), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_647), .A2(n_610), .B1(n_636), .B2(n_627), .C(n_640), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_644), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_659), .A2(n_656), .B1(n_650), .B2(n_653), .C(n_654), .Y(n_665) );
AO22x1_ASAP7_75t_L g666 ( .A1(n_664), .A2(n_655), .B1(n_635), .B2(n_629), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_657), .A2(n_627), .B(n_631), .Y(n_667) );
INVx2_ASAP7_75t_SL g668 ( .A(n_658), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_668), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_665), .Y(n_670) );
OR4x2_ASAP7_75t_L g671 ( .A(n_666), .B(n_659), .C(n_661), .D(n_663), .Y(n_671) );
XNOR2xp5_ASAP7_75t_L g672 ( .A(n_670), .B(n_669), .Y(n_672) );
XOR2x2_ASAP7_75t_L g673 ( .A(n_671), .B(n_667), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_672), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_673), .B(n_660), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_675), .B1(n_671), .B2(n_662), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_642), .B1(n_608), .B2(n_618), .C(n_612), .Y(n_678) );
endmodule