module real_jpeg_11634_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_82),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_82),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_7),
.B(n_138),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_102),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_7),
.B(n_66),
.C(n_85),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_36),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_7),
.A2(n_69),
.B(n_166),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_27),
.B(n_35),
.C(n_193),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_102),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_8),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_30),
.B1(n_65),
.B2(n_66),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_42),
.B1(n_65),
.B2(n_66),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_48),
.B1(n_65),
.B2(n_66),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_15),
.B(n_28),
.Y(n_62)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_104),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_90),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_21),
.A2(n_22),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_57),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_57),
.C(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_26),
.A2(n_31),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g60 ( 
.A1(n_27),
.A2(n_46),
.A3(n_50),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_31),
.A2(n_40),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_32),
.B(n_41),
.Y(n_121)
);

NOR2x1_ASAP7_75t_R g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_34),
.A2(n_37),
.B(n_102),
.Y(n_193)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_38),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_38),
.B(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B(n_51),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_44),
.A2(n_49),
.B1(n_53),
.B2(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_53),
.B(n_102),
.C(n_103),
.Y(n_101)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_75),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_64),
.A2(n_69),
.B1(n_75),
.B2(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_71),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_66),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_65),
.B(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_75),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_69),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_70),
.A2(n_71),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_70),
.B(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_71),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_75),
.A2(n_172),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_75),
.B(n_102),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_75),
.A2(n_140),
.B(n_180),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_76),
.B(n_90),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_80),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_83),
.A2(n_89),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_87),
.A2(n_93),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_87),
.B(n_102),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_94),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_98),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_91),
.B(n_95),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_96),
.A2(n_97),
.B(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_99),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_123),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_115),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_144),
.B(n_224),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_141),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_128),
.B(n_141),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_134),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_132),
.B(n_134),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.C(n_139),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_219),
.B(n_223),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_204),
.B(n_218),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_188),
.B(n_203),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_168),
.B(n_187),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_151),
.B1(n_155),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_152),
.A2(n_154),
.B(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_176),
.B(n_186),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_174),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_181),
.B(n_185),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_190),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_198),
.C(n_202),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_194),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_206),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_214),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);


endmodule