module real_aes_7975_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g455 ( .A1(n_0), .A2(n_156), .B(n_456), .C(n_459), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_1), .B(n_450), .Y(n_460) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
INVx1_ASAP7_75t_L g154 ( .A(n_3), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_4), .B(n_157), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_5), .A2(n_445), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_6), .A2(n_179), .B(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_7), .A2(n_38), .B1(n_144), .B2(n_202), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_8), .A2(n_9), .B1(n_707), .B2(n_708), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_8), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_9), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_10), .B(n_179), .Y(n_187) );
AND2x6_ASAP7_75t_L g159 ( .A(n_11), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_12), .A2(n_159), .B(n_436), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_13), .B(n_39), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_13), .B(n_39), .Y(n_119) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
INVx1_ASAP7_75t_L g135 ( .A(n_15), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_16), .B(n_140), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_17), .B(n_157), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_18), .B(n_131), .Y(n_189) );
AO32x2_ASAP7_75t_L g240 ( .A1(n_19), .A2(n_130), .A3(n_173), .B1(n_179), .B2(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_20), .A2(n_30), .B1(n_121), .B2(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_20), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_21), .B(n_144), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_22), .B(n_131), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_23), .A2(n_55), .B1(n_144), .B2(n_202), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_24), .A2(n_81), .B1(n_140), .B2(n_144), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_25), .B(n_144), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_26), .A2(n_173), .B(n_436), .C(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_27), .A2(n_173), .B(n_436), .C(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_29), .B(n_175), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_30), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_30), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_31), .A2(n_445), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_32), .B(n_175), .Y(n_217) );
INVx2_ASAP7_75t_L g142 ( .A(n_33), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_34), .A2(n_442), .B(n_485), .C(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_35), .B(n_144), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_36), .B(n_175), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_37), .B(n_224), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_40), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_41), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_42), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_43), .B(n_157), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_44), .B(n_445), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_45), .A2(n_442), .B(n_485), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_46), .B(n_144), .Y(n_182) );
INVx1_ASAP7_75t_L g457 ( .A(n_47), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_48), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_49), .A2(n_90), .B1(n_202), .B2(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g510 ( .A(n_50), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_51), .B(n_144), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_52), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_53), .B(n_445), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_54), .B(n_152), .Y(n_186) );
AOI22xp33_ASAP7_75t_SL g193 ( .A1(n_56), .A2(n_60), .B1(n_140), .B2(n_144), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_57), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_58), .B(n_144), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_59), .B(n_144), .Y(n_221) );
INVx1_ASAP7_75t_L g160 ( .A(n_61), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_62), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_63), .B(n_450), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_64), .A2(n_146), .B(n_152), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_65), .B(n_144), .Y(n_155) );
INVx1_ASAP7_75t_L g134 ( .A(n_66), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_67), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_68), .B(n_157), .Y(n_488) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_69), .A2(n_173), .A3(n_179), .B1(n_200), .B2(n_205), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_70), .B(n_158), .Y(n_501) );
INVx1_ASAP7_75t_L g169 ( .A(n_71), .Y(n_169) );
INVx1_ASAP7_75t_L g212 ( .A(n_72), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_73), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_74), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_75), .A2(n_436), .B(n_438), .C(n_442), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_76), .B(n_140), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_77), .Y(n_519) );
INVx1_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_79), .A2(n_103), .B1(n_112), .B2(n_736), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_80), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_82), .B(n_202), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_83), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_84), .B(n_140), .Y(n_216) );
INVx2_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_86), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_87), .B(n_172), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_88), .B(n_140), .Y(n_183) );
INVx2_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
OR2x2_ASAP7_75t_L g116 ( .A(n_89), .B(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g724 ( .A(n_89), .B(n_716), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_91), .A2(n_101), .B1(n_140), .B2(n_141), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_92), .B(n_445), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_93), .Y(n_487) );
INVxp67_ASAP7_75t_L g522 ( .A(n_94), .Y(n_522) );
XNOR2xp5_ASAP7_75t_L g725 ( .A(n_95), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_96), .B(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_97), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g439 ( .A(n_98), .Y(n_439) );
INVx1_ASAP7_75t_L g497 ( .A(n_99), .Y(n_497) );
AND2x2_ASAP7_75t_L g512 ( .A(n_100), .B(n_175), .Y(n_512) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g736 ( .A(n_105), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g427 ( .A(n_108), .B(n_117), .Y(n_427) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_108), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO221x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_718), .B1(n_721), .B2(n_730), .C(n_732), .Y(n_112) );
OAI222xp33_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_706), .B1(n_709), .B2(n_713), .C1(n_714), .C2(n_717), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B1(n_426), .B2(n_428), .Y(n_114) );
INVx2_ASAP7_75t_L g711 ( .A(n_115), .Y(n_711) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g716 ( .A(n_117), .Y(n_716) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_120), .A2(n_428), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_122), .A2(n_123), .B1(n_727), .B2(n_729), .Y(n_726) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR5x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_317), .C(n_375), .D(n_411), .E(n_418), .Y(n_123) );
NAND3xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_263), .C(n_287), .Y(n_124) );
AOI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_195), .B1(n_229), .B2(n_234), .C(n_244), .Y(n_125) );
OAI21xp5_ASAP7_75t_SL g397 ( .A1(n_126), .A2(n_398), .B(n_400), .Y(n_397) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_176), .Y(n_126) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_127), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
INVx2_ASAP7_75t_L g233 ( .A(n_128), .Y(n_233) );
AND2x2_ASAP7_75t_L g246 ( .A(n_128), .B(n_178), .Y(n_246) );
AND2x2_ASAP7_75t_L g300 ( .A(n_128), .B(n_177), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_128), .B(n_163), .Y(n_315) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_161), .Y(n_128) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_129), .A2(n_164), .B(n_174), .Y(n_163) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_130), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_132), .B(n_133), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_150), .B(n_159), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_143), .C(n_146), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_139), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_139), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
INVx1_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx3_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_144), .Y(n_441) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
AND2x6_ASAP7_75t_L g436 ( .A(n_145), .B(n_437), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g438 ( .A1(n_146), .A2(n_439), .B(n_440), .C(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_147), .A2(n_215), .B(n_216), .Y(n_214) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g469 ( .A(n_148), .Y(n_469) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx1_ASAP7_75t_L g224 ( .A(n_149), .Y(n_224) );
INVx1_ASAP7_75t_L g437 ( .A(n_149), .Y(n_437) );
AND2x2_ASAP7_75t_L g446 ( .A(n_149), .B(n_153), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_155), .C(n_156), .Y(n_150) );
O2A1O1Ixp5_ASAP7_75t_L g168 ( .A1(n_151), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_151), .A2(n_468), .B(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_156), .A2(n_185), .B(n_186), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_156), .A2(n_172), .B1(n_192), .B2(n_193), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_156), .A2(n_172), .B1(n_242), .B2(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_157), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_157), .A2(n_182), .B(n_183), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_SL g210 ( .A1(n_157), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_157), .B(n_522), .Y(n_521) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_158), .A2(n_172), .B1(n_201), .B2(n_204), .Y(n_200) );
BUFx3_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_159), .A2(n_181), .B(n_184), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .B(n_214), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_159), .A2(n_220), .B(n_225), .Y(n_219) );
INVx4_ASAP7_75t_SL g443 ( .A(n_159), .Y(n_443) );
AND2x4_ASAP7_75t_L g445 ( .A(n_159), .B(n_446), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_159), .B(n_446), .Y(n_498) );
AND2x2_ASAP7_75t_L g333 ( .A(n_162), .B(n_274), .Y(n_333) );
AND2x2_ASAP7_75t_L g366 ( .A(n_162), .B(n_178), .Y(n_366) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g273 ( .A(n_163), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g286 ( .A(n_163), .B(n_178), .Y(n_286) );
AND2x2_ASAP7_75t_L g293 ( .A(n_163), .B(n_274), .Y(n_293) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_163), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_163), .B(n_177), .Y(n_309) );
INVx1_ASAP7_75t_L g340 ( .A(n_163), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_173), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_171), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g458 ( .A(n_172), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g190 ( .A(n_173), .B(n_191), .C(n_194), .Y(n_190) );
INVx2_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_175), .A2(n_209), .B(n_217), .Y(n_208) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_175), .A2(n_219), .B(n_228), .Y(n_218) );
INVx1_ASAP7_75t_L g475 ( .A(n_175), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_175), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_175), .A2(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g316 ( .A(n_176), .Y(n_316) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_188), .Y(n_176) );
INVx2_ASAP7_75t_L g272 ( .A(n_177), .Y(n_272) );
AND2x2_ASAP7_75t_L g294 ( .A(n_177), .B(n_233), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_177), .B(n_340), .Y(n_345) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_178), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g417 ( .A(n_178), .B(n_381), .Y(n_417) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_187), .Y(n_178) );
INVx4_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_179), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_179), .A2(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g231 ( .A(n_188), .Y(n_231) );
INVx3_ASAP7_75t_L g332 ( .A(n_188), .Y(n_332) );
OR2x2_ASAP7_75t_L g362 ( .A(n_188), .B(n_363), .Y(n_362) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_188), .B(n_272), .Y(n_388) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g275 ( .A(n_189), .Y(n_275) );
AO21x1_ASAP7_75t_L g274 ( .A1(n_191), .A2(n_194), .B(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_194), .A2(n_434), .B(n_447), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_194), .B(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g450 ( .A(n_194), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_194), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_194), .A2(n_496), .B(n_503), .Y(n_495) );
AOI33xp33_ASAP7_75t_L g408 ( .A1(n_195), .A2(n_246), .A3(n_260), .B1(n_332), .B2(n_409), .B3(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
OR2x2_ASAP7_75t_L g261 ( .A(n_197), .B(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_197), .B(n_258), .Y(n_320) );
OR2x2_ASAP7_75t_L g373 ( .A(n_197), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g299 ( .A(n_198), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g324 ( .A(n_198), .B(n_206), .Y(n_324) );
AND2x2_ASAP7_75t_L g391 ( .A(n_198), .B(n_236), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_198), .A2(n_291), .B(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
INVx1_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
AND2x2_ASAP7_75t_L g270 ( .A(n_199), .B(n_240), .Y(n_270) );
AND2x2_ASAP7_75t_L g319 ( .A(n_199), .B(n_239), .Y(n_319) );
INVx2_ASAP7_75t_L g459 ( .A(n_203), .Y(n_459) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_203), .Y(n_489) );
INVx1_ASAP7_75t_L g472 ( .A(n_205), .Y(n_472) );
INVx2_ASAP7_75t_SL g361 ( .A(n_206), .Y(n_361) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
INVx2_ASAP7_75t_L g281 ( .A(n_207), .Y(n_281) );
INVx1_ASAP7_75t_L g412 ( .A(n_207), .Y(n_412) );
AND2x2_ASAP7_75t_L g425 ( .A(n_207), .B(n_306), .Y(n_425) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
OR2x2_ASAP7_75t_L g258 ( .A(n_208), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_218), .Y(n_236) );
AND2x2_ASAP7_75t_L g253 ( .A(n_218), .B(n_239), .Y(n_253) );
INVx1_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
INVx1_ASAP7_75t_L g266 ( .A(n_218), .Y(n_266) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_240), .Y(n_291) );
INVx2_ASAP7_75t_L g307 ( .A(n_218), .Y(n_307) );
AND2x2_ASAP7_75t_L g400 ( .A(n_218), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_218), .B(n_281), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
INVx1_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_231), .B(n_315), .Y(n_381) );
INVx1_ASAP7_75t_SL g341 ( .A(n_232), .Y(n_341) );
INVx2_ASAP7_75t_L g262 ( .A(n_233), .Y(n_262) );
AND2x2_ASAP7_75t_L g331 ( .A(n_233), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g347 ( .A(n_233), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
INVx1_ASAP7_75t_L g409 ( .A(n_235), .Y(n_409) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g367 ( .A(n_237), .B(n_357), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_237), .A2(n_378), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g280 ( .A(n_238), .B(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
INVx1_ASAP7_75t_L g329 ( .A(n_238), .Y(n_329) );
OR2x2_ASAP7_75t_L g393 ( .A(n_239), .B(n_252), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_239), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g306 ( .A(n_240), .B(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B1(n_254), .B2(n_256), .Y(n_244) );
OR2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_273), .Y(n_323) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_246), .A2(n_365), .B1(n_367), .B2(n_368), .C1(n_369), .C2(n_372), .Y(n_364) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g311 ( .A(n_250), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_252), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_252), .Y(n_336) );
AND2x2_ASAP7_75t_L g384 ( .A(n_252), .B(n_253), .Y(n_384) );
INVx1_ASAP7_75t_L g402 ( .A(n_252), .Y(n_402) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g368 ( .A(n_255), .B(n_294), .Y(n_368) );
AND2x2_ASAP7_75t_L g410 ( .A(n_255), .B(n_286), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_257), .B(n_305), .Y(n_392) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_258), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g285 ( .A(n_262), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g353 ( .A(n_262), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B(n_271), .C(n_276), .Y(n_263) );
INVxp67_ASAP7_75t_L g277 ( .A(n_264), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_265), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_265), .B(n_312), .Y(n_407) );
BUFx3_ASAP7_75t_L g371 ( .A(n_266), .Y(n_371) );
INVx1_ASAP7_75t_L g278 ( .A(n_267), .Y(n_278) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g297 ( .A(n_269), .B(n_291), .Y(n_297) );
INVx1_ASAP7_75t_SL g337 ( .A(n_270), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g327 ( .A(n_272), .Y(n_327) );
AND2x2_ASAP7_75t_L g350 ( .A(n_272), .B(n_333), .Y(n_350) );
INVx1_ASAP7_75t_SL g321 ( .A(n_273), .Y(n_321) );
INVx1_ASAP7_75t_L g348 ( .A(n_274), .Y(n_348) );
AOI31xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .A3(n_279), .B(n_282), .Y(n_276) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g369 ( .A(n_280), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g343 ( .A(n_281), .Y(n_343) );
BUFx2_ASAP7_75t_L g357 ( .A(n_281), .Y(n_357) );
AND2x2_ASAP7_75t_L g385 ( .A(n_281), .B(n_306), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g358 ( .A(n_285), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_286), .B(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g406 ( .A(n_286), .B(n_332), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B(n_295), .C(n_310), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_292), .A2(n_319), .B1(n_320), .B2(n_321), .C(n_322), .Y(n_318) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g326 ( .A(n_293), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g363 ( .A(n_294), .Y(n_363) );
OAI32xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .A3(n_301), .B1(n_303), .B2(n_308), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_297), .A2(n_350), .B(n_351), .C(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_305), .A2(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_312), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g360 ( .A(n_312), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g377 ( .A(n_314), .Y(n_377) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND4xp25_ASAP7_75t_SL g317 ( .A(n_318), .B(n_330), .C(n_349), .D(n_364), .Y(n_317) );
AND2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g378 ( .A(n_319), .B(n_371), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_321), .B(n_353), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_325), .B2(n_328), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_323), .A2(n_374), .B1(n_405), .B2(n_407), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g411 ( .A1(n_323), .A2(n_412), .B(n_413), .C(n_416), .Y(n_411) );
INVx2_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_326), .A2(n_360), .B1(n_377), .B2(n_378), .C1(n_379), .C2(n_382), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_334), .C(n_338), .Y(n_330) );
INVx1_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_335), .A2(n_339), .B1(n_342), .B2(n_344), .Y(n_338) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g365 ( .A(n_347), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g423 ( .A(n_350), .Y(n_423) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_359), .B2(n_362), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_357), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
INVx1_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_368), .Y(n_422) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND5xp2_ASAP7_75t_L g375 ( .A(n_376), .B(n_383), .C(n_397), .D(n_403), .E(n_408), .Y(n_375) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_386), .C(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI31xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .A3(n_393), .B(n_394), .Y(n_389) );
INVx1_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI222xp33_ASAP7_75t_L g418 ( .A1(n_405), .A2(n_407), .B1(n_419), .B2(n_422), .C1(n_423), .C2(n_424), .Y(n_418) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g712 ( .A(n_426), .Y(n_712) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR3x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_614), .C(n_663), .Y(n_428) );
NAND5xp2_ASAP7_75t_L g429 ( .A(n_430), .B(n_548), .C(n_577), .D(n_585), .E(n_600), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_476), .B(n_492), .C(n_532), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_461), .Y(n_431) );
AND2x2_ASAP7_75t_L g543 ( .A(n_432), .B(n_540), .Y(n_543) );
AND2x2_ASAP7_75t_L g576 ( .A(n_432), .B(n_462), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_432), .B(n_480), .Y(n_669) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_449), .Y(n_432) );
INVx2_ASAP7_75t_L g479 ( .A(n_433), .Y(n_479) );
BUFx2_ASAP7_75t_L g643 ( .A(n_433), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .Y(n_434) );
INVx5_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_SL g452 ( .A1(n_443), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_443), .A2(n_454), .B(n_519), .C(n_520), .Y(n_518) );
BUFx2_ASAP7_75t_L g465 ( .A(n_445), .Y(n_465) );
AND2x2_ASAP7_75t_L g461 ( .A(n_449), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
AND2x2_ASAP7_75t_L g627 ( .A(n_449), .B(n_540), .Y(n_627) );
AND2x2_ASAP7_75t_L g682 ( .A(n_449), .B(n_479), .Y(n_682) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_460), .Y(n_449) );
INVx2_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g599 ( .A(n_461), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_461), .B(n_480), .Y(n_646) );
INVx5_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
AND2x4_ASAP7_75t_L g561 ( .A(n_462), .B(n_541), .Y(n_561) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_462), .Y(n_583) );
AND2x2_ASAP7_75t_L g658 ( .A(n_462), .B(n_643), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_462), .B(n_481), .Y(n_661) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_466), .B(n_472), .Y(n_463) );
INVx2_ASAP7_75t_L g471 ( .A(n_469), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_471), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_471), .A2(n_489), .B(n_510), .C(n_511), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_476), .B(n_541), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_476), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
AND2x2_ASAP7_75t_L g566 ( .A(n_478), .B(n_541), .Y(n_566) );
AND2x2_ASAP7_75t_L g584 ( .A(n_478), .B(n_481), .Y(n_584) );
INVx1_ASAP7_75t_L g604 ( .A(n_478), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_478), .B(n_540), .Y(n_649) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_478), .Y(n_691) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_479), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_480), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_480), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_480), .A2(n_536), .B(n_597), .C(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g603 ( .A(n_480), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g612 ( .A(n_480), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g616 ( .A(n_480), .B(n_540), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_480), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g631 ( .A(n_480), .B(n_541), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_480), .B(n_682), .Y(n_681) );
INVx5_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g545 ( .A(n_481), .Y(n_545) );
AND2x2_ASAP7_75t_L g586 ( .A(n_481), .B(n_539), .Y(n_586) );
AND2x2_ASAP7_75t_L g598 ( .A(n_481), .B(n_573), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_481), .B(n_627), .Y(n_645) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_513), .Y(n_492) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
OR2x2_ASAP7_75t_L g536 ( .A(n_494), .B(n_505), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_494), .B(n_543), .C(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_494), .B(n_515), .Y(n_553) );
OR2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_556), .Y(n_568) );
AND2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_524), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_494), .B(n_705), .Y(n_704) );
INVx5_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_495), .B(n_515), .Y(n_571) );
AND2x2_ASAP7_75t_L g610 ( .A(n_495), .B(n_525), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_495), .B(n_524), .Y(n_638) );
OR2x2_ASAP7_75t_L g641 ( .A(n_495), .B(n_524), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_499), .Y(n_496) );
INVx5_ASAP7_75t_SL g556 ( .A(n_505), .Y(n_556) );
OR2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_514), .Y(n_562) );
AND2x2_ASAP7_75t_L g578 ( .A(n_505), .B(n_579), .Y(n_578) );
AOI321xp33_ASAP7_75t_L g585 ( .A1(n_505), .A2(n_586), .A3(n_587), .B1(n_588), .B2(n_594), .C(n_596), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_505), .B(n_513), .Y(n_595) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_505), .Y(n_608) );
OR2x2_ASAP7_75t_L g655 ( .A(n_505), .B(n_553), .Y(n_655) );
AND2x2_ASAP7_75t_L g677 ( .A(n_505), .B(n_574), .Y(n_677) );
AND2x2_ASAP7_75t_L g696 ( .A(n_505), .B(n_515), .Y(n_696) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .Y(n_505) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_515), .B(n_524), .Y(n_537) );
AND2x2_ASAP7_75t_L g546 ( .A(n_515), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g573 ( .A(n_515), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_515), .B(n_574), .Y(n_579) );
INVxp67_ASAP7_75t_L g609 ( .A(n_515), .Y(n_609) );
OR2x2_ASAP7_75t_L g651 ( .A(n_515), .B(n_556), .Y(n_651) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_515) );
OR2x2_ASAP7_75t_L g533 ( .A(n_524), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_SL g547 ( .A(n_524), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_524), .B(n_536), .Y(n_580) );
AND2x2_ASAP7_75t_L g629 ( .A(n_524), .B(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_L g667 ( .A(n_524), .B(n_556), .Y(n_667) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_525), .B(n_556), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B(n_538), .C(n_542), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_533), .A2(n_535), .B1(n_660), .B2(n_662), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_535), .A2(n_558), .B1(n_613), .B2(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_SL g687 ( .A(n_536), .Y(n_687) );
INVx1_ASAP7_75t_SL g587 ( .A(n_537), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_539), .B(n_559), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g600 ( .A1(n_539), .A2(n_580), .B1(n_587), .B2(n_601), .C1(n_605), .C2(n_611), .Y(n_600) );
AND2x2_ASAP7_75t_L g690 ( .A(n_539), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_540), .B(n_560), .Y(n_635) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_540), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_540), .B(n_584), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_540), .B(n_691), .Y(n_701) );
INVx1_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_541), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_543), .A2(n_684), .B(n_685), .C(n_688), .Y(n_683) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_545), .B(n_607), .C(n_610), .Y(n_606) );
OR2x2_ASAP7_75t_L g634 ( .A(n_545), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_545), .B(n_561), .Y(n_662) );
OR2x2_ASAP7_75t_L g567 ( .A(n_547), .B(n_568), .Y(n_567) );
AOI211xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_551), .B(n_557), .C(n_569), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_550), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_552), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g570 ( .A(n_555), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_556), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g624 ( .A(n_556), .B(n_574), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_556), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_556), .B(n_573), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_562), .B1(n_563), .B2(n_567), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_559), .B(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_561), .B(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_SL g625 ( .A1(n_562), .A2(n_626), .B1(n_628), .B2(n_630), .C(n_632), .Y(n_625) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g680 ( .A(n_565), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_565), .B(n_682), .Y(n_693) );
INVx1_ASAP7_75t_L g613 ( .A(n_566), .Y(n_613) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_568), .A2(n_651), .B(n_674), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B(n_575), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g617 ( .A(n_578), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_579), .A2(n_665), .B1(n_668), .B2(n_670), .C(n_673), .Y(n_664) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_587), .A2(n_677), .B1(n_678), .B2(n_680), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g653 ( .A(n_589), .Y(n_653) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp67_ASAP7_75t_SL g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g657 ( .A(n_593), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g622 ( .A(n_598), .Y(n_622) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_603), .B(n_627), .Y(n_679) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_609), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_610), .B(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g702 ( .A(n_610), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI211xp5_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_617), .B(n_618), .C(n_652), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_625), .C(n_644), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g705 ( .A(n_629), .Y(n_705) );
AND2x2_ASAP7_75t_L g642 ( .A(n_631), .B(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_640), .B2(n_642), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g650 ( .A(n_638), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g703 ( .A(n_639), .Y(n_703) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI31xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .A3(n_647), .B(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_659), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_676), .C(n_683), .D(n_697), .E(n_700), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_675), .A2(n_701), .B1(n_702), .B2(n_704), .Y(n_700) );
INVx1_ASAP7_75t_SL g699 ( .A(n_677), .Y(n_699) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_692), .B(n_694), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g713 ( .A(n_706), .Y(n_713) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g731 ( .A(n_719), .Y(n_731) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g735 ( .A(n_724), .Y(n_735) );
INVx1_ASAP7_75t_L g729 ( .A(n_727), .Y(n_729) );
BUFx3_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
endmodule