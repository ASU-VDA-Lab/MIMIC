module fake_jpeg_28327_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_45),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_22),
.B1(n_29),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_32),
.B1(n_19),
.B2(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_22),
.B1(n_17),
.B2(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_71),
.B1(n_18),
.B2(n_20),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_22),
.B1(n_29),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_58),
.B1(n_32),
.B2(n_20),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_27),
.B1(n_36),
.B2(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_73),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_21),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_30),
.B(n_23),
.C(n_28),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_34),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_17),
.B1(n_19),
.B2(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_34),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_33),
.B1(n_32),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_89),
.B1(n_110),
.B2(n_114),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_97),
.B(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_105),
.B1(n_115),
.B2(n_50),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_87),
.B1(n_93),
.B2(n_108),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_20),
.B1(n_18),
.B2(n_26),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_92),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_53),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_107),
.B(n_30),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_26),
.B1(n_11),
.B2(n_16),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_100),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_23),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_25),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_54),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_49),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_49),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_52),
.A2(n_25),
.B1(n_30),
.B2(n_16),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_113),
.Y(n_143)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_56),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_30),
.B1(n_15),
.B2(n_13),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_118),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_68),
.B1(n_50),
.B2(n_48),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_123),
.B1(n_127),
.B2(n_93),
.Y(n_148)
);

NOR2x1_ASAP7_75t_R g121 ( 
.A(n_91),
.B(n_54),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_128),
.B(n_140),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_81),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_79),
.A2(n_74),
.B1(n_63),
.B2(n_59),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_0),
.B(n_2),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_63),
.B1(n_69),
.B2(n_76),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_113),
.B1(n_105),
.B2(n_76),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_76),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_129),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_2),
.B(n_3),
.Y(n_179)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_99),
.B1(n_113),
.B2(n_78),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_103),
.C(n_96),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_144),
.C(n_122),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_152),
.B1(n_162),
.B2(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_88),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_111),
.B(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_172),
.B(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_88),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_90),
.B1(n_84),
.B2(n_89),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_165),
.B1(n_173),
.B2(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_159),
.B(n_164),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_87),
.B1(n_86),
.B2(n_107),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_118),
.A2(n_95),
.B1(n_100),
.B2(n_81),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_145),
.C(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_107),
.B1(n_97),
.B2(n_111),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_138),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_104),
.A3(n_97),
.B1(n_107),
.B2(n_88),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_101),
.B1(n_80),
.B2(n_112),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_106),
.B1(n_97),
.B2(n_108),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_78),
.B1(n_115),
.B2(n_102),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_120),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_123),
.A2(n_101),
.B1(n_62),
.B2(n_15),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_121),
.B1(n_139),
.B2(n_126),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_140),
.B(n_138),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_140),
.B(n_128),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_181),
.B(n_192),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_207),
.B1(n_174),
.B2(n_160),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_185),
.A2(n_186),
.B1(n_199),
.B2(n_209),
.Y(n_237)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_140),
.C(n_138),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_195),
.C(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_193),
.B(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_137),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_177),
.C(n_170),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_145),
.B1(n_117),
.B2(n_130),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

CKINVDCx6p67_ASAP7_75t_R g197 ( 
.A(n_152),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_149),
.B(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_120),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_13),
.B1(n_12),
.B2(n_6),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_13),
.B1(n_12),
.B2(n_6),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_176),
.B1(n_175),
.B2(n_148),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_224),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_163),
.C(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_163),
.C(n_155),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_190),
.C(n_180),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_197),
.B1(n_188),
.B2(n_8),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_155),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_182),
.B(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_171),
.C(n_179),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_231),
.C(n_233),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_168),
.C(n_161),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_172),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_161),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_235),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_3),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_4),
.C(n_6),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_238),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

AOI321xp33_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_201),
.A3(n_184),
.B1(n_185),
.B2(n_183),
.C(n_200),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_248),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_252),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_210),
.B(n_202),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_208),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_258),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_197),
.B1(n_205),
.B2(n_206),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_257),
.B1(n_227),
.B2(n_222),
.Y(n_272)
);

OAI322xp33_ASAP7_75t_L g256 ( 
.A1(n_212),
.A2(n_191),
.A3(n_204),
.B1(n_187),
.B2(n_209),
.C1(n_211),
.C2(n_197),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_245),
.C(n_242),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_260),
.A2(n_216),
.B1(n_213),
.B2(n_229),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_259),
.A2(n_223),
.B(n_224),
.Y(n_264)
);

OAI21x1_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_273),
.B(n_239),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_267),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_270),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_225),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_236),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_275),
.C(n_242),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_259),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_4),
.C(n_7),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_4),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_277),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_243),
.A2(n_9),
.B1(n_10),
.B2(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_246),
.Y(n_289)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_248),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_255),
.B1(n_244),
.B2(n_257),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_263),
.B(n_264),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_284),
.B(n_253),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_292),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_260),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_287),
.B(n_266),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_247),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_271),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_273),
.B(n_249),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.C(n_304),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_281),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_252),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_284),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_240),
.B(n_270),
.Y(n_301)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_9),
.B1(n_10),
.B2(n_240),
.C(n_293),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_R g307 ( 
.A(n_305),
.B(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_294),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_313),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_288),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_288),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_286),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_302),
.B(n_303),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_312),
.B(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_279),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_319),
.B(n_320),
.C(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_292),
.Y(n_321)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_324),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_325),
.C(n_318),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_326),
.Y(n_329)
);


endmodule