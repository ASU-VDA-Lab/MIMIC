module fake_jpeg_30444_n_282 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_220;
wire n_137;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_1),
.Y(n_75)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_35),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_38),
.B1(n_18),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_61),
.B1(n_64),
.B2(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_22),
.B1(n_36),
.B2(n_34),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_57),
.A2(n_70),
.B(n_86),
.Y(n_116)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_31),
.B1(n_35),
.B2(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_62),
.B(n_63),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_35),
.B1(n_26),
.B2(n_37),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_26),
.B1(n_36),
.B2(n_34),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_52),
.B1(n_41),
.B2(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_83),
.B1(n_46),
.B2(n_21),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_53),
.B1(n_47),
.B2(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_72),
.B1(n_67),
.B2(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_71),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_47),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_21),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_21),
.B1(n_24),
.B2(n_19),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_66),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_70),
.C(n_87),
.Y(n_145)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_91),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_53),
.B1(n_44),
.B2(n_21),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_102),
.B1(n_104),
.B2(n_108),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_44),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_95),
.Y(n_134)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_56),
.B(n_86),
.Y(n_130)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_81),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_59),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_118),
.B1(n_60),
.B2(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_8),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_70),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_118)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_56),
.Y(n_125)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_128),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_143),
.B(n_113),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_142),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_70),
.B(n_87),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_148),
.B(n_90),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_81),
.B(n_69),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_146),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_91),
.C(n_88),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_89),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_94),
.B(n_80),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_93),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_56),
.B(n_78),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_56),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_99),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_117),
.B1(n_104),
.B2(n_102),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_156),
.B1(n_177),
.B2(n_138),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_172),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_89),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_99),
.B(n_103),
.C(n_98),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_97),
.B1(n_105),
.B2(n_78),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_106),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_97),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_175),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_96),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_178),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_112),
.B1(n_120),
.B2(n_105),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_101),
.B(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_126),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

NAND4xp25_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_191),
.C(n_192),
.D(n_155),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_168),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_172),
.B1(n_154),
.B2(n_166),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_189),
.B1(n_196),
.B2(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_130),
.B1(n_134),
.B2(n_146),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_141),
.C(n_147),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_134),
.A3(n_138),
.B1(n_147),
.B2(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_147),
.B1(n_131),
.B2(n_123),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_139),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_180),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_131),
.B1(n_123),
.B2(n_136),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_187),
.C(n_186),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_213),
.C(n_215),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_133),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_160),
.B1(n_155),
.B2(n_179),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_222),
.B1(n_223),
.B2(n_200),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_220),
.B(n_221),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_178),
.C(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_133),
.Y(n_218)
);

OAI322xp33_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_163),
.A3(n_161),
.B1(n_153),
.B2(n_177),
.C1(n_164),
.C2(n_157),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_219),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_161),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_181),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_199),
.C(n_196),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.C(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_231),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_204),
.C(n_181),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_201),
.C(n_192),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_192),
.B(n_195),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_220),
.B(n_222),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_203),
.C(n_198),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_195),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_205),
.C(n_217),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_248),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_228),
.B(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_245),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_223),
.B1(n_221),
.B2(n_208),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_246),
.B1(n_250),
.B2(n_162),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_208),
.B1(n_214),
.B2(n_216),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_193),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_203),
.C(n_198),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_235),
.C(n_227),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_255),
.C(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_229),
.C(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_193),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_258),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_157),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_123),
.C(n_88),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_240),
.B1(n_244),
.B2(n_239),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_264),
.Y(n_270)
);

AND3x1_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_137),
.C(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_171),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_169),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_136),
.B1(n_137),
.B2(n_119),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_255),
.B(n_257),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_268),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_260),
.C(n_261),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_270),
.C(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_15),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.C(n_276),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_278),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_270),
.Y(n_282)
);


endmodule