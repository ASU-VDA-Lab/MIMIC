module fake_netlist_6_2911_n_1830 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1830);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1830;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_934;
wire n_482;
wire n_204;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_48),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_27),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_89),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_25),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_40),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_70),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_73),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_80),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_126),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_100),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_51),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_19),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_29),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_21),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_42),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_68),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_115),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_45),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_37),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_51),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_147),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_24),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_16),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_2),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_39),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_34),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_53),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_49),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_26),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_47),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_139),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_65),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_95),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_140),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_4),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_125),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_82),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_63),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_32),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_49),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_34),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_48),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_12),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_83),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_129),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_36),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_67),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_52),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_93),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_62),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_78),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_103),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_13),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_26),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_88),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_54),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_46),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_43),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_157),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_86),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_79),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_52),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_87),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_99),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_110),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_17),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_104),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_84),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_106),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_38),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_20),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_161),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_141),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_53),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_156),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_5),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_54),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_76),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_127),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_6),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_40),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_60),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_109),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_11),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_143),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_153),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_92),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_111),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_101),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_61),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_158),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_23),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_41),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_91),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_145),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_4),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_22),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_28),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_15),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_120),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_98),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_112),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_14),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_21),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_59),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_36),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_61),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_9),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_108),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_155),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_28),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_60),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_46),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_45),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_55),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_31),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_19),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_102),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_192),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_174),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_174),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_176),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_169),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_205),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_176),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_189),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_182),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_189),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_264),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_227),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_201),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_277),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_272),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_183),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_186),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_227),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_227),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_267),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_188),
.Y(n_351)
);

INVx4_ASAP7_75t_R g352 ( 
.A(n_277),
.Y(n_352)
);

BUFx2_ASAP7_75t_SL g353 ( 
.A(n_224),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_166),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_320),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_190),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_201),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_208),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_208),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_165),
.B(n_184),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_224),
.B(n_0),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_193),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_168),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_267),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_209),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_257),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_170),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_209),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_216),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_216),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_227),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_225),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_225),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_231),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_165),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_196),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_171),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_172),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_197),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_203),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_175),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_231),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_239),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_239),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_267),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_245),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_234),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_245),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_250),
.B(n_1),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_227),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_215),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_259),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_177),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_217),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_228),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_237),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_251),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_241),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_241),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_241),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_252),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_250),
.B(n_1),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_241),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_262),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_341),
.A2(n_270),
.B(n_206),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_259),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_361),
.B(n_234),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_173),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_173),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_349),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_387),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_371),
.A2(n_211),
.B(n_194),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_241),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_289),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_402),
.B(n_234),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_343),
.B(n_326),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_270),
.B(n_206),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_289),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_332),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_337),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_357),
.B(n_289),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_365),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_369),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_370),
.B(n_289),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_374),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_384),
.B(n_289),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_360),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_353),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_329),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_352),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_329),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_334),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_334),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_328),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_338),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_338),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_406),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_194),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_345),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_419),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_R g484 ( 
.A(n_410),
.B(n_345),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_475),
.B(n_350),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

BUFx4f_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_477),
.A2(n_471),
.B1(n_478),
.B2(n_474),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_420),
.B(n_364),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_420),
.Y(n_491)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_346),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_420),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

OAI22xp33_ASAP7_75t_L g498 ( 
.A1(n_475),
.A2(n_232),
.B1(n_355),
.B2(n_311),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_476),
.A2(n_300),
.B1(n_323),
.B2(n_293),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_410),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_296),
.B1(n_279),
.B2(n_325),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_268),
.C(n_261),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_466),
.B(n_346),
.Y(n_507)
);

INVxp33_ASAP7_75t_SL g508 ( 
.A(n_422),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_211),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_466),
.B(n_351),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_475),
.B(n_351),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_466),
.B(n_356),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_466),
.A2(n_296),
.B1(n_279),
.B2(n_325),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_441),
.Y(n_517)
);

NOR2x1p5_ASAP7_75t_L g518 ( 
.A(n_475),
.B(n_473),
.Y(n_518)
);

INVx8_ASAP7_75t_L g519 ( 
.A(n_466),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_410),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_406),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_410),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_406),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_445),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_470),
.B(n_356),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_471),
.B(n_261),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_444),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

BUFx12f_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_470),
.B(n_362),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_268),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_445),
.B(n_362),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_470),
.B(n_376),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_445),
.B(n_376),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_385),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_437),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_470),
.B(n_379),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_437),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_447),
.B(n_379),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_391),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_444),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_447),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_430),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_471),
.B(n_276),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_467),
.B(n_391),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_433),
.A2(n_296),
.B1(n_214),
.B2(n_220),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_448),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_437),
.Y(n_563)
);

AO21x2_ASAP7_75t_L g564 ( 
.A1(n_417),
.A2(n_282),
.B(n_276),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_446),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_411),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_419),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_467),
.B(n_468),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_419),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_430),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_468),
.B(n_395),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_419),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_468),
.B(n_395),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_471),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_477),
.B(n_396),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_446),
.Y(n_579)
);

AOI21x1_ASAP7_75t_L g580 ( 
.A1(n_417),
.A2(n_284),
.B(n_282),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_476),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_477),
.B(n_396),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_419),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_430),
.Y(n_584)
);

CKINVDCx11_ASAP7_75t_R g585 ( 
.A(n_411),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_433),
.B(n_397),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_423),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_477),
.B(n_397),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_430),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_433),
.A2(n_296),
.B1(n_214),
.B2(n_220),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_474),
.B(n_473),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_446),
.Y(n_593)
);

BUFx4f_ASAP7_75t_L g594 ( 
.A(n_474),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_449),
.B(n_401),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_453),
.B(n_401),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_453),
.B(n_404),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_452),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_453),
.B(n_404),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_443),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_417),
.A2(n_296),
.B1(n_210),
.B2(n_302),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_423),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_452),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_478),
.B(n_354),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_423),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_476),
.A2(n_316),
.B1(n_266),
.B2(n_271),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_449),
.B(n_363),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_416),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_423),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_478),
.B(n_393),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_416),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_423),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_423),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_423),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_416),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_452),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_423),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_451),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_448),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_453),
.B(n_244),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_461),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_434),
.B(n_288),
.C(n_284),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_416),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_473),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_620),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_576),
.B(n_474),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_481),
.A2(n_474),
.B1(n_473),
.B2(n_469),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_576),
.B(n_474),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_564),
.A2(n_434),
.B1(n_474),
.B2(n_473),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_624),
.B(n_473),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_481),
.B(n_473),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_564),
.A2(n_434),
.B1(n_473),
.B2(n_460),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_577),
.B(n_367),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_488),
.B(n_594),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_488),
.B(n_411),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_568),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_558),
.B(n_377),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_568),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_569),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_562),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g644 ( 
.A(n_490),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_564),
.A2(n_493),
.B1(n_624),
.B2(n_528),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_569),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_493),
.A2(n_472),
.B1(n_469),
.B2(n_381),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_528),
.A2(n_460),
.B1(n_448),
.B2(n_436),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_571),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_508),
.B(n_378),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_507),
.B(n_453),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_SL g652 ( 
.A(n_491),
.B(n_340),
.C(n_335),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_533),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_512),
.B(n_448),
.Y(n_654)
);

NAND2x1_ASAP7_75t_L g655 ( 
.A(n_483),
.B(n_416),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_508),
.B(n_344),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_533),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_514),
.B(n_448),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_587),
.B(n_347),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_519),
.B(n_234),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_570),
.B(n_554),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_489),
.A2(n_472),
.B1(n_469),
.B2(n_330),
.Y(n_663)
);

NAND2x1_ASAP7_75t_L g664 ( 
.A(n_483),
.B(n_504),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_623),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_494),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_490),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_552),
.B(n_539),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_479),
.Y(n_669)
);

BUFx4f_ASAP7_75t_L g670 ( 
.A(n_531),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_581),
.B(n_460),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_594),
.B(n_469),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_486),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_573),
.A2(n_472),
.B1(n_409),
.B2(n_436),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_486),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_581),
.B(n_622),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_552),
.B(n_472),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_499),
.A2(n_273),
.B1(n_274),
.B2(n_278),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_603),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_495),
.A2(n_460),
.B1(n_436),
.B2(n_409),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_483),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_519),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_586),
.B(n_409),
.Y(n_683)
);

AND2x2_ASAP7_75t_SL g684 ( 
.A(n_602),
.B(n_212),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_491),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_574),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_495),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_542),
.B(n_409),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_586),
.B(n_436),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_603),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_574),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_543),
.B(n_234),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_497),
.A2(n_297),
.B(n_185),
.C(n_200),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_544),
.B(n_461),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_531),
.A2(n_557),
.B1(n_538),
.B2(n_551),
.Y(n_695)
);

AND2x6_ASAP7_75t_SL g696 ( 
.A(n_550),
.B(n_184),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_519),
.A2(n_408),
.B(n_405),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_575),
.A2(n_260),
.B1(n_269),
.B2(n_460),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_497),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_583),
.B(n_442),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_583),
.B(n_442),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_588),
.B(n_442),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_588),
.B(n_442),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_603),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_543),
.B(n_443),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_610),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_L g707 ( 
.A(n_500),
.B(n_461),
.C(n_457),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_610),
.B(n_442),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_597),
.B(n_451),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_521),
.B(n_524),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_502),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_502),
.A2(n_442),
.B1(n_246),
.B2(n_263),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_613),
.B(n_442),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_613),
.B(n_442),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_562),
.B(n_621),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_598),
.B(n_451),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_621),
.B(n_288),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_600),
.B(n_578),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_615),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_505),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_518),
.A2(n_212),
.B1(n_263),
.B2(n_246),
.Y(n_722)
);

BUFx8_ASAP7_75t_L g723 ( 
.A(n_534),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_505),
.A2(n_200),
.B(n_210),
.C(n_303),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_534),
.B(n_457),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_615),
.B(n_405),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_619),
.B(n_405),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_603),
.B(n_443),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_619),
.B(n_405),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_567),
.B(n_457),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_522),
.B(n_405),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_522),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_603),
.B(n_443),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_519),
.B(n_317),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_499),
.A2(n_283),
.B1(n_286),
.B2(n_295),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_525),
.B(n_408),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_525),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_606),
.B(n_443),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_529),
.Y(n_739)
);

BUFx6f_ASAP7_75t_SL g740 ( 
.A(n_531),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_609),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_519),
.B(n_317),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_529),
.B(n_408),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_545),
.B(n_408),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_606),
.B(n_443),
.Y(n_745)
);

AOI221xp5_ASAP7_75t_L g746 ( 
.A1(n_498),
.A2(n_280),
.B1(n_213),
.B2(n_253),
.C(n_275),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_545),
.B(n_408),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_547),
.B(n_548),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_582),
.B(n_457),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_606),
.B(n_623),
.Y(n_750)
);

NAND2x1_ASAP7_75t_L g751 ( 
.A(n_483),
.B(n_416),
.Y(n_751)
);

BUFx5_ASAP7_75t_L g752 ( 
.A(n_547),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_548),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_609),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_549),
.B(n_412),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_549),
.B(n_563),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_563),
.B(n_412),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_606),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_537),
.B(n_458),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_565),
.B(n_412),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_565),
.B(n_412),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_482),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_484),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_500),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_623),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_L g766 ( 
.A(n_480),
.B(n_510),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_518),
.B(n_412),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_503),
.A2(n_465),
.B1(n_454),
.B2(n_463),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_537),
.B(n_596),
.Y(n_769)
);

NAND2x1_ASAP7_75t_L g770 ( 
.A(n_504),
.B(n_416),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_609),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_482),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_606),
.B(n_443),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_623),
.B(n_443),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_612),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_589),
.B(n_513),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_612),
.Y(n_778)
);

O2A1O1Ixp5_ASAP7_75t_L g779 ( 
.A1(n_580),
.A2(n_465),
.B(n_463),
.C(n_454),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_485),
.B(n_458),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_504),
.B(n_443),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_496),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_530),
.B(n_458),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_504),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_616),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_616),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_496),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_616),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_516),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_531),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_531),
.B(n_414),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_509),
.B(n_443),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_608),
.B(n_458),
.C(n_310),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_688),
.B(n_668),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_692),
.A2(n_705),
.B(n_781),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_710),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_715),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_666),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_670),
.B(n_684),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_709),
.B(n_538),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_679),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_681),
.A2(n_614),
.B(n_509),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_769),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_681),
.A2(n_614),
.B(n_509),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_784),
.B(n_752),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_677),
.B(n_763),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_720),
.B(n_611),
.Y(n_807)
);

AOI21x1_ASAP7_75t_L g808 ( 
.A1(n_692),
.A2(n_580),
.B(n_517),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_748),
.A2(n_592),
.B(n_503),
.Y(n_809)
);

BUFx4f_ASAP7_75t_L g810 ( 
.A(n_694),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_716),
.B(n_538),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_718),
.A2(n_607),
.B(n_540),
.C(n_546),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_777),
.A2(n_535),
.B1(n_614),
.B2(n_557),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_756),
.A2(n_592),
.B(n_510),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_784),
.A2(n_592),
.B(n_418),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_731),
.A2(n_592),
.B(n_510),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_659),
.A2(n_557),
.B1(n_538),
.B2(n_592),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_627),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_676),
.B(n_538),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_764),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_662),
.B(n_557),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_784),
.A2(n_418),
.B(n_414),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_752),
.B(n_557),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_752),
.B(n_625),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_723),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_638),
.A2(n_456),
.B(n_462),
.C(n_450),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_640),
.A2(n_510),
.B1(n_480),
.B2(n_625),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_682),
.A2(n_418),
.B(n_414),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_682),
.A2(n_661),
.B(n_697),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_752),
.B(n_625),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_638),
.A2(n_480),
.B1(n_510),
.B2(n_607),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_682),
.A2(n_418),
.B(n_414),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_730),
.A2(n_591),
.B(n_561),
.Y(n_833)
);

HAxp5_ASAP7_75t_L g834 ( 
.A(n_678),
.B(n_202),
.CON(n_834),
.SN(n_834)
);

INVx11_ASAP7_75t_L g835 ( 
.A(n_723),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_752),
.B(n_506),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_764),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_752),
.B(n_506),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_752),
.B(n_533),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_684),
.A2(n_515),
.B1(n_501),
.B2(n_510),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_695),
.A2(n_301),
.B(n_290),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_633),
.B(n_506),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_661),
.A2(n_418),
.B(n_414),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_723),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_633),
.B(n_511),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_734),
.A2(n_424),
.B(n_421),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_734),
.A2(n_424),
.B(n_421),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_742),
.A2(n_424),
.B(n_421),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_669),
.A2(n_480),
.B1(n_510),
.B2(n_280),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_644),
.B(n_636),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_679),
.B(n_533),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_742),
.A2(n_424),
.B(n_421),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_783),
.A2(n_672),
.B1(n_749),
.B2(n_629),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_685),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_736),
.A2(n_480),
.B(n_431),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_743),
.A2(n_424),
.B(n_421),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_669),
.B(n_511),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_744),
.A2(n_425),
.B(n_533),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_683),
.B(n_585),
.Y(n_859)
);

OAI321xp33_ASAP7_75t_L g860 ( 
.A1(n_746),
.A2(n_235),
.A3(n_230),
.B1(n_229),
.B2(n_243),
.C(n_223),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_693),
.A2(n_462),
.B(n_450),
.C(n_456),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_673),
.B(n_511),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_679),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_672),
.A2(n_480),
.B1(n_254),
.B2(n_238),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_747),
.A2(n_480),
.B(n_431),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_673),
.B(n_527),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_679),
.B(n_536),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_675),
.B(n_527),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_626),
.A2(n_255),
.B1(n_179),
.B2(n_180),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_650),
.B(n_450),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_645),
.A2(n_631),
.B1(n_670),
.B2(n_634),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_755),
.A2(n_431),
.B(n_516),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_690),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_644),
.B(n_527),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_689),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_759),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_639),
.A2(n_290),
.B(n_301),
.C(n_307),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_715),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_675),
.B(n_555),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_687),
.A2(n_249),
.B(n_185),
.C(n_213),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_757),
.A2(n_761),
.B(n_760),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_667),
.B(n_555),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_690),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_690),
.B(n_536),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_690),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_670),
.A2(n_326),
.B1(n_318),
.B2(n_308),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_641),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_687),
.B(n_555),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_699),
.B(n_556),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_637),
.A2(n_425),
.B(n_536),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_L g891 ( 
.A1(n_647),
.A2(n_312),
.B(n_304),
.Y(n_891)
);

AND2x6_ASAP7_75t_L g892 ( 
.A(n_699),
.B(n_536),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_711),
.A2(n_248),
.B(n_223),
.C(n_229),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_762),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_711),
.B(n_556),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_790),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_721),
.B(n_732),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_721),
.B(n_556),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_637),
.A2(n_425),
.B(n_536),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_767),
.A2(n_431),
.B(n_517),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_722),
.A2(n_618),
.B(n_617),
.C(n_604),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_715),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_705),
.A2(n_523),
.B(n_520),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_732),
.B(n_584),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_762),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_628),
.A2(n_425),
.B(n_572),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_630),
.A2(n_425),
.B(n_572),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_791),
.A2(n_431),
.B(n_520),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_653),
.A2(n_572),
.B(n_492),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_SL g910 ( 
.A(n_656),
.B(n_178),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_654),
.A2(n_526),
.B(n_523),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_658),
.A2(n_532),
.B(n_526),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_704),
.B(n_572),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_643),
.B(n_307),
.Y(n_914)
);

OAI21xp33_ASAP7_75t_L g915 ( 
.A1(n_663),
.A2(n_319),
.B(n_314),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_651),
.A2(n_318),
.B(n_308),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_657),
.A2(n_572),
.B(n_492),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_704),
.B(n_584),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_693),
.A2(n_456),
.B(n_462),
.C(n_439),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_773),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_737),
.B(n_584),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_724),
.A2(n_432),
.B(n_439),
.C(n_604),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_642),
.A2(n_618),
.B(n_617),
.C(n_599),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_704),
.B(n_532),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_696),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_737),
.B(n_739),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_773),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_643),
.B(n_230),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_646),
.A2(n_560),
.B(n_599),
.C(n_595),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_704),
.B(n_541),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_664),
.A2(n_492),
.B(n_487),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_726),
.A2(n_492),
.B(n_487),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_727),
.A2(n_590),
.B(n_487),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_780),
.B(n_321),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_717),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_739),
.B(n_541),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_782),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_793),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_729),
.A2(n_750),
.B(n_781),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_790),
.A2(n_236),
.B1(n_265),
.B2(n_256),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_750),
.A2(n_248),
.B(n_235),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_792),
.A2(n_487),
.B(n_590),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_782),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_753),
.B(n_553),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_753),
.B(n_553),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_758),
.B(n_559),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_717),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_674),
.B(n_322),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_717),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_652),
.B(n_324),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_758),
.B(n_559),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_792),
.A2(n_590),
.B(n_595),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_787),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_671),
.A2(n_590),
.B(n_593),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_758),
.B(n_560),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_665),
.B(n_566),
.Y(n_956)
);

O2A1O1Ixp5_ASAP7_75t_L g957 ( 
.A1(n_775),
.A2(n_593),
.B(n_579),
.C(n_566),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_758),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_649),
.A2(n_455),
.B(n_465),
.C(n_459),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_660),
.B(n_455),
.Y(n_960)
);

CKINVDCx10_ASAP7_75t_R g961 ( 
.A(n_740),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_700),
.A2(n_455),
.B(n_465),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_686),
.B(n_455),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_701),
.A2(n_590),
.B(n_601),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_787),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_691),
.B(n_455),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_706),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_719),
.A2(n_459),
.B(n_465),
.C(n_463),
.Y(n_968)
);

OAI321xp33_ASAP7_75t_L g969 ( 
.A1(n_735),
.A2(n_309),
.A3(n_243),
.B1(n_249),
.B2(n_315),
.C(n_253),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_665),
.B(n_459),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_765),
.B(n_443),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_712),
.A2(n_299),
.B1(n_187),
.B2(n_191),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_775),
.A2(n_313),
.B(n_315),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_853),
.A2(n_632),
.B(n_725),
.C(n_698),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_801),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_798),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_810),
.B(n_765),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_812),
.A2(n_707),
.B(n_714),
.C(n_703),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_829),
.A2(n_766),
.B(n_680),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_794),
.B(n_806),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_796),
.B(n_648),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_806),
.B(n_741),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_810),
.B(n_635),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_818),
.Y(n_984)
);

OA22x2_ASAP7_75t_L g985 ( 
.A1(n_876),
.A2(n_302),
.B1(n_297),
.B2(n_303),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_825),
.B(n_702),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_805),
.A2(n_766),
.B(n_751),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_870),
.B(n_754),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_971),
.A2(n_713),
.B(n_708),
.C(n_738),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_798),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_796),
.B(n_202),
.Y(n_991)
);

AOI33xp33_ASAP7_75t_L g992 ( 
.A1(n_859),
.A2(n_305),
.A3(n_313),
.B1(n_285),
.B2(n_281),
.B3(n_275),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_L g993 ( 
.A(n_948),
.B(n_771),
.C(n_788),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_850),
.B(n_807),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_875),
.B(n_202),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_854),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_799),
.A2(n_740),
.B1(n_258),
.B2(n_281),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_799),
.A2(n_740),
.B1(n_786),
.B2(n_785),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_948),
.A2(n_778),
.B(n_776),
.C(n_772),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_841),
.A2(n_305),
.B1(n_258),
.B2(n_285),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_SL g1001 ( 
.A1(n_925),
.A2(n_291),
.B1(n_309),
.B2(n_242),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_934),
.B(n_789),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_934),
.B(n_789),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_887),
.B(n_728),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_SL g1005 ( 
.A(n_910),
.B(n_306),
.C(n_181),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_808),
.A2(n_745),
.B(n_774),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_800),
.A2(n_745),
.B1(n_774),
.B2(n_733),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_805),
.A2(n_770),
.B(n_655),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_881),
.A2(n_738),
.B(n_733),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_SL g1010 ( 
.A1(n_820),
.A2(n_291),
.B1(n_222),
.B2(n_221),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_850),
.B(n_728),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_801),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_967),
.B(n_459),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_833),
.A2(n_202),
.B1(n_178),
.B2(n_219),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_807),
.A2(n_779),
.B(n_768),
.C(n_459),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_938),
.B(n_195),
.Y(n_1016)
);

NOR2xp67_ASAP7_75t_R g1017 ( 
.A(n_935),
.B(n_463),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_894),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_SL g1019 ( 
.A1(n_941),
.A2(n_432),
.B(n_463),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_803),
.B(n_875),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_823),
.A2(n_590),
.B(n_601),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_SL g1022 ( 
.A(n_950),
.B(n_915),
.C(n_891),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_835),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_811),
.A2(n_294),
.B1(n_218),
.B2(n_199),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_815),
.A2(n_601),
.B(n_416),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_813),
.A2(n_207),
.B(n_226),
.C(n_233),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_874),
.B(n_413),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_905),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_947),
.B(n_198),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_SL g1030 ( 
.A(n_950),
.B(n_292),
.C(n_287),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_SL g1031 ( 
.A(n_817),
.B(n_247),
.C(n_240),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_928),
.B(n_178),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_928),
.B(n_204),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_874),
.B(n_413),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_834),
.A2(n_440),
.B(n_415),
.C(n_413),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_882),
.B(n_415),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_920),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_939),
.A2(n_428),
.B(n_427),
.C(n_407),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_871),
.A2(n_464),
.B1(n_443),
.B2(n_428),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_797),
.B(n_204),
.Y(n_1040)
);

CKINVDCx8_ASAP7_75t_R g1041 ( 
.A(n_961),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_927),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_834),
.A2(n_440),
.B(n_415),
.C(n_407),
.Y(n_1043)
);

AO22x1_ASAP7_75t_L g1044 ( 
.A1(n_837),
.A2(n_204),
.B1(n_219),
.B2(n_440),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_882),
.B(n_428),
.Y(n_1045)
);

BUFx8_ASAP7_75t_L g1046 ( 
.A(n_914),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_802),
.A2(n_804),
.B(n_824),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_937),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_914),
.Y(n_1049)
);

BUFx8_ASAP7_75t_SL g1050 ( 
.A(n_844),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_830),
.A2(n_601),
.B(n_426),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_896),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_814),
.A2(n_428),
.B(n_407),
.C(n_438),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_969),
.B(n_860),
.C(n_886),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_896),
.B(n_2),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_943),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_949),
.A2(n_219),
.B1(n_464),
.B2(n_438),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_SL g1058 ( 
.A(n_940),
.B(n_916),
.C(n_869),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_464),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_953),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_801),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_836),
.A2(n_601),
.B(n_426),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_821),
.B(n_438),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_965),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_797),
.B(n_163),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_878),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_819),
.B(n_438),
.C(n_429),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_809),
.A2(n_464),
.B1(n_429),
.B2(n_427),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_878),
.A2(n_464),
.B1(n_429),
.B2(n_427),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_902),
.B(n_429),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_902),
.Y(n_1071)
);

BUFx4f_ASAP7_75t_L g1072 ( 
.A(n_801),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_936),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_897),
.B(n_427),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_944),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_945),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_926),
.B(n_407),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_863),
.B(n_3),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_873),
.B(n_162),
.Y(n_1079)
);

INVx5_ASAP7_75t_L g1080 ( 
.A(n_873),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_960),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_873),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_863),
.B(n_5),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_880),
.A2(n_435),
.B(n_426),
.C(n_10),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_963),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_827),
.A2(n_464),
.B1(n_426),
.B2(n_435),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_966),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_972),
.A2(n_831),
.B1(n_864),
.B2(n_971),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_826),
.A2(n_464),
.B(n_426),
.C(n_435),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_956),
.B(n_464),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_959),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_816),
.A2(n_464),
.B(n_426),
.C(n_435),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_968),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_883),
.B(n_7),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_956),
.B(n_464),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_873),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_885),
.B(n_150),
.Y(n_1097)
);

AND2x2_ASAP7_75t_SL g1098 ( 
.A(n_840),
.B(n_885),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_840),
.A2(n_464),
.B1(n_435),
.B2(n_426),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_838),
.A2(n_464),
.B(n_144),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_903),
.A2(n_142),
.B(n_137),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_795),
.A2(n_136),
.B1(n_134),
.B2(n_131),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_885),
.B(n_7),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_880),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_883),
.B(n_8),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_923),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_929),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_839),
.A2(n_858),
.B(n_828),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_885),
.B(n_128),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_L g1110 ( 
.A1(n_893),
.A2(n_12),
.B(n_14),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_893),
.A2(n_877),
.B1(n_861),
.B2(n_919),
.C(n_922),
.Y(n_1111)
);

INVxp33_ASAP7_75t_SL g1112 ( 
.A(n_970),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_842),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_973),
.A2(n_116),
.B1(n_113),
.B2(n_97),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_958),
.B(n_90),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_924),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_892),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_855),
.A2(n_865),
.B(n_908),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_845),
.B(n_18),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_849),
.B(n_85),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_849),
.A2(n_22),
.B(n_25),
.Y(n_1121)
);

BUFx8_ASAP7_75t_L g1122 ( 
.A(n_976),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_990),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1022),
.A2(n_994),
.B1(n_1112),
.B2(n_1005),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_979),
.A2(n_974),
.B(n_1002),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_980),
.A2(n_839),
.B1(n_851),
.B2(n_889),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_996),
.B(n_851),
.Y(n_1127)
);

OAI22x1_ASAP7_75t_L g1128 ( 
.A1(n_1055),
.A2(n_913),
.B1(n_884),
.B2(n_867),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_978),
.A2(n_901),
.B(n_957),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_984),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1003),
.A2(n_832),
.B(n_856),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1009),
.A2(n_822),
.B(n_872),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1108),
.A2(n_906),
.B(n_907),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_982),
.B(n_857),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_981),
.B(n_862),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_983),
.A2(n_912),
.B(n_911),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1050),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_982),
.B(n_868),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1098),
.A2(n_900),
.B(n_843),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1006),
.A2(n_899),
.B(n_890),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1026),
.A2(n_1111),
.B(n_1118),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1022),
.A2(n_962),
.B(n_954),
.C(n_847),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1098),
.A2(n_846),
.B(n_852),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1073),
.B(n_895),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1018),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1025),
.A2(n_1051),
.B(n_1062),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1052),
.B(n_867),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1075),
.B(n_866),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1049),
.B(n_918),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1118),
.A2(n_848),
.B(n_884),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1028),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_995),
.B(n_918),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_987),
.A2(n_952),
.B(n_924),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1101),
.A2(n_930),
.B(n_955),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1110),
.A2(n_955),
.B1(n_951),
.B2(n_946),
.C(n_930),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1046),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1046),
.Y(n_1157)
);

OAI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1005),
.A2(n_879),
.B1(n_888),
.B2(n_898),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1007),
.A2(n_909),
.B(n_917),
.Y(n_1159)
);

AOI221x1_ASAP7_75t_L g1160 ( 
.A1(n_1054),
.A2(n_904),
.B1(n_921),
.B2(n_933),
.C(n_932),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1037),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1088),
.A2(n_964),
.B(n_942),
.C(n_931),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_986),
.B(n_892),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1008),
.A2(n_892),
.B(n_77),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1020),
.B(n_27),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1054),
.A2(n_1030),
.B(n_1016),
.C(n_1040),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_999),
.A2(n_892),
.B(n_74),
.C(n_72),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1072),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1020),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1061),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1015),
.A2(n_892),
.B(n_71),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1021),
.A2(n_66),
.B(n_30),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_SL g1173 ( 
.A(n_1041),
.B(n_29),
.Y(n_1173)
);

AO21x1_ASAP7_75t_L g1174 ( 
.A1(n_998),
.A2(n_30),
.B(n_33),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1089),
.A2(n_33),
.A3(n_35),
.B(n_37),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1030),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1042),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1019),
.A2(n_42),
.B(n_43),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_1023),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1106),
.A2(n_44),
.B(n_47),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1058),
.A2(n_50),
.B(n_55),
.C(n_57),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1058),
.A2(n_50),
.B(n_57),
.C(n_58),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_993),
.A2(n_58),
.B(n_62),
.C(n_1121),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1092),
.A2(n_1039),
.A3(n_1068),
.B(n_1038),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_989),
.A2(n_1095),
.B(n_1090),
.Y(n_1185)
);

AOI221xp5_ASAP7_75t_L g1186 ( 
.A1(n_1014),
.A2(n_1010),
.B1(n_1001),
.B2(n_1000),
.C(n_1044),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1107),
.A2(n_1102),
.A3(n_1091),
.B(n_1093),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1053),
.A2(n_1067),
.B(n_1031),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1100),
.A2(n_1013),
.B(n_1070),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1048),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_L g1191 ( 
.A1(n_1011),
.A2(n_1119),
.B(n_977),
.C(n_988),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_986),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1063),
.A2(n_1081),
.B(n_1087),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1056),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_1014),
.A2(n_1000),
.B1(n_991),
.B2(n_1031),
.C(n_1104),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1076),
.B(n_1085),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1055),
.A2(n_1035),
.B(n_1043),
.C(n_1103),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1027),
.A2(n_1034),
.B(n_1086),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1099),
.A2(n_1074),
.B(n_1077),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1064),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1080),
.A2(n_1036),
.B(n_1113),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_1061),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1117),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1099),
.A2(n_1116),
.B(n_1045),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_997),
.A2(n_992),
.B(n_1105),
.C(n_1094),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1080),
.A2(n_1004),
.B(n_1072),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1060),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1071),
.B(n_986),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1078),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1080),
.A2(n_1120),
.B(n_1115),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1078),
.A2(n_1094),
.B(n_1105),
.C(n_1083),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_985),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1080),
.A2(n_1067),
.B(n_1029),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1059),
.B(n_997),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1065),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1083),
.A2(n_1024),
.B1(n_1066),
.B2(n_1109),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1017),
.A2(n_1061),
.B(n_1082),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_975),
.B(n_1012),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1084),
.A2(n_1057),
.B(n_1114),
.C(n_1069),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1061),
.A2(n_1082),
.B(n_1096),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_985),
.A2(n_1117),
.B(n_1097),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1082),
.A2(n_1096),
.B(n_1079),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1082),
.A2(n_594),
.B(n_682),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1096),
.Y(n_1225)
);

NAND3x1_ASAP7_75t_L g1226 ( 
.A(n_1096),
.B(n_499),
.C(n_650),
.Y(n_1226)
);

AO32x2_ASAP7_75t_L g1227 ( 
.A1(n_998),
.A2(n_871),
.A3(n_886),
.B1(n_1039),
.B2(n_722),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_984),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_997),
.A2(n_663),
.B(n_647),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_976),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_976),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1117),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_979),
.A2(n_978),
.B(n_1015),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_984),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1050),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1049),
.B(n_986),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_980),
.B(n_794),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1089),
.A2(n_841),
.A3(n_916),
.B(n_871),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1022),
.A2(n_656),
.B1(n_650),
.B2(n_636),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_974),
.A2(n_812),
.B(n_672),
.C(n_978),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_994),
.B(n_494),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_984),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1090),
.A2(n_871),
.B(n_1095),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_984),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1022),
.A2(n_812),
.B(n_853),
.C(n_777),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1022),
.A2(n_948),
.B1(n_1054),
.B2(n_850),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1080),
.B(n_1072),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1022),
.A2(n_656),
.B1(n_650),
.B2(n_636),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_976),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_974),
.A2(n_812),
.B(n_672),
.C(n_978),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1049),
.B(n_986),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1112),
.B(n_810),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_984),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1047),
.A2(n_1108),
.B(n_903),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1089),
.A2(n_1092),
.B(n_1111),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1022),
.A2(n_656),
.B1(n_650),
.B2(n_636),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1117),
.Y(n_1264)
);

AOI221x1_ASAP7_75t_L g1265 ( 
.A1(n_1054),
.A2(n_1022),
.B1(n_1058),
.B2(n_1031),
.C(n_1110),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1041),
.Y(n_1267)
);

INVx3_ASAP7_75t_SL g1268 ( 
.A(n_1023),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1047),
.A2(n_1108),
.B(n_903),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_980),
.B(n_794),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_979),
.A2(n_594),
.B(n_682),
.Y(n_1271)
);

AO32x2_ASAP7_75t_L g1272 ( 
.A1(n_998),
.A2(n_871),
.A3(n_886),
.B1(n_1039),
.B2(n_722),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_980),
.B(n_794),
.Y(n_1273)
);

OAI21xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1249),
.A2(n_1171),
.B(n_1186),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1195),
.A2(n_1176),
.B1(n_1165),
.B2(n_1263),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1253),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1242),
.A2(n_1251),
.B1(n_1229),
.B2(n_1124),
.Y(n_1277)
);

BUFx10_ASAP7_75t_L g1278 ( 
.A(n_1137),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1240),
.A2(n_1273),
.B1(n_1270),
.B2(n_1210),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1196),
.A2(n_1229),
.B1(n_1226),
.B2(n_1256),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1228),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1236),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1250),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1245),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1231),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1247),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1267),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1174),
.A2(n_1273),
.B1(n_1270),
.B2(n_1240),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1122),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1122),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1259),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1244),
.B(n_1197),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1250),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1248),
.A2(n_1212),
.B1(n_1169),
.B2(n_1206),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1151),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1216),
.A2(n_1238),
.B1(n_1255),
.B2(n_1192),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1161),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1197),
.B(n_1152),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1171),
.A2(n_1222),
.B1(n_1234),
.B2(n_1213),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1179),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1217),
.A2(n_1123),
.B1(n_1147),
.B2(n_1198),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1234),
.A2(n_1199),
.B1(n_1215),
.B2(n_1135),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1168),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1238),
.A2(n_1255),
.B1(n_1209),
.B2(n_1173),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1204),
.Y(n_1306)
);

INVx6_ASAP7_75t_L g1307 ( 
.A(n_1149),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1177),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1265),
.A2(n_1215),
.B1(n_1222),
.B2(n_1157),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1268),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1199),
.A2(n_1125),
.B1(n_1193),
.B2(n_1188),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1190),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1156),
.A2(n_1188),
.B1(n_1149),
.B2(n_1262),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1134),
.A2(n_1138),
.B1(n_1230),
.B2(n_1148),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1237),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1194),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1225),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1201),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1223),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1262),
.A2(n_1139),
.B1(n_1208),
.B2(n_1136),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1145),
.A2(n_1128),
.B1(n_1144),
.B2(n_1127),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1143),
.A2(n_1200),
.B1(n_1214),
.B2(n_1129),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1219),
.B(n_1181),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1170),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1203),
.Y(n_1325)
);

INVx6_ASAP7_75t_L g1326 ( 
.A(n_1163),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1220),
.A2(n_1183),
.B1(n_1166),
.B2(n_1141),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1187),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1182),
.B(n_1243),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1163),
.A2(n_1178),
.B1(n_1211),
.B2(n_1180),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1233),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1126),
.A2(n_1172),
.B1(n_1164),
.B2(n_1264),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1233),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1191),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1264),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1175),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1129),
.A2(n_1126),
.B1(n_1158),
.B2(n_1202),
.Y(n_1337)
);

CKINVDCx8_ASAP7_75t_R g1338 ( 
.A(n_1221),
.Y(n_1338)
);

BUFx4_ASAP7_75t_R g1339 ( 
.A(n_1254),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1175),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1205),
.A2(n_1185),
.B1(n_1132),
.B2(n_1131),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1175),
.Y(n_1342)
);

BUFx2_ASAP7_75t_R g1343 ( 
.A(n_1167),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1207),
.A2(n_1159),
.B1(n_1272),
.B2(n_1227),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1160),
.A2(n_1218),
.B1(n_1246),
.B2(n_1271),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1187),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1187),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1153),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1140),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1241),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1154),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1241),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1189),
.A2(n_1150),
.B1(n_1133),
.B2(n_1266),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1142),
.A2(n_1235),
.B1(n_1261),
.B2(n_1258),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1232),
.A2(n_1257),
.B(n_1252),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1239),
.A2(n_1272),
.B1(n_1227),
.B2(n_1260),
.Y(n_1356)
);

INVx3_ASAP7_75t_SL g1357 ( 
.A(n_1155),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1184),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1224),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_R g1360 ( 
.A1(n_1227),
.A2(n_1272),
.B1(n_1155),
.B2(n_1184),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1184),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1162),
.B(n_1146),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1269),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1122),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1130),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1240),
.B(n_1270),
.Y(n_1367)
);

INVx5_ASAP7_75t_L g1368 ( 
.A(n_1168),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1253),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1242),
.A2(n_910),
.B1(n_1263),
.B2(n_1251),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1267),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1130),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1165),
.A2(n_910),
.B1(n_500),
.B2(n_330),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1240),
.B(n_1270),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1130),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1168),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1122),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1130),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1267),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1253),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1267),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1242),
.A2(n_650),
.B1(n_656),
.B2(n_910),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1122),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1168),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1130),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1390)
);

CKINVDCx11_ASAP7_75t_R g1391 ( 
.A(n_1267),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1122),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1267),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1231),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1122),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1240),
.B(n_1270),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1122),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1130),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1250),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1168),
.Y(n_1402)
);

BUFx8_ASAP7_75t_SL g1403 ( 
.A(n_1137),
.Y(n_1403)
);

BUFx2_ASAP7_75t_SL g1404 ( 
.A(n_1179),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1267),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1231),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1267),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1054),
.B2(n_1195),
.Y(n_1409)
);

BUFx2_ASAP7_75t_SL g1410 ( 
.A(n_1179),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1411)
);

AO21x1_ASAP7_75t_L g1412 ( 
.A1(n_1327),
.A2(n_1277),
.B(n_1370),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1394),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1357),
.B(n_1361),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1354),
.A2(n_1353),
.B(n_1341),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1367),
.B(n_1375),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1311),
.A2(n_1355),
.B(n_1274),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1396),
.B(n_1279),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1346),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1301),
.A2(n_1275),
.B(n_1294),
.C(n_1384),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_SL g1421 ( 
.A1(n_1329),
.A2(n_1321),
.B(n_1328),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1386),
.A2(n_1275),
.B(n_1365),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1373),
.A2(n_1374),
.B1(n_1376),
.B2(n_1400),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1347),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1319),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1336),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1339),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1285),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1340),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1351),
.Y(n_1430)
);

NAND4xp25_ASAP7_75t_L g1431 ( 
.A(n_1365),
.B(n_1384),
.C(n_1390),
.D(n_1398),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_R g1432 ( 
.A(n_1300),
.B(n_1371),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1352),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1292),
.B(n_1298),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1353),
.A2(n_1341),
.B(n_1322),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1350),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1350),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1374),
.A2(n_1398),
.B(n_1390),
.C(n_1400),
.Y(n_1438)
);

AOI221xp5_ASAP7_75t_L g1439 ( 
.A1(n_1376),
.A2(n_1409),
.B1(n_1408),
.B2(n_1380),
.C(n_1288),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1351),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1360),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_SL g1442 ( 
.A1(n_1321),
.A2(n_1409),
.B(n_1380),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1333),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1334),
.A2(n_1339),
.B1(n_1307),
.B2(n_1408),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1322),
.A2(n_1349),
.B(n_1362),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1302),
.B(n_1299),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1304),
.B(n_1314),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1276),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1280),
.A2(n_1334),
.B1(n_1309),
.B2(n_1307),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1281),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1282),
.Y(n_1451)
);

NAND2x1_ASAP7_75t_L g1452 ( 
.A(n_1319),
.B(n_1311),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1344),
.B(n_1284),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1286),
.B(n_1291),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1366),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1372),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1333),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1377),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1381),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1349),
.A2(n_1337),
.B(n_1320),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1389),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1348),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1399),
.B(n_1320),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1295),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1297),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1308),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1312),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1337),
.A2(n_1356),
.B(n_1288),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1325),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1316),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1318),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1406),
.B(n_1305),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1356),
.B(n_1363),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1323),
.A2(n_1359),
.B(n_1345),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1342),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1324),
.A2(n_1332),
.B(n_1331),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1342),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1306),
.A2(n_1283),
.B(n_1401),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1319),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1307),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1330),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_SL g1483 ( 
.A1(n_1335),
.A2(n_1315),
.B(n_1401),
.C(n_1293),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1338),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1313),
.B(n_1317),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_R g1486 ( 
.A(n_1382),
.B(n_1290),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1296),
.B(n_1383),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1293),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1326),
.B(n_1303),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1369),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1303),
.A2(n_1343),
.B(n_1368),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1368),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1368),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1368),
.A2(n_1364),
.B(n_1395),
.Y(n_1494)
);

BUFx12f_ASAP7_75t_L g1495 ( 
.A(n_1287),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1364),
.A2(n_1395),
.B1(n_1310),
.B2(n_1289),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1378),
.B(n_1388),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1378),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1402),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1364),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1395),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1404),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1310),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1475),
.B(n_1410),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1426),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1420),
.A2(n_1387),
.B(n_1397),
.C(n_1289),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1432),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1438),
.A2(n_1422),
.B(n_1439),
.C(n_1431),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1412),
.B(n_1397),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1423),
.A2(n_1300),
.B(n_1371),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1479),
.B(n_1379),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_SL g1512 ( 
.A1(n_1484),
.A2(n_1392),
.B(n_1387),
.C(n_1379),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1475),
.B(n_1392),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1469),
.B(n_1278),
.Y(n_1514)
);

AO22x2_ASAP7_75t_L g1515 ( 
.A1(n_1441),
.A2(n_1417),
.B1(n_1477),
.B2(n_1482),
.Y(n_1515)
);

AO32x1_ASAP7_75t_L g1516 ( 
.A1(n_1446),
.A2(n_1393),
.A3(n_1287),
.B1(n_1405),
.B2(n_1391),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1421),
.A2(n_1278),
.B(n_1391),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1413),
.B(n_1393),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1411),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1494),
.B(n_1385),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1477),
.B(n_1385),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1484),
.A2(n_1405),
.B(n_1407),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1485),
.B(n_1407),
.Y(n_1523)
);

NAND4xp25_ASAP7_75t_L g1524 ( 
.A(n_1447),
.B(n_1403),
.C(n_1418),
.D(n_1472),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1441),
.B(n_1403),
.Y(n_1525)
);

CKINVDCx6p67_ASAP7_75t_R g1526 ( 
.A(n_1495),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1485),
.B(n_1453),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1434),
.B(n_1416),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1415),
.A2(n_1435),
.B(n_1460),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1494),
.B(n_1430),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1446),
.A2(n_1468),
.B(n_1444),
.C(n_1415),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1532)
);

AND4x1_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1449),
.C(n_1501),
.D(n_1500),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1427),
.A2(n_1496),
.B1(n_1502),
.B2(n_1501),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1454),
.B(n_1474),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1428),
.B(n_1461),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1430),
.B(n_1440),
.Y(n_1537)
);

AO22x2_ASAP7_75t_L g1538 ( 
.A1(n_1482),
.A2(n_1442),
.B1(n_1421),
.B2(n_1426),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1468),
.A2(n_1435),
.B(n_1452),
.C(n_1491),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1474),
.B(n_1414),
.Y(n_1540)
);

AND2x6_ASAP7_75t_L g1541 ( 
.A(n_1463),
.B(n_1425),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1460),
.A2(n_1445),
.B(n_1429),
.Y(n_1542)
);

AOI211xp5_ASAP7_75t_L g1543 ( 
.A1(n_1487),
.A2(n_1483),
.B(n_1490),
.C(n_1500),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_SL g1544 ( 
.A1(n_1442),
.A2(n_1427),
.B(n_1464),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1427),
.A2(n_1487),
.B1(n_1448),
.B2(n_1474),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1463),
.A2(n_1414),
.B1(n_1470),
.B2(n_1459),
.C(n_1450),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1429),
.A2(n_1419),
.B(n_1424),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1450),
.B(n_1451),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1451),
.B(n_1455),
.Y(n_1549)
);

O2A1O1Ixp33_ASAP7_75t_SL g1550 ( 
.A1(n_1498),
.A2(n_1492),
.B(n_1493),
.C(n_1443),
.Y(n_1550)
);

AO21x2_ASAP7_75t_L g1551 ( 
.A1(n_1419),
.A2(n_1424),
.B(n_1437),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1456),
.B(n_1458),
.Y(n_1552)
);

AOI221xp5_ASAP7_75t_L g1553 ( 
.A1(n_1458),
.A2(n_1467),
.B1(n_1471),
.B2(n_1465),
.C(n_1470),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_SL g1554 ( 
.A(n_1476),
.B(n_1427),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1459),
.A2(n_1471),
.B1(n_1467),
.B2(n_1466),
.C(n_1465),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1491),
.A2(n_1478),
.B(n_1499),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1547),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1547),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1547),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1510),
.A2(n_1476),
.B1(n_1473),
.B2(n_1495),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1551),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1509),
.A2(n_1480),
.B1(n_1503),
.B2(n_1481),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1505),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1505),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1535),
.B(n_1433),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1551),
.Y(n_1566)
);

BUFx4f_ASAP7_75t_SL g1567 ( 
.A(n_1526),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1520),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1509),
.A2(n_1480),
.B1(n_1503),
.B2(n_1481),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1540),
.B(n_1542),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_1523),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1530),
.B(n_1462),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1529),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1462),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1437),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1548),
.B(n_1549),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1530),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1529),
.B(n_1436),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1524),
.A2(n_1480),
.B1(n_1481),
.B2(n_1476),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1537),
.B(n_1440),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1552),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1527),
.B(n_1532),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1515),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1519),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1515),
.A2(n_1481),
.B1(n_1489),
.B2(n_1488),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1557),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1570),
.B(n_1539),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1570),
.B(n_1539),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1558),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1559),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1573),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1570),
.B(n_1573),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1578),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1563),
.B(n_1515),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1573),
.B(n_1554),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1564),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1568),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1577),
.B(n_1537),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1561),
.A2(n_1531),
.B(n_1556),
.Y(n_1601)
);

OAI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1560),
.A2(n_1508),
.B(n_1506),
.C(n_1579),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1560),
.A2(n_1508),
.B1(n_1531),
.B2(n_1506),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1575),
.B(n_1537),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1583),
.A2(n_1538),
.B1(n_1526),
.B2(n_1520),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1522),
.C(n_1543),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1561),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1571),
.A2(n_1546),
.B1(n_1534),
.B2(n_1528),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1563),
.B(n_1553),
.Y(n_1611)
);

AND2x4_ASAP7_75t_SL g1612 ( 
.A(n_1580),
.B(n_1520),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1583),
.A2(n_1538),
.B1(n_1504),
.B2(n_1518),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1591),
.Y(n_1614)
);

OR2x2_ASAP7_75t_SL g1615 ( 
.A(n_1596),
.B(n_1514),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_R g1617 ( 
.A(n_1613),
.B(n_1486),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1591),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1612),
.B(n_1568),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1612),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1610),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1599),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1612),
.B(n_1568),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1591),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1611),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1598),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1598),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1588),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1588),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1586),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1604),
.A2(n_1533),
.B(n_1585),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1586),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1589),
.B(n_1572),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1603),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1588),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1589),
.B(n_1574),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1595),
.B(n_1584),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1590),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1589),
.B(n_1584),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1590),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1604),
.A2(n_1517),
.B1(n_1541),
.B2(n_1544),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1595),
.B(n_1582),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1589),
.B(n_1574),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1612),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1636),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1627),
.B(n_1594),
.Y(n_1653)
);

AO32x1_ASAP7_75t_L g1654 ( 
.A1(n_1623),
.A2(n_1604),
.A3(n_1610),
.B1(n_1599),
.B2(n_1586),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1614),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1612),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1616),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1636),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1593),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1605),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1627),
.B(n_1594),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1623),
.B(n_1593),
.Y(n_1662)
);

AOI31xp33_ASAP7_75t_L g1663 ( 
.A1(n_1622),
.A2(n_1602),
.A3(n_1610),
.B(n_1512),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1614),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1618),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1567),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1618),
.Y(n_1667)
);

NOR2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1646),
.B(n_1525),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1628),
.Y(n_1669)
);

NAND4xp75_ASAP7_75t_L g1670 ( 
.A(n_1637),
.B(n_1593),
.C(n_1516),
.D(n_1521),
.Y(n_1670)
);

AOI222xp33_ASAP7_75t_L g1671 ( 
.A1(n_1648),
.A2(n_1602),
.B1(n_1613),
.B2(n_1507),
.C1(n_1606),
.C2(n_1616),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1636),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1619),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1626),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1626),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1638),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1621),
.B(n_1605),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1638),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1638),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1628),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1634),
.B(n_1600),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1646),
.A2(n_1607),
.B(n_1602),
.C(n_1512),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1641),
.Y(n_1689)
);

NAND2x1_ASAP7_75t_L g1690 ( 
.A(n_1619),
.B(n_1599),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1644),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1634),
.B(n_1600),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1644),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1629),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1656),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1674),
.B(n_1639),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1655),
.Y(n_1697)
);

XNOR2xp5_ASAP7_75t_L g1698 ( 
.A(n_1668),
.B(n_1607),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1657),
.B(n_1629),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1655),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1674),
.B(n_1639),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1653),
.B(n_1615),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1640),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1694),
.B(n_1630),
.Y(n_1705)
);

OAI211xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1671),
.A2(n_1607),
.B(n_1606),
.C(n_1647),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1694),
.B(n_1630),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1653),
.B(n_1615),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1685),
.B(n_1632),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1661),
.B(n_1632),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1664),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1661),
.B(n_1649),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1659),
.B(n_1645),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1659),
.B(n_1645),
.Y(n_1715)
);

AO21x1_ASAP7_75t_L g1716 ( 
.A1(n_1663),
.A2(n_1647),
.B(n_1590),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1664),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_SL g1719 ( 
.A1(n_1662),
.A2(n_1651),
.B1(n_1620),
.B2(n_1649),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_SL g1720 ( 
.A(n_1687),
.B(n_1599),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1673),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1687),
.B(n_1617),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1673),
.B(n_1582),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1601),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1665),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1682),
.B(n_1601),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1685),
.B(n_1631),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1667),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1656),
.B(n_1677),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1656),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1697),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1698),
.B(n_1671),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1722),
.A2(n_1666),
.B1(n_1601),
.B2(n_1662),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1701),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1722),
.A2(n_1670),
.B1(n_1601),
.B2(n_1656),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1663),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1695),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1699),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1703),
.A2(n_1670),
.B1(n_1651),
.B2(n_1620),
.Y(n_1740)
);

XOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1708),
.B(n_1513),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1713),
.B(n_1690),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1706),
.A2(n_1654),
.B(n_1689),
.C(n_1516),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1715),
.A2(n_1730),
.B1(n_1729),
.B2(n_1651),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_L g1745 ( 
.A(n_1720),
.B(n_1689),
.C(n_1691),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1714),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1711),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1706),
.A2(n_1654),
.B(n_1516),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1705),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1716),
.B(n_1691),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1705),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1707),
.A2(n_1690),
.B1(n_1625),
.B2(n_1619),
.Y(n_1754)
);

OAI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1719),
.A2(n_1693),
.B1(n_1654),
.B2(n_1688),
.C(n_1667),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1700),
.A2(n_1601),
.B1(n_1707),
.B2(n_1709),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1736),
.A2(n_1710),
.B1(n_1712),
.B2(n_1654),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1739),
.B(n_1732),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1738),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1739),
.Y(n_1760)
);

AOI31xp33_ASAP7_75t_L g1761 ( 
.A1(n_1737),
.A2(n_1702),
.A3(n_1704),
.B(n_1700),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1742),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1749),
.A2(n_1740),
.B1(n_1733),
.B2(n_1745),
.Y(n_1763)
);

OAI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1743),
.A2(n_1709),
.B1(n_1727),
.B2(n_1693),
.C(n_1725),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1735),
.B(n_1750),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1747),
.B(n_1693),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1753),
.B(n_1717),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1744),
.A2(n_1746),
.B1(n_1754),
.B2(n_1751),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1731),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1746),
.B(n_1723),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1751),
.A2(n_1601),
.B1(n_1677),
.B2(n_1728),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1734),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1741),
.B(n_1718),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1727),
.Y(n_1774)
);

OAI21xp33_ASAP7_75t_SL g1775 ( 
.A1(n_1756),
.A2(n_1679),
.B(n_1660),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1733),
.A2(n_1654),
.B1(n_1724),
.B2(n_1726),
.C(n_1688),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1763),
.A2(n_1758),
.B1(n_1768),
.B2(n_1764),
.C(n_1775),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1760),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1759),
.B(n_1752),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1765),
.Y(n_1780)
);

AO22x1_ASAP7_75t_L g1781 ( 
.A1(n_1758),
.A2(n_1688),
.B1(n_1654),
.B2(n_1677),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1761),
.B(n_1756),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1771),
.A2(n_1742),
.B1(n_1755),
.B2(n_1677),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1762),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1770),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1757),
.B(n_1536),
.C(n_1652),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1773),
.B(n_1619),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1766),
.B(n_1679),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1780),
.Y(n_1789)
);

NAND4xp75_ASAP7_75t_L g1790 ( 
.A(n_1782),
.B(n_1767),
.C(n_1772),
.D(n_1769),
.Y(n_1790)
);

OAI21xp33_ASAP7_75t_L g1791 ( 
.A1(n_1777),
.A2(n_1774),
.B(n_1767),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_SL g1792 ( 
.A(n_1779),
.B(n_1776),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1783),
.A2(n_1675),
.B1(n_1676),
.B2(n_1684),
.C(n_1652),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1785),
.B(n_1681),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1784),
.Y(n_1795)
);

NOR3x1_ASAP7_75t_L g1796 ( 
.A(n_1787),
.B(n_1675),
.C(n_1676),
.Y(n_1796)
);

NAND4xp25_ASAP7_75t_SL g1797 ( 
.A(n_1786),
.B(n_1516),
.C(n_1686),
.D(n_1692),
.Y(n_1797)
);

NAND4xp25_ASAP7_75t_L g1798 ( 
.A(n_1778),
.B(n_1569),
.C(n_1562),
.D(n_1683),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1791),
.A2(n_1783),
.B1(n_1781),
.B2(n_1788),
.C(n_1684),
.Y(n_1799)
);

OA211x2_ASAP7_75t_L g1800 ( 
.A1(n_1792),
.A2(n_1555),
.B(n_1576),
.C(n_1625),
.Y(n_1800)
);

AOI322xp5_ASAP7_75t_L g1801 ( 
.A1(n_1789),
.A2(n_1592),
.A3(n_1595),
.B1(n_1603),
.B2(n_1597),
.C1(n_1692),
.C2(n_1686),
.Y(n_1801)
);

O2A1O1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1795),
.A2(n_1684),
.B(n_1652),
.C(n_1658),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1793),
.A2(n_1625),
.B(n_1597),
.C(n_1592),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1799),
.A2(n_1794),
.B1(n_1798),
.B2(n_1790),
.C(n_1797),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1800),
.A2(n_1631),
.B1(n_1633),
.B2(n_1642),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1803),
.A2(n_1796),
.B(n_1658),
.C(n_1672),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1801),
.A2(n_1802),
.B(n_1672),
.C(n_1658),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1799),
.A2(n_1680),
.B1(n_1678),
.B2(n_1672),
.C(n_1597),
.Y(n_1808)
);

OAI21xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1799),
.A2(n_1681),
.B(n_1683),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1805),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1804),
.A2(n_1680),
.B1(n_1678),
.B2(n_1517),
.Y(n_1811)
);

XNOR2xp5_ASAP7_75t_L g1812 ( 
.A(n_1808),
.B(n_1511),
.Y(n_1812)
);

NOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1678),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1806),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1810),
.B(n_1809),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1814),
.A2(n_1680),
.B(n_1603),
.C(n_1592),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1811),
.B(n_1640),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1815),
.Y(n_1818)
);

NAND4xp25_ASAP7_75t_L g1819 ( 
.A(n_1818),
.B(n_1817),
.C(n_1816),
.D(n_1813),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1812),
.B(n_1625),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1819),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1821),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1820),
.A2(n_1642),
.B1(n_1633),
.B2(n_1595),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1822),
.B(n_1823),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1822),
.A2(n_1650),
.B(n_1643),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1824),
.A2(n_1650),
.B(n_1643),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1825),
.B(n_1511),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1827),
.Y(n_1828)
);

OAI221xp5_ASAP7_75t_R g1829 ( 
.A1(n_1828),
.A2(n_1608),
.B1(n_1609),
.B2(n_1599),
.C(n_1550),
.Y(n_1829)
);

AOI211xp5_ASAP7_75t_L g1830 ( 
.A1(n_1829),
.A2(n_1497),
.B(n_1457),
.C(n_1443),
.Y(n_1830)
);


endmodule