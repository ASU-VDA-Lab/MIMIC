module fake_ariane_1061_n_187 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_187);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_187;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_118;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_3),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_3),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_4),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_4),
.Y(n_65)
);

AND3x1_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_6),
.C(n_7),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_8),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_42),
.B1(n_47),
.B2(n_46),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_52),
.B1(n_51),
.B2(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

OAI221xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_43),
.B1(n_47),
.B2(n_42),
.C(n_9),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_66),
.B1(n_57),
.B2(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_75),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_78),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_79),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_79),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_79),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_100),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_97),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_99),
.B(n_83),
.C(n_96),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_97),
.B(n_91),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_115),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_81),
.B(n_105),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_111),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_118),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_120),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_127),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_116),
.C(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_104),
.B1(n_110),
.B2(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_124),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_125),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_129),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_129),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_130),
.C(n_56),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_123),
.Y(n_156)
);

NAND2x1_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_128),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_58),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_156),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_157),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_132),
.B(n_128),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_117),
.B(n_133),
.Y(n_167)
);

NAND4xp25_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_56),
.C(n_89),
.D(n_64),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_64),
.Y(n_169)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_153),
.B(n_77),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_133),
.B(n_117),
.C(n_55),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_96),
.C(n_88),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_55),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_77),
.B1(n_95),
.B2(n_55),
.Y(n_176)
);

AND4x1_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_55),
.C(n_77),
.D(n_13),
.Y(n_177)
);

NOR3x1_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_164),
.C(n_77),
.Y(n_178)
);

AOI222xp33_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_95),
.B1(n_93),
.B2(n_14),
.C1(n_18),
.C2(n_20),
.Y(n_179)
);

NAND2x1p5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_93),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_173),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_176),
.B1(n_172),
.B2(n_177),
.Y(n_183)
);

AOI211xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_170),
.B(n_12),
.C(n_23),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_180),
.B(n_93),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_184),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_183),
.B1(n_25),
.B2(n_30),
.Y(n_187)
);


endmodule