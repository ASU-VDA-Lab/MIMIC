module fake_jpeg_25050_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_63),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_52),
.B1(n_61),
.B2(n_50),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_88),
.B1(n_58),
.B2(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.Y(n_92)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_57),
.B1(n_50),
.B2(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_102),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_85),
.B1(n_79),
.B2(n_83),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_70),
.B(n_49),
.C(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_60),
.B1(n_59),
.B2(n_55),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_54),
.B1(n_46),
.B2(n_56),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_59),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_115),
.B1(n_118),
.B2(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_47),
.B1(n_19),
.B2(n_20),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_17),
.B1(n_43),
.B2(n_40),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_122),
.B1(n_108),
.B2(n_4),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_95),
.B1(n_103),
.B2(n_107),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_96),
.C(n_107),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_96),
.B(n_2),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_117),
.B(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_15),
.C(n_39),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_45),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_134),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_126),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_117),
.B(n_115),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_2),
.B(n_5),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_141),
.B1(n_10),
.B2(n_12),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_9),
.Y(n_144)
);

AO32x1_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_29),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_14),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_34),
.B1(n_18),
.B2(n_21),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_146),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_159),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_143),
.C(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_155),
.C(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_153),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_148),
.B(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_154),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_154),
.C(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_149),
.C(n_150),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_36),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_144),
.C(n_23),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_37),
.B(n_32),
.Y(n_170)
);


endmodule