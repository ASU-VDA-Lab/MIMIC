module fake_netlist_5_1436_n_1254 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1254);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1254;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_731;
wire n_371;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_582;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_577;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_384;
wire n_1061;
wire n_462;
wire n_1193;
wire n_1113;
wire n_1226;
wire n_722;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_1251;

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_208),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_80),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_188),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_42),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_336),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_147),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_17),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_190),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_300),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_213),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_53),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_273),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_225),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_85),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_127),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_121),
.B(n_142),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_278),
.Y(n_361)
);

BUFx8_ASAP7_75t_SL g362 ( 
.A(n_269),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_151),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_83),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_141),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_272),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_133),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_251),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_81),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_181),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_217),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_43),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_34),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_104),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_329),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_201),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_293),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_335),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_135),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_224),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_18),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_232),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_282),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_36),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_252),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_191),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_86),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_87),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_315),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_136),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_19),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_7),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_182),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_292),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_294),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_199),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_157),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_57),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_77),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_140),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_289),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_44),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_154),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_178),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_149),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_155),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_46),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_100),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_3),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_82),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_114),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_254),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_138),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_197),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_110),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_70),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_94),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_226),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_277),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_331),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_200),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_123),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_132),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_337),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_174),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_20),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_73),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_284),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_274),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_50),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_63),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_161),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_156),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_95),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_192),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_306),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_341),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_44),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_108),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_316),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_51),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_139),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_270),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_184),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_266),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_320),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_183),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_158),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_159),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_290),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_253),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_103),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_80),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_120),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_249),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_143),
.B(n_338),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_55),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_56),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_3),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_45),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_204),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_260),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_99),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_210),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_126),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_187),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_311),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_58),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_84),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_291),
.Y(n_471)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_106),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_302),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_206),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_288),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_137),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_102),
.Y(n_477)
);

BUFx5_ASAP7_75t_L g478 ( 
.A(n_227),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_205),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_340),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_152),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_257),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_134),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_49),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_308),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_146),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_408),
.B(n_0),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

BUFx8_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_394),
.B(n_0),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_348),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_344),
.A2(n_356),
.B(n_354),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_348),
.Y(n_493)
);

CKINVDCx6p67_ASAP7_75t_R g494 ( 
.A(n_373),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_348),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_348),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_410),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_351),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_386),
.B(n_401),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

OA21x2_ASAP7_75t_L g504 ( 
.A1(n_357),
.A2(n_1),
.B(n_2),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_397),
.B(n_1),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_352),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_351),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_343),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_2),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_469),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_369),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_472),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_472),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_4),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_400),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_517)
);

INVxp33_ASAP7_75t_SL g518 ( 
.A(n_372),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_377),
.B(n_5),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_403),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_391),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_382),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_427),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_355),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_472),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_359),
.B(n_8),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_377),
.B(n_9),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_443),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_431),
.B(n_9),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_464),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_391),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_346),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_485),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_409),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_450),
.B(n_10),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_362),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_454),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_478),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_450),
.B(n_406),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_434),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_434),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_364),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_385),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_478),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_365),
.B(n_11),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_366),
.B(n_11),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_461),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_367),
.A2(n_374),
.B(n_371),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_484),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_380),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_345),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_406),
.B(n_12),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_392),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_389),
.B(n_13),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_540),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_518),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_523),
.B(n_342),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_522),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_523),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_537),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_493),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_500),
.B(n_350),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_496),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_535),
.Y(n_570)
);

BUFx4f_ASAP7_75t_L g571 ( 
.A(n_492),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_498),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_559),
.B(n_363),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_535),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_500),
.B(n_395),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_507),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_R g577 ( 
.A(n_559),
.B(n_358),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_547),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_489),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_489),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_495),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_494),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_500),
.B(n_398),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_497),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_538),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_491),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_544),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_491),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_500),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_508),
.B(n_456),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_508),
.B(n_479),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_488),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_508),
.Y(n_596)
);

AOI22x1_ASAP7_75t_SL g597 ( 
.A1(n_517),
.A2(n_399),
.B1(n_417),
.B2(n_393),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_534),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_534),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_534),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_R g601 ( 
.A(n_551),
.B(n_361),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_534),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_R g603 ( 
.A(n_551),
.B(n_368),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_543),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_525),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_556),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_503),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_503),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_506),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_506),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_515),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_607),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_608),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_601),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_569),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_606),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_567),
.B(n_492),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_604),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_604),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_569),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_573),
.B(n_543),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_570),
.B(n_490),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_574),
.B(n_531),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_568),
.B(n_505),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_501),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_590),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_601),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_592),
.B(n_558),
.C(n_539),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_554),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_593),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_582),
.B(n_531),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_594),
.B(n_510),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_585),
.B(n_554),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_610),
.B(n_516),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_589),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_571),
.B(n_513),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_577),
.B(n_487),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_572),
.B(n_514),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_575),
.B(n_521),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_584),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_603),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_612),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_599),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_605),
.B(n_526),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_529),
.Y(n_652)
);

BUFx6f_ASAP7_75t_SL g653 ( 
.A(n_563),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_588),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_530),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_501),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_600),
.B(n_502),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_602),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_502),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_583),
.B(n_558),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_561),
.B(n_511),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_579),
.B(n_539),
.C(n_528),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_564),
.B(n_542),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_566),
.B(n_548),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_597),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_563),
.B(n_515),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_581),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_595),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_569),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g672 ( 
.A(n_586),
.B(n_528),
.C(n_519),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_573),
.B(n_515),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_563),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_567),
.B(n_525),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_580),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_586),
.B(n_519),
.C(n_560),
.Y(n_677)
);

OR2x2_ASAP7_75t_SL g678 ( 
.A(n_586),
.B(n_524),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_567),
.B(n_525),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_573),
.B(n_511),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_614),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_653),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_648),
.B(n_383),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_645),
.B(n_549),
.Y(n_684)
);

AND2x6_ASAP7_75t_SL g685 ( 
.A(n_660),
.B(n_532),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_651),
.B(n_421),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_656),
.B(n_549),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_673),
.B(n_550),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_669),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_676),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_680),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_631),
.B(n_635),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_630),
.A2(n_424),
.B1(n_440),
.B2(n_430),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_675),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_631),
.B(n_550),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_648),
.B(n_445),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_675),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_640),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_662),
.B(n_616),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_626),
.B(n_641),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_629),
.B(n_524),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_627),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_641),
.A2(n_457),
.B(n_360),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_650),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_620),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_625),
.B(n_463),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_659),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_644),
.B(n_533),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_679),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_679),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_621),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_628),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_639),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_632),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_653),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_647),
.B(n_467),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_652),
.B(n_533),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_636),
.A2(n_619),
.B1(n_504),
.B2(n_672),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_615),
.B(n_541),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_678),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_642),
.B(n_447),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_637),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_654),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_618),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_632),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_652),
.B(n_536),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_677),
.A2(n_349),
.B1(n_353),
.B2(n_347),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_655),
.B(n_536),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_613),
.B(n_509),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_667),
.B(n_504),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_643),
.Y(n_732)
);

CKINVDCx8_ASAP7_75t_R g733 ( 
.A(n_658),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_633),
.B(n_432),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_666),
.B(n_527),
.Y(n_735)
);

NOR2x1_ASAP7_75t_R g736 ( 
.A(n_668),
.B(n_442),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_638),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_674),
.B(n_541),
.Y(n_738)
);

INVx5_ASAP7_75t_L g739 ( 
.A(n_659),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_670),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_664),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_649),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_664),
.B(n_458),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_665),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_622),
.B(n_411),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_SL g747 ( 
.A1(n_661),
.A2(n_517),
.B1(n_520),
.B2(n_557),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_657),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_671),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_663),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_646),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_624),
.B(n_459),
.Y(n_753)
);

NOR2x2_ASAP7_75t_L g754 ( 
.A(n_666),
.B(n_520),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_614),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_680),
.B(n_512),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_623),
.B(n_370),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_676),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_614),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_623),
.B(n_375),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_707),
.B(n_739),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_722),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_692),
.B(n_441),
.Y(n_763)
);

AOI221x1_ASAP7_75t_L g764 ( 
.A1(n_703),
.A2(n_449),
.B1(n_455),
.B2(n_446),
.C(n_444),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_752),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_695),
.A2(n_465),
.B(n_462),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_684),
.A2(n_475),
.B(n_378),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_721),
.A2(n_557),
.B(n_379),
.C(n_381),
.Y(n_768)
);

INVx3_ASAP7_75t_SL g769 ( 
.A(n_682),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_707),
.B(n_376),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_741),
.B(n_384),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_681),
.Y(n_772)
);

BUFx12f_ASAP7_75t_L g773 ( 
.A(n_715),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_745),
.B(n_387),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_732),
.B(n_388),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_727),
.B(n_390),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_690),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_707),
.B(n_552),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_740),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_752),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_718),
.A2(n_402),
.B1(n_404),
.B2(n_396),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_688),
.A2(n_407),
.B1(n_412),
.B2(n_405),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_755),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_686),
.B(n_413),
.Y(n_784)
);

NAND2x2_ASAP7_75t_L g785 ( 
.A(n_742),
.B(n_414),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_758),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_717),
.A2(n_416),
.B(n_415),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_689),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_753),
.A2(n_419),
.B(n_420),
.C(n_418),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_726),
.A2(n_425),
.B(n_423),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_694),
.B(n_426),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_697),
.B(n_709),
.Y(n_792)
);

OA22x2_ASAP7_75t_L g793 ( 
.A1(n_750),
.A2(n_555),
.B1(n_553),
.B2(n_436),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_759),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_708),
.A2(n_478),
.B(n_438),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_710),
.B(n_433),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_758),
.Y(n_797)
);

CKINVDCx10_ASAP7_75t_R g798 ( 
.A(n_754),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_729),
.A2(n_452),
.B(n_451),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_712),
.Y(n_800)
);

AO32x1_ASAP7_75t_L g801 ( 
.A1(n_744),
.A2(n_478),
.A3(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_702),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_713),
.B(n_466),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_752),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_743),
.A2(n_470),
.B1(n_471),
.B2(n_468),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_706),
.A2(n_474),
.B1(n_476),
.B2(n_473),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_711),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_687),
.A2(n_480),
.B1(n_481),
.B2(n_477),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_748),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_725),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_691),
.A2(n_483),
.B(n_482),
.C(n_546),
.Y(n_811)
);

AO21x1_ASAP7_75t_L g812 ( 
.A1(n_731),
.A2(n_16),
.B(n_17),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_757),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_738),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_724),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_SL g816 ( 
.A(n_739),
.B(n_22),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_760),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_720),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_714),
.Y(n_819)
);

OAI21xp33_ASAP7_75t_SL g820 ( 
.A1(n_756),
.A2(n_26),
.B(n_27),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_704),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_701),
.B(n_27),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_751),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_749),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_730),
.B(n_88),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_705),
.B(n_28),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_SL g827 ( 
.A1(n_747),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_737),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_746),
.A2(n_90),
.B(n_89),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_699),
.A2(n_92),
.B(n_91),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_698),
.B(n_93),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_730),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_723),
.B(n_96),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_705),
.B(n_29),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_683),
.A2(n_98),
.B(n_97),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_696),
.A2(n_105),
.B(n_101),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_716),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_837)
);

XNOR2xp5_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_107),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_733),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_735),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_734),
.B(n_32),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_685),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_735),
.Y(n_843)
);

OAI21xp33_ASAP7_75t_L g844 ( 
.A1(n_736),
.A2(n_36),
.B(n_37),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_681),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_SL g846 ( 
.A1(n_700),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_721),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_719),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_722),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_SL g850 ( 
.A1(n_743),
.A2(n_111),
.B(n_112),
.C(n_109),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_719),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_722),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_722),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_700),
.A2(n_115),
.B1(n_116),
.B2(n_113),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_SL g855 ( 
.A1(n_743),
.A2(n_118),
.B(n_119),
.C(n_117),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_722),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_681),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_721),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_700),
.B(n_46),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_722),
.B(n_47),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_700),
.B(n_48),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_719),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_719),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_722),
.B(n_49),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_741),
.B(n_50),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_681),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_721),
.A2(n_124),
.B1(n_125),
.B2(n_122),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_700),
.B(n_52),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_741),
.B(n_54),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_741),
.B(n_54),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_700),
.B(n_55),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_700),
.B(n_56),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_721),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_873)
);

BUFx2_ASAP7_75t_SL g874 ( 
.A(n_722),
.Y(n_874)
);

OAI22x1_ASAP7_75t_L g875 ( 
.A1(n_693),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_875)
);

BUFx10_ASAP7_75t_L g876 ( 
.A(n_841),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

OAI21x1_ASAP7_75t_SL g878 ( 
.A1(n_812),
.A2(n_129),
.B(n_128),
.Y(n_878)
);

AO21x2_ASAP7_75t_L g879 ( 
.A1(n_826),
.A2(n_131),
.B(n_130),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_788),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_762),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_762),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_802),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_765),
.Y(n_884)
);

BUFx2_ASAP7_75t_R g885 ( 
.A(n_874),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_765),
.Y(n_886)
);

CKINVDCx8_ASAP7_75t_R g887 ( 
.A(n_762),
.Y(n_887)
);

AO21x2_ASAP7_75t_L g888 ( 
.A1(n_834),
.A2(n_763),
.B(n_795),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_851),
.B(n_62),
.Y(n_889)
);

CKINVDCx10_ASAP7_75t_R g890 ( 
.A(n_798),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_780),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_862),
.B(n_64),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_852),
.Y(n_893)
);

CKINVDCx6p67_ASAP7_75t_R g894 ( 
.A(n_769),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_772),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_792),
.B(n_64),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_859),
.A2(n_145),
.B(n_144),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_852),
.Y(n_898)
);

AOI22x1_ASAP7_75t_L g899 ( 
.A1(n_875),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_804),
.B(n_832),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_783),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_784),
.B(n_65),
.Y(n_902)
);

AOI22x1_ASAP7_75t_L g903 ( 
.A1(n_766),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_903)
);

AOI22x1_ASAP7_75t_L g904 ( 
.A1(n_835),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_904)
);

OAI21x1_ASAP7_75t_SL g905 ( 
.A1(n_836),
.A2(n_150),
.B(n_148),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_780),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_853),
.B(n_153),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_814),
.B(n_71),
.Y(n_908)
);

OAI21x1_ASAP7_75t_SL g909 ( 
.A1(n_813),
.A2(n_162),
.B(n_160),
.Y(n_909)
);

BUFx2_ASAP7_75t_SL g910 ( 
.A(n_853),
.Y(n_910)
);

NOR2x1_ASAP7_75t_L g911 ( 
.A(n_828),
.B(n_163),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_794),
.Y(n_912)
);

AO21x2_ASAP7_75t_L g913 ( 
.A1(n_861),
.A2(n_165),
.B(n_164),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_868),
.A2(n_167),
.B(n_166),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_866),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_824),
.A2(n_169),
.B(n_168),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_800),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_839),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_797),
.B(n_170),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_845),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_780),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_779),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_871),
.A2(n_172),
.B(n_171),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_786),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_764),
.A2(n_175),
.B(n_173),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_810),
.A2(n_177),
.B(n_176),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_856),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_807),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_848),
.B(n_72),
.Y(n_929)
);

CKINVDCx11_ASAP7_75t_R g930 ( 
.A(n_773),
.Y(n_930)
);

CKINVDCx6p67_ASAP7_75t_R g931 ( 
.A(n_821),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_872),
.A2(n_180),
.B(n_179),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_777),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_857),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_863),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_809),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_823),
.B(n_73),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_818),
.Y(n_938)
);

AO21x2_ASAP7_75t_L g939 ( 
.A1(n_850),
.A2(n_186),
.B(n_185),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_793),
.Y(n_940)
);

INVx8_ASAP7_75t_L g941 ( 
.A(n_825),
.Y(n_941)
);

CKINVDCx6p67_ASAP7_75t_R g942 ( 
.A(n_843),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_815),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_771),
.B(n_74),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_819),
.Y(n_945)
);

BUFx2_ASAP7_75t_R g946 ( 
.A(n_785),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_825),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_860),
.Y(n_949)
);

OR3x4_ASAP7_75t_SL g950 ( 
.A(n_827),
.B(n_75),
.C(n_76),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_840),
.B(n_193),
.Y(n_951)
);

OR3x4_ASAP7_75t_SL g952 ( 
.A(n_842),
.B(n_75),
.C(n_76),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_855),
.A2(n_195),
.B(n_194),
.Y(n_953)
);

AOI22x1_ASAP7_75t_L g954 ( 
.A1(n_822),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_791),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_789),
.A2(n_767),
.B(n_796),
.Y(n_956)
);

INVx6_ASAP7_75t_L g957 ( 
.A(n_864),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_803),
.B(n_78),
.C(n_79),
.Y(n_958)
);

AOI22x1_ASAP7_75t_L g959 ( 
.A1(n_838),
.A2(n_81),
.B1(n_196),
.B2(n_198),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_865),
.B(n_339),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_774),
.B(n_776),
.Y(n_961)
);

BUFx2_ASAP7_75t_SL g962 ( 
.A(n_761),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_816),
.B(n_833),
.Y(n_963)
);

BUFx12f_ASAP7_75t_L g964 ( 
.A(n_778),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_775),
.A2(n_790),
.B(n_787),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_831),
.A2(n_202),
.B(n_203),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_869),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_829),
.A2(n_207),
.B(n_209),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_870),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_820),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_770),
.B(n_211),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_846),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_830),
.A2(n_212),
.B(n_214),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_817),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_854),
.A2(n_215),
.B(n_216),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_837),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_805),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_867),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_801),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_806),
.Y(n_980)
);

BUFx8_ASAP7_75t_L g981 ( 
.A(n_844),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_808),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_847),
.Y(n_983)
);

AO21x2_ASAP7_75t_L g984 ( 
.A1(n_799),
.A2(n_221),
.B(n_222),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_858),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_781),
.Y(n_986)
);

AO21x2_ASAP7_75t_L g987 ( 
.A1(n_811),
.A2(n_223),
.B(n_228),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_895),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_895),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_917),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_883),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_928),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_917),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_920),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_893),
.Y(n_995)
);

CKINVDCx11_ASAP7_75t_R g996 ( 
.A(n_930),
.Y(n_996)
);

OAI22xp33_ASAP7_75t_L g997 ( 
.A1(n_902),
.A2(n_782),
.B1(n_768),
.B2(n_873),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_980),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_998)
);

INVx6_ASAP7_75t_L g999 ( 
.A(n_933),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_955),
.B(n_233),
.Y(n_1000)
);

OAI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_948),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_918),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_978),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_934),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_981),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_982),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_894),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_880),
.Y(n_1008)
);

BUFx2_ASAP7_75t_R g1009 ( 
.A(n_877),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_983),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_1010)
);

BUFx8_ASAP7_75t_L g1011 ( 
.A(n_936),
.Y(n_1011)
);

BUFx10_ASAP7_75t_L g1012 ( 
.A(n_889),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_938),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_922),
.B(n_250),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_924),
.Y(n_1015)
);

AO21x1_ASAP7_75t_L g1016 ( 
.A1(n_944),
.A2(n_255),
.B(n_256),
.Y(n_1016)
);

CKINVDCx11_ASAP7_75t_R g1017 ( 
.A(n_887),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_983),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_961),
.B(n_262),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_969),
.B(n_263),
.Y(n_1020)
);

AO21x1_ASAP7_75t_L g1021 ( 
.A1(n_960),
.A2(n_264),
.B(n_265),
.Y(n_1021)
);

CKINVDCx11_ASAP7_75t_R g1022 ( 
.A(n_931),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_912),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_885),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_943),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_901),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_881),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_882),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_935),
.B(n_267),
.Y(n_1029)
);

INVx6_ASAP7_75t_L g1030 ( 
.A(n_948),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_896),
.B(n_268),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_915),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_892),
.B(n_271),
.Y(n_1033)
);

AOI222xp33_ASAP7_75t_L g1034 ( 
.A1(n_981),
.A2(n_275),
.B1(n_276),
.B2(n_279),
.C1(n_280),
.C2(n_281),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_937),
.B(n_283),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_957),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_947),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_945),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_951),
.Y(n_1039)
);

BUFx2_ASAP7_75t_SL g1040 ( 
.A(n_948),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_976),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_908),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_986),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_957),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_898),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_974),
.B(n_295),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_900),
.B(n_296),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_986),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_985),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_900),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_940),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_971),
.A2(n_305),
.B1(n_307),
.B2(n_309),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_876),
.B(n_310),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_884),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_SL g1055 ( 
.A1(n_959),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_949),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_886),
.Y(n_1057)
);

INVx6_ASAP7_75t_L g1058 ( 
.A(n_927),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_970),
.A2(n_318),
.B(n_319),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_942),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_SL g1061 ( 
.A1(n_899),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_891),
.B(n_324),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_899),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_1063)
);

INVxp67_ASAP7_75t_SL g1064 ( 
.A(n_891),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_906),
.Y(n_1065)
);

OAI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_941),
.A2(n_328),
.B1(n_330),
.B2(n_332),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_916),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_996),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_1007),
.B(n_958),
.C(n_952),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_991),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_1040),
.B(n_910),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_1002),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_1044),
.B(n_910),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_R g1074 ( 
.A(n_1015),
.B(n_1056),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1042),
.B(n_929),
.Y(n_1075)
);

CKINVDCx16_ASAP7_75t_R g1076 ( 
.A(n_1008),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1033),
.B(n_967),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_1017),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_1013),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_988),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_1022),
.B(n_964),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_989),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_989),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_1009),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1034),
.A2(n_904),
.B1(n_954),
.B2(n_932),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_1058),
.Y(n_1086)
);

AO32x2_ASAP7_75t_L g1087 ( 
.A1(n_1043),
.A2(n_950),
.A3(n_954),
.B1(n_979),
.B2(n_903),
.Y(n_1087)
);

INVxp33_ASAP7_75t_SL g1088 ( 
.A(n_1045),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_990),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_997),
.A2(n_923),
.B1(n_963),
.B2(n_903),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1035),
.B(n_911),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1051),
.B(n_919),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_990),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_995),
.B(n_921),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_993),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1047),
.B(n_921),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_993),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_1011),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1044),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1041),
.B(n_962),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1058),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1011),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1059),
.A2(n_956),
.B(n_965),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1012),
.A2(n_972),
.B1(n_909),
.B2(n_878),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1063),
.A2(n_972),
.B1(n_909),
.B2(n_878),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1024),
.B(n_1019),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1050),
.B(n_966),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_1053),
.B(n_946),
.C(n_890),
.Y(n_1108)
);

CKINVDCx8_ASAP7_75t_R g1109 ( 
.A(n_1028),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1060),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1036),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_992),
.B(n_907),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1061),
.A2(n_972),
.B1(n_977),
.B2(n_905),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1027),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_994),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1030),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1014),
.B(n_914),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1039),
.B(n_888),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1026),
.B(n_897),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_1067),
.A2(n_953),
.A3(n_939),
.B(n_925),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1055),
.A2(n_905),
.B1(n_925),
.B2(n_987),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_SL g1122 ( 
.A(n_1020),
.B(n_913),
.C(n_879),
.Y(n_1122)
);

NOR4xp25_ASAP7_75t_L g1123 ( 
.A(n_1048),
.B(n_1001),
.C(n_1066),
.D(n_1046),
.Y(n_1123)
);

BUFx4f_ASAP7_75t_SL g1124 ( 
.A(n_995),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1032),
.B(n_984),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_999),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1054),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1037),
.B(n_975),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1023),
.B(n_973),
.Y(n_1129)
);

CKINVDCx16_ASAP7_75t_R g1130 ( 
.A(n_1029),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1004),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1038),
.B(n_926),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1025),
.B(n_968),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1080),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1085),
.A2(n_1005),
.B1(n_1052),
.B2(n_1016),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1082),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1083),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1089),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_L g1139 ( 
.A(n_1100),
.B(n_1031),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1093),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1095),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1097),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1115),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1091),
.B(n_1064),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1077),
.B(n_1057),
.Y(n_1145)
);

NOR2x1p5_ASAP7_75t_L g1146 ( 
.A(n_1068),
.B(n_1000),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1109),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1131),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1123),
.B(n_1021),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1079),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1103),
.B(n_1067),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1130),
.A2(n_1106),
.B1(n_1087),
.B2(n_1117),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1096),
.B(n_1065),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1092),
.B(n_1112),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1118),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1129),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1133),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1128),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1107),
.B(n_1062),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1119),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1101),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1078),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1125),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_L g1164 ( 
.A(n_1127),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1154),
.B(n_1076),
.Y(n_1165)
);

AND2x2_ASAP7_75t_SL g1166 ( 
.A(n_1159),
.B(n_1090),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1150),
.B(n_1111),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1155),
.B(n_1104),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1135),
.A2(n_1113),
.B1(n_1105),
.B2(n_998),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1134),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1144),
.B(n_1070),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1136),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1137),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1145),
.B(n_1075),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1148),
.B(n_1126),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1138),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_SL g1177 ( 
.A(n_1151),
.B(n_1071),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1160),
.B(n_1120),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1140),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1156),
.B(n_1132),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1153),
.B(n_1069),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1158),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1141),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1163),
.B(n_1122),
.Y(n_1184)
);

OAI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1135),
.A2(n_1006),
.B1(n_1003),
.B2(n_1049),
.C(n_1018),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1143),
.B(n_1121),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1142),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1177),
.B(n_1157),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_R g1189 ( 
.A(n_1170),
.B(n_1147),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1172),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1173),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1182),
.B(n_1151),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1182),
.B(n_1151),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1176),
.B(n_1152),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1179),
.B(n_1152),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1183),
.B(n_1143),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1187),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1178),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1184),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1180),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1180),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1190),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1199),
.A2(n_1185),
.B1(n_1149),
.B2(n_1168),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1191),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1197),
.Y(n_1205)
);

NAND4xp25_ASAP7_75t_L g1206 ( 
.A(n_1194),
.B(n_1184),
.C(n_1181),
.D(n_1168),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1196),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1200),
.B(n_1174),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1201),
.B(n_1171),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1194),
.B(n_1186),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1195),
.B(n_1186),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1188),
.B(n_1165),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1203),
.A2(n_1195),
.B(n_1149),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1202),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1202),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1206),
.A2(n_1166),
.B1(n_1169),
.B2(n_1188),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1210),
.A2(n_1192),
.B(n_1193),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1211),
.A2(n_1169),
.B1(n_1185),
.B2(n_1139),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1212),
.A2(n_1146),
.B(n_1147),
.C(n_1167),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1209),
.B(n_1162),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1214),
.Y(n_1221)
);

INVxp67_ASAP7_75t_SL g1222 ( 
.A(n_1215),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1213),
.A2(n_1204),
.B(n_1205),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1216),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1218),
.A2(n_1189),
.B(n_1188),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1224),
.Y(n_1226)
);

AOI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1223),
.A2(n_1225),
.B(n_1219),
.C(n_1217),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1221),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1222),
.B(n_1220),
.Y(n_1229)
);

XNOR2x2_ASAP7_75t_L g1230 ( 
.A(n_1223),
.B(n_1074),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1221),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1231),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1228),
.Y(n_1233)
);

AOI221x1_ASAP7_75t_SL g1234 ( 
.A1(n_1227),
.A2(n_1208),
.B1(n_1207),
.B2(n_1175),
.C(n_1198),
.Y(n_1234)
);

NOR3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1233),
.B(n_1162),
.C(n_1084),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1232),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1236),
.Y(n_1237)
);

NOR2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1237),
.B(n_1229),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_1238),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1238),
.Y(n_1240)
);

NAND4xp25_ASAP7_75t_L g1241 ( 
.A(n_1240),
.B(n_1234),
.C(n_1226),
.D(n_1102),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1239),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1242),
.B(n_1228),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1241),
.A2(n_1230),
.B1(n_1235),
.B2(n_1124),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1243),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1244),
.B(n_1161),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1245),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_1246),
.A2(n_1099),
.B1(n_1110),
.B2(n_1114),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1247),
.A2(n_1098),
.B1(n_1072),
.B2(n_999),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1248),
.B(n_1086),
.Y(n_1250)
);

OAI221xp5_ASAP7_75t_R g1251 ( 
.A1(n_1249),
.A2(n_1108),
.B1(n_1081),
.B2(n_1088),
.C(n_1010),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1250),
.A2(n_1116),
.B1(n_1150),
.B2(n_1094),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1251),
.B(n_1073),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1253),
.A2(n_1252),
.B1(n_1127),
.B2(n_1164),
.Y(n_1254)
);


endmodule