module fake_jpeg_5923_n_160 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_160);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_25),
.B1(n_23),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_27),
.B1(n_25),
.B2(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_26),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_17),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_13),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_28),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_17),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_67),
.Y(n_83)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_65),
.Y(n_88)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22x1_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_51),
.B1(n_41),
.B2(n_37),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_75),
.B(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_40),
.Y(n_92)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_32),
.C(n_34),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_34),
.C(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_57),
.Y(n_86)
);

OR2x6_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_31),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_46),
.B1(n_50),
.B2(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_24),
.B1(n_15),
.B2(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_80),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_24),
.B1(n_15),
.B2(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_86),
.B1(n_68),
.B2(n_69),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_70),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_104),
.B1(n_107),
.B2(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_69),
.B1(n_60),
.B2(n_73),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_60),
.C(n_68),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_99),
.C(n_97),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_61),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_83),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_71),
.B1(n_67),
.B2(n_56),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_119),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_115),
.A2(n_101),
.B1(n_100),
.B2(n_91),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_94),
.B(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_127),
.B(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_90),
.C(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_65),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_63),
.B1(n_42),
.B2(n_53),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_110),
.B1(n_113),
.B2(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_116),
.B1(n_112),
.B2(n_125),
.Y(n_144)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_127),
.B1(n_122),
.B2(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_141),
.B(n_132),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_120),
.B(n_124),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_123),
.C(n_121),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_143),
.C(n_145),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_40),
.C(n_24),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_141),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_139),
.A2(n_131),
.B1(n_10),
.B2(n_7),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_143),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_146),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_0),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_154),
.C(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_6),
.C(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_6),
.Y(n_160)
);


endmodule