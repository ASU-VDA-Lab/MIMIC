module fake_netlist_1_9924_n_624 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_624);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_624;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_18), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_62), .Y(n_74) );
HB1xp67_ASAP7_75t_L g75 ( .A(n_61), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_42), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_2), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_44), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_69), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_26), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_16), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_14), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_40), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_28), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_29), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_17), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
BUFx2_ASAP7_75t_L g91 ( .A(n_53), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_38), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_67), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_23), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_9), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_68), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_27), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_43), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_16), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_1), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_52), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_50), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_47), .B(n_58), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_39), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_63), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_14), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_51), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_60), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_18), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_110), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_110), .Y(n_121) );
OR2x2_ASAP7_75t_L g122 ( .A(n_111), .B(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_110), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_110), .Y(n_125) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_80), .B(n_72), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_91), .B(n_0), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_102), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_91), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_75), .B(n_3), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_102), .B(n_79), .Y(n_134) );
BUFx8_ASAP7_75t_L g135 ( .A(n_105), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_102), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_79), .B(n_32), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_111), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_87), .B(n_31), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_78), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_73), .B(n_3), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_85), .B(n_4), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_73), .B(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_93), .B(n_5), .Y(n_148) );
NAND2xp33_ASAP7_75t_R g149 ( .A(n_82), .B(n_35), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_85), .B(n_5), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_98), .B(n_6), .Y(n_152) );
OAI21x1_ASAP7_75t_L g153 ( .A1(n_87), .A2(n_37), .B(n_66), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_83), .B(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_103), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_104), .B(n_7), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_120), .B(n_100), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_120), .B(n_140), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_127), .Y(n_163) );
OR2x6_ASAP7_75t_L g164 ( .A(n_122), .B(n_108), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_135), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_119), .B(n_117), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
BUFx10_ASAP7_75t_L g172 ( .A(n_126), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_146), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_121), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVxp67_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_147), .B(n_117), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_119), .B(n_97), .Y(n_181) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_126), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_129), .B(n_108), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_129), .B(n_131), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_131), .B(n_106), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_147), .B(n_104), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_121), .B(n_100), .Y(n_192) );
INVx6_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_146), .B(n_88), .Y(n_195) );
OR2x6_ASAP7_75t_L g196 ( .A(n_122), .B(n_92), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_151), .B(n_84), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_118), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_123), .A2(n_77), .B1(n_84), .B2(n_88), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_151), .B(n_77), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_123), .B(n_92), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_118), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_118), .Y(n_203) );
AND3x4_ASAP7_75t_L g204 ( .A(n_126), .B(n_116), .C(n_109), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_132), .B(n_94), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_133), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_130), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_132), .B(n_101), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_193), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_206), .B(n_142), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_198), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_203), .Y(n_216) );
AND2x4_ASAP7_75t_SL g217 ( .A(n_172), .B(n_115), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_202), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_202), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_163), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_187), .B(n_137), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
OR2x6_ASAP7_75t_L g225 ( .A(n_193), .B(n_153), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_160), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_206), .B(n_141), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_158), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_174), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_187), .B(n_142), .Y(n_231) );
INVx5_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_212), .B(n_95), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_167), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_180), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_175), .B(n_138), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_175), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_178), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_161), .Y(n_241) );
BUFx4f_ASAP7_75t_SL g242 ( .A(n_159), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_197), .B(n_141), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_169), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_178), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_171), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_176), .B(n_156), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_168), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_177), .Y(n_252) );
INVxp67_ASAP7_75t_SL g253 ( .A(n_184), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_197), .B(n_138), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_179), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_189), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_211), .B(n_156), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_164), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_166), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_181), .B(n_155), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_208), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_181), .B(n_155), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_166), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_159), .B(n_125), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_164), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_168), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_182), .A2(n_134), .B1(n_136), .B2(n_154), .Y(n_269) );
NOR2xp67_ASAP7_75t_L g270 ( .A(n_194), .B(n_136), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_215), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_221), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_221), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_222), .B(n_194), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_215), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_250), .B(n_195), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_239), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_228), .B(n_190), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_239), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_250), .B(n_164), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_216), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_258), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_259), .B(n_196), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_238), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_228), .B(n_195), .Y(n_286) );
AO22x1_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_204), .B1(n_178), .B2(n_191), .Y(n_287) );
AOI222xp33_ASAP7_75t_L g288 ( .A1(n_242), .A2(n_182), .B1(n_162), .B2(n_200), .C1(n_183), .C2(n_172), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_237), .B(n_196), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_222), .B(n_200), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_248), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_248), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_218), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_248), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_243), .A2(n_178), .B1(n_191), .B2(n_204), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_216), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_214), .B(n_205), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_218), .Y(n_298) );
BUFx4_ASAP7_75t_SL g299 ( .A(n_227), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_237), .B(n_205), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_253), .A2(n_196), .B1(n_183), .B2(n_192), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_241), .A2(n_201), .B(n_210), .C(n_170), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_266), .B(n_201), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_225), .A2(n_207), .B(n_170), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_225), .A2(n_207), .B(n_153), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_226), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_241), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
INVx4_ASAP7_75t_L g310 ( .A(n_232), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_266), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_244), .Y(n_312) );
AOI22xp33_ASAP7_75t_SL g313 ( .A1(n_217), .A2(n_255), .B1(n_249), .B2(n_268), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_226), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_226), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_285), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_299), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_286), .B(n_247), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_304), .B(n_243), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_301), .A2(n_253), .B1(n_243), .B2(n_254), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_289), .A2(n_247), .B1(n_254), .B2(n_243), .Y(n_322) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_289), .A2(n_231), .B1(n_223), .B2(n_257), .C1(n_254), .C2(n_261), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
CKINVDCx6p67_ASAP7_75t_R g325 ( .A(n_272), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_297), .A2(n_261), .B(n_263), .C(n_233), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_231), .B1(n_223), .B2(n_254), .C1(n_263), .C2(n_217), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_279), .A2(n_267), .B1(n_246), .B2(n_244), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_277), .B(n_265), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
INVx6_ASAP7_75t_L g331 ( .A(n_310), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_309), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_295), .A2(n_267), .B1(n_252), .B2(n_256), .Y(n_333) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_304), .B(n_217), .Y(n_334) );
AOI22xp33_ASAP7_75t_SL g335 ( .A1(n_274), .A2(n_76), .B1(n_265), .B2(n_191), .Y(n_335) );
CKINVDCx6p67_ASAP7_75t_R g336 ( .A(n_284), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_271), .A2(n_256), .B1(n_252), .B2(n_246), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_281), .A2(n_245), .B1(n_225), .B2(n_270), .Y(n_338) );
CKINVDCx12_ASAP7_75t_R g339 ( .A(n_281), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_302), .A2(n_269), .B(n_225), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_293), .Y(n_341) );
OAI22xp5_ASAP7_75t_SL g342 ( .A1(n_313), .A2(n_96), .B1(n_199), .B2(n_225), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_287), .A2(n_199), .B1(n_201), .B2(n_152), .C(n_157), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_290), .A2(n_220), .B(n_219), .C(n_125), .Y(n_344) );
OAI22xp5_ASAP7_75t_SL g345 ( .A1(n_334), .A2(n_284), .B1(n_283), .B2(n_311), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_320), .A2(n_276), .B1(n_296), .B2(n_282), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g347 ( .A1(n_327), .A2(n_288), .B(n_277), .C(n_283), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_321), .B(n_271), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_329), .B(n_304), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_323), .A2(n_304), .B1(n_191), .B2(n_312), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_276), .B1(n_282), .B2(n_296), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_340), .A2(n_306), .B(n_225), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
AO221x2_ASAP7_75t_L g354 ( .A1(n_342), .A2(n_287), .B1(n_113), .B2(n_114), .C(n_112), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_329), .B(n_308), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_331), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_322), .A2(n_308), .B1(n_312), .B2(n_125), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_334), .A2(n_191), .B1(n_275), .B2(n_270), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_335), .A2(n_310), .B1(n_220), .B2(n_219), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_328), .A2(n_124), .B1(n_314), .B2(n_307), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_319), .A2(n_310), .B1(n_292), .B2(n_291), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_325), .A2(n_149), .B1(n_273), .B2(n_310), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_338), .A2(n_305), .B(n_128), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_321), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_326), .B(n_298), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_351), .A2(n_341), .B(n_337), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_357), .B(n_336), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
OA21x2_ASAP7_75t_L g374 ( .A1(n_352), .A2(n_341), .B(n_128), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_355), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_348), .B(n_321), .Y(n_376) );
INVx5_ASAP7_75t_SL g377 ( .A(n_348), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_347), .A2(n_343), .B1(n_316), .B2(n_332), .C(n_333), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_351), .A2(n_325), .B1(n_336), .B2(n_317), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_355), .Y(n_380) );
OA21x2_ASAP7_75t_L g381 ( .A1(n_369), .A2(n_128), .B(n_112), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_350), .A2(n_319), .B1(n_339), .B2(n_317), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_356), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_356), .B(n_319), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_361), .A2(n_344), .B1(n_331), .B2(n_113), .C(n_114), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_134), .B1(n_139), .B2(n_143), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_367), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_357), .B(n_298), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_346), .A2(n_124), .B1(n_136), .B2(n_150), .C(n_130), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_368), .B(n_105), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_298), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_367), .B(n_303), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_346), .A2(n_124), .B1(n_136), .B2(n_130), .C(n_107), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_367), .B(n_315), .Y(n_395) );
AO21x2_ASAP7_75t_L g396 ( .A1(n_366), .A2(n_315), .B(n_314), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_348), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_354), .B(n_74), .C(n_99), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_349), .B(n_315), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
INVx4_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
OAI21xp33_ASAP7_75t_SL g402 ( .A1(n_368), .A2(n_307), .B(n_303), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_383), .B(n_353), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_376), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_388), .B(n_354), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_377), .A2(n_354), .B1(n_345), .B2(n_363), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_401), .B(n_362), .Y(n_409) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_401), .B(n_360), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_390), .B(n_398), .C(n_378), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_380), .B(n_366), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_372), .B(n_345), .Y(n_414) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_379), .A2(n_365), .A3(n_363), .B1(n_359), .B2(n_358), .Y(n_415) );
OAI31xp33_ASAP7_75t_L g416 ( .A1(n_385), .A2(n_359), .A3(n_362), .B(n_358), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_382), .B(n_364), .C(n_8), .D(n_9), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_380), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_376), .B(n_366), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_400), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_397), .B(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_391), .B(n_134), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_373), .A2(n_273), .B1(n_307), .B2(n_303), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_397), .A2(n_166), .B(n_209), .C(n_188), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_384), .B(n_7), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_391), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_377), .A2(n_314), .B1(n_273), .B2(n_292), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
NOR3xp33_ASAP7_75t_L g431 ( .A(n_394), .B(n_294), .C(n_213), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_386), .B(n_166), .C(n_186), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_377), .B(n_8), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_387), .B(n_134), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g436 ( .A1(n_402), .A2(n_185), .B(n_188), .C(n_209), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_377), .A2(n_139), .B1(n_143), .B2(n_134), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_392), .B(n_10), .Y(n_438) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_387), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g441 ( .A(n_401), .B(n_371), .C(n_389), .Y(n_441) );
AOI31xp67_ASAP7_75t_L g442 ( .A1(n_403), .A2(n_264), .A3(n_236), .B(n_262), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_399), .A2(n_139), .B1(n_143), .B2(n_213), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_393), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_393), .B(n_11), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_403), .B(n_134), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_381), .A2(n_213), .B1(n_229), .B2(n_230), .C(n_294), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_396), .B(n_134), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_405), .B(n_396), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_440), .B(n_396), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_436), .A2(n_381), .B(n_374), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_423), .B(n_374), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_430), .B(n_381), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_404), .B(n_374), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_432), .B(n_374), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_412), .B(n_12), .Y(n_458) );
NAND4xp25_ASAP7_75t_SL g459 ( .A(n_408), .B(n_13), .C(n_15), .D(n_20), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_419), .B(n_13), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_408), .A2(n_139), .B1(n_143), .B2(n_134), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_417), .B(n_15), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_423), .B(n_186), .Y(n_463) );
AOI332xp33_ASAP7_75t_L g464 ( .A1(n_428), .A2(n_234), .A3(n_235), .B1(n_236), .B2(n_240), .B3(n_251), .C1(n_262), .C2(n_143), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_413), .B(n_209), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_422), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_421), .B(n_186), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_421), .B(n_186), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_439), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_411), .A2(n_139), .B(n_143), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_413), .B(n_209), .Y(n_471) );
AND4x1_ASAP7_75t_L g472 ( .A(n_416), .B(n_21), .C(n_22), .D(n_25), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_418), .A2(n_143), .B1(n_139), .B2(n_294), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_409), .B(n_280), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_448), .A2(n_188), .B(n_185), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_444), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_420), .B(n_188), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_445), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_409), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_442), .Y(n_480) );
NOR3xp33_ASAP7_75t_SL g481 ( .A(n_427), .B(n_143), .C(n_139), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_406), .A2(n_414), .B1(n_441), .B2(n_410), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_415), .B(n_291), .C(n_292), .D(n_251), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_434), .B(n_34), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_449), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_438), .B(n_185), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_449), .B(n_429), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_435), .B(n_41), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_441), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_446), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_435), .B(n_45), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_429), .B(n_426), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_446), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g495 ( .A1(n_447), .A2(n_273), .B(n_291), .C(n_294), .Y(n_495) );
OAI31xp33_ASAP7_75t_L g496 ( .A1(n_447), .A2(n_245), .A3(n_229), .B(n_230), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_425), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_46), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_431), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_437), .B(n_224), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_455), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_452), .A2(n_273), .B(n_229), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_469), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_456), .B(n_48), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_459), .A2(n_224), .B1(n_278), .B2(n_280), .Y(n_506) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_482), .A2(n_245), .A3(n_230), .B(n_56), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_490), .B(n_234), .C(n_262), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_476), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_469), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_479), .B(n_280), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_466), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_466), .Y(n_513) );
AOI21xp33_ASAP7_75t_SL g514 ( .A1(n_482), .A2(n_49), .B(n_55), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_453), .B(n_57), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_478), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_451), .B(n_64), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_458), .A2(n_236), .B(n_251), .C(n_240), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_462), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_493), .B(n_280), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_454), .B(n_65), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_488), .B(n_70), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_467), .B(n_224), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_465), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_457), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_460), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_467), .Y(n_527) );
NAND3x1_ASAP7_75t_L g528 ( .A(n_453), .B(n_280), .C(n_278), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_491), .B(n_224), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_468), .B(n_224), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_500), .A2(n_280), .B1(n_278), .B2(n_207), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_494), .B(n_240), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_450), .B(n_234), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_471), .B(n_235), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_471), .B(n_235), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_485), .B(n_264), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_485), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_500), .B(n_278), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_497), .B(n_278), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_264), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_487), .B(n_278), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_468), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_477), .B(n_232), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_484), .B(n_232), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_480), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_474), .B(n_232), .Y(n_547) );
AOI32xp33_ASAP7_75t_L g548 ( .A1(n_519), .A2(n_484), .A3(n_461), .B1(n_499), .B2(n_498), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_504), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_504), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_526), .B(n_484), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_509), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_510), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_525), .B(n_486), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_512), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_513), .B(n_472), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_543), .B(n_474), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_546), .Y(n_560) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_543), .B(n_461), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_547), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_524), .Y(n_563) );
XNOR2x2_ASAP7_75t_L g564 ( .A(n_515), .B(n_473), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_506), .A2(n_474), .B1(n_495), .B2(n_481), .Y(n_565) );
AOI31xp33_ASAP7_75t_SL g566 ( .A1(n_527), .A2(n_475), .A3(n_501), .B(n_464), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_540), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_505), .A2(n_483), .B1(n_470), .B2(n_499), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_537), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_533), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_528), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_514), .A2(n_489), .B1(n_492), .B2(n_496), .C(n_260), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_515), .B(n_492), .Y(n_574) );
XNOR2xp5_ASAP7_75t_L g575 ( .A(n_547), .B(n_489), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_508), .A2(n_232), .B(n_207), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_506), .A2(n_232), .B1(n_260), .B2(n_528), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_534), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_538), .A2(n_232), .B1(n_260), .B2(n_547), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_517), .B(n_260), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
OA22x2_ASAP7_75t_L g582 ( .A1(n_545), .A2(n_260), .B1(n_541), .B2(n_544), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_523), .B(n_530), .Y(n_583) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_507), .A2(n_511), .B(n_521), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_541), .Y(n_585) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_538), .B(n_522), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_529), .Y(n_587) );
OAI21xp5_ASAP7_75t_SL g588 ( .A1(n_531), .A2(n_518), .B(n_503), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_531), .A2(n_539), .B(n_532), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_539), .A2(n_459), .B(n_514), .C(n_379), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_542), .B(n_490), .C(n_482), .Y(n_591) );
AO22x2_ASAP7_75t_L g592 ( .A1(n_536), .A2(n_513), .B1(n_512), .B2(n_516), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_514), .A2(n_459), .B(n_379), .C(n_418), .Y(n_593) );
OAI221xp5_ASAP7_75t_SL g594 ( .A1(n_548), .A2(n_593), .B1(n_590), .B2(n_561), .C(n_568), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_592), .A2(n_582), .B(n_565), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_592), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_550), .B(n_553), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_558), .A2(n_552), .B1(n_591), .B2(n_568), .Y(n_598) );
XOR2x2_ASAP7_75t_L g599 ( .A(n_564), .B(n_575), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_558), .A2(n_584), .B(n_552), .C(n_562), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_549), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_586), .A2(n_571), .B1(n_583), .B2(n_559), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_588), .A2(n_572), .B(n_571), .C(n_549), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_583), .A2(n_570), .B1(n_581), .B2(n_578), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
INVx5_ASAP7_75t_L g606 ( .A(n_599), .Y(n_606) );
O2A1O1Ixp5_ASAP7_75t_L g607 ( .A1(n_594), .A2(n_555), .B(n_560), .C(n_567), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_596), .B(n_551), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_601), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g610 ( .A1(n_603), .A2(n_566), .B(n_577), .C(n_589), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_600), .A2(n_573), .B(n_576), .C(n_551), .Y(n_611) );
OAI211xp5_ASAP7_75t_SL g612 ( .A1(n_595), .A2(n_579), .B(n_556), .C(n_585), .Y(n_612) );
NOR2x2_ASAP7_75t_L g613 ( .A(n_606), .B(n_598), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_606), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_608), .Y(n_615) );
OAI322xp33_ASAP7_75t_L g616 ( .A1(n_611), .A2(n_597), .A3(n_554), .B1(n_587), .B2(n_569), .C1(n_574), .C2(n_563), .Y(n_616) );
OA21x2_ASAP7_75t_L g617 ( .A1(n_614), .A2(n_607), .B(n_609), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_615), .A2(n_606), .B1(n_612), .B2(n_610), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_618), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_617), .A2(n_613), .B1(n_597), .B2(n_616), .Y(n_620) );
NOR2xp67_ASAP7_75t_L g621 ( .A(n_619), .B(n_573), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_621), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_622), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_623), .A2(n_620), .B(n_580), .Y(n_624) );
endmodule