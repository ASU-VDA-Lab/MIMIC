module fake_aes_9711_n_484 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_484);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_484;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g66 ( .A(n_52), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_50), .Y(n_67) );
INVxp67_ASAP7_75t_L g68 ( .A(n_19), .Y(n_68) );
CKINVDCx16_ASAP7_75t_R g69 ( .A(n_31), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_27), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_55), .Y(n_71) );
INVx2_ASAP7_75t_L g72 ( .A(n_44), .Y(n_72) );
INVxp67_ASAP7_75t_SL g73 ( .A(n_60), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_51), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_21), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_48), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_29), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_20), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_63), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_11), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_17), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_37), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_33), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_26), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_30), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_62), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_3), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_54), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_1), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_6), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_6), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_46), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_53), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_2), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_10), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_13), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_56), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_66), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_66), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_75), .B(n_0), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_100), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_81), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_100), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_84), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_100), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_100), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
NOR2xp33_ASAP7_75t_R g120 ( .A(n_69), .B(n_34), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_83), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_68), .B(n_0), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_100), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_82), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_88), .B(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_74), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_94), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_76), .A2(n_36), .B(n_64), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_79), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_90), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_99), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_93), .B(n_4), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_132), .B(n_67), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_135), .B(n_85), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_138), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
OAI21xp33_ASAP7_75t_L g145 ( .A1(n_103), .A2(n_101), .B(n_78), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_135), .B(n_93), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_131), .B(n_86), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_138), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_135), .B(n_101), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_103), .B(n_78), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_104), .B(n_97), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_133), .B(n_91), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
AOI22x1_ASAP7_75t_L g168 ( .A1(n_104), .A2(n_137), .B1(n_136), .B2(n_134), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_133), .B(n_89), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_106), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_125), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_124), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_106), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_110), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_124), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_124), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_105), .B(n_92), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_107), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_126), .B(n_95), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_126), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_171), .Y(n_182) );
NOR2xp67_ASAP7_75t_L g183 ( .A(n_155), .B(n_105), .Y(n_183) );
INVx3_ASAP7_75t_SL g184 ( .A(n_141), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_179), .B(n_109), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
CKINVDCx8_ASAP7_75t_R g190 ( .A(n_161), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_179), .B(n_109), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_181), .B(n_121), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
BUFx4f_ASAP7_75t_SL g194 ( .A(n_161), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_181), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_141), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_178), .B(n_136), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_178), .B(n_134), .Y(n_201) );
O2A1O1Ixp5_ASAP7_75t_L g202 ( .A1(n_173), .A2(n_115), .B(n_129), .C(n_127), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_141), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_148), .B(n_139), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_130), .B(n_129), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_180), .B(n_119), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_164), .B(n_119), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_153), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
NOR2xp33_ASAP7_75t_R g211 ( .A(n_149), .B(n_112), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_174), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_141), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_178), .B(n_122), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_174), .Y(n_218) );
INVx5_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_170), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_170), .Y(n_223) );
NOR3xp33_ASAP7_75t_SL g224 ( .A(n_145), .B(n_127), .C(n_122), .Y(n_224) );
INVx5_ASAP7_75t_L g225 ( .A(n_149), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_180), .Y(n_226) );
AO22x1_ASAP7_75t_L g227 ( .A1(n_158), .A2(n_73), .B1(n_77), .B2(n_98), .Y(n_227) );
INVx6_ASAP7_75t_L g228 ( .A(n_147), .Y(n_228) );
NOR2xp33_ASAP7_75t_R g229 ( .A(n_149), .B(n_128), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_160), .B(n_115), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_207), .B(n_230), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_189), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_190), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_228), .Y(n_235) );
BUFx4_ASAP7_75t_SL g236 ( .A(n_198), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_184), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_200), .A2(n_217), .B(n_201), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_228), .Y(n_241) );
OR2x2_ASAP7_75t_SL g242 ( .A(n_192), .B(n_130), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_189), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_188), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_186), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_185), .B(n_160), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_191), .Y(n_249) );
NAND3xp33_ASAP7_75t_SL g250 ( .A(n_211), .B(n_120), .C(n_87), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_185), .B(n_160), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_199), .A2(n_166), .B(n_162), .C(n_147), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_185), .B(n_168), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_219), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
INVxp67_ASAP7_75t_SL g257 ( .A(n_186), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_194), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_193), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_187), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_198), .B(n_162), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_205), .B1(n_195), .B2(n_208), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_213), .A2(n_162), .B1(n_147), .B2(n_170), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_193), .B(n_147), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_193), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_193), .A2(n_170), .B1(n_166), .B2(n_175), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_210), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_219), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_216), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_246), .A2(n_249), .B1(n_263), .B2(n_231), .Y(n_273) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_253), .A2(n_206), .B(n_202), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_248), .B(n_183), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_261), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_233), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_233), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_240), .A2(n_183), .B(n_187), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_262), .B(n_227), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_234), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_264), .A2(n_197), .B1(n_224), .B2(n_203), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_248), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_265), .A2(n_219), .B1(n_209), .B2(n_215), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_236), .Y(n_285) );
INVx8_ASAP7_75t_L g286 ( .A(n_265), .Y(n_286) );
AOI211xp5_ASAP7_75t_L g287 ( .A1(n_250), .A2(n_229), .B(n_123), .C(n_96), .Y(n_287) );
AND2x2_ASAP7_75t_SL g288 ( .A(n_248), .B(n_218), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_244), .Y(n_289) );
OAI21xp33_ASAP7_75t_SL g290 ( .A1(n_244), .A2(n_204), .B(n_209), .Y(n_290) );
NAND2xp33_ASAP7_75t_R g291 ( .A(n_251), .B(n_196), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_245), .B(n_232), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_252), .B(n_212), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_251), .B(n_212), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_273), .B(n_268), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_279), .A2(n_253), .B(n_268), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g298 ( .A1(n_287), .A2(n_259), .B1(n_123), .B2(n_235), .C(n_241), .Y(n_298) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_291), .A2(n_267), .B(n_243), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_280), .A2(n_270), .B1(n_271), .B2(n_242), .Y(n_300) );
OAI22xp33_ASAP7_75t_SL g301 ( .A1(n_285), .A2(n_96), .B1(n_102), .B2(n_271), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_292), .A2(n_106), .B1(n_114), .B2(n_175), .C(n_215), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_276), .A2(n_114), .B1(n_204), .B2(n_222), .C(n_110), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_210), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_276), .B(n_225), .Y(n_305) );
OAI33xp33_ASAP7_75t_L g306 ( .A1(n_293), .A2(n_110), .A3(n_111), .B1(n_102), .B2(n_222), .B3(n_242), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_272), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_278), .Y(n_308) );
OAI21x1_ASAP7_75t_SL g309 ( .A1(n_278), .A2(n_173), .B(n_269), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_272), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_283), .A2(n_254), .B1(n_266), .B2(n_225), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_274), .A2(n_130), .B(n_111), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_283), .A2(n_225), .B1(n_223), .B2(n_220), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_285), .A2(n_237), .B1(n_239), .B2(n_238), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_289), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_295), .B(n_289), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_308), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_310), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_298), .B(n_290), .C(n_124), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_315), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_315), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_304), .Y(n_324) );
OAI31xp33_ASAP7_75t_L g325 ( .A1(n_301), .A2(n_275), .A3(n_282), .B(n_284), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_304), .B(n_288), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_306), .A2(n_275), .B1(n_294), .B2(n_286), .C(n_281), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_296), .B(n_288), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_310), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_312), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_312), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_307), .B(n_274), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_307), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_310), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g336 ( .A1(n_302), .A2(n_108), .B1(n_113), .B2(n_281), .C(n_223), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_310), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_300), .B(n_124), .C(n_113), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_311), .A2(n_257), .B1(n_237), .B2(n_247), .Y(n_340) );
OAI33xp33_ASAP7_75t_L g341 ( .A1(n_305), .A2(n_177), .A3(n_140), .B1(n_144), .B2(n_146), .B3(n_150), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_336), .A2(n_299), .B(n_297), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_323), .B(n_274), .Y(n_343) );
NOR3xp33_ASAP7_75t_L g344 ( .A(n_327), .B(n_314), .C(n_108), .Y(n_344) );
AOI322xp5_ASAP7_75t_L g345 ( .A1(n_318), .A2(n_4), .A3(n_5), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_10), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_325), .A2(n_313), .B1(n_303), .B2(n_309), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_323), .B(n_274), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_317), .B(n_130), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_318), .A2(n_108), .B1(n_124), .B2(n_173), .C(n_221), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_328), .B(n_7), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_321), .B(n_8), .Y(n_352) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_320), .B(n_143), .C(n_151), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_333), .B(n_143), .C(n_151), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_324), .B(n_12), .Y(n_355) );
AOI322xp5_ASAP7_75t_L g356 ( .A1(n_328), .A2(n_13), .A3(n_15), .B1(n_16), .B2(n_18), .C1(n_140), .C2(n_146), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_22), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_23), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_316), .B(n_25), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_316), .B(n_28), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_332), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_329), .B(n_218), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_330), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_335), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_326), .B(n_218), .Y(n_366) );
XOR2xp5_ASAP7_75t_L g367 ( .A(n_335), .B(n_256), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_319), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_326), .B(n_32), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
AOI221x1_ASAP7_75t_L g371 ( .A1(n_331), .A2(n_151), .B1(n_143), .B2(n_156), .C(n_172), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_218), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_337), .Y(n_374) );
NAND2xp33_ASAP7_75t_R g375 ( .A(n_337), .B(n_35), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_351), .B(n_337), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_351), .B(n_339), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_SL g378 ( .A1(n_345), .A2(n_338), .B(n_339), .C(n_340), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_373), .Y(n_380) );
INVx4_ASAP7_75t_L g381 ( .A(n_365), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_360), .B(n_38), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_365), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_360), .B(n_39), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_362), .B(n_40), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_364), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_362), .B(n_41), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_345), .B(n_167), .C(n_150), .D(n_146), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_343), .B(n_42), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_370), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_374), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_344), .A2(n_341), .B1(n_256), .B2(n_214), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_347), .B(n_43), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_347), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_45), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_369), .B(n_47), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_369), .B(n_49), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_366), .B(n_57), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_355), .B(n_58), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_358), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_348), .B(n_59), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_367), .B(n_61), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_348), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_357), .B(n_65), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_363), .B(n_140), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_358), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_389), .B(n_356), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_390), .A2(n_342), .B1(n_346), .B2(n_359), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_381), .B(n_353), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_397), .B(n_361), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_403), .A2(n_375), .B1(n_354), .B2(n_372), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_397), .B(n_342), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_406), .B(n_349), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_409), .B(n_367), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
AOI21xp5_ASAP7_75t_SL g421 ( .A1(n_387), .A2(n_371), .B(n_256), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_381), .A2(n_371), .B1(n_260), .B2(n_269), .Y(n_422) );
XOR2x2_ASAP7_75t_L g423 ( .A(n_381), .B(n_258), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
NAND3x2_ASAP7_75t_L g425 ( .A(n_394), .B(n_143), .C(n_176), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_392), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_379), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_379), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_260), .B1(n_258), .B2(n_255), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_376), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_399), .A2(n_260), .B1(n_255), .B2(n_220), .Y(n_434) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_400), .A2(n_163), .B(n_152), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_378), .A2(n_157), .B1(n_151), .B2(n_156), .C(n_143), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_411), .A2(n_410), .B1(n_396), .B2(n_391), .C(n_402), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_412), .A2(n_383), .B1(n_405), .B2(n_407), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_419), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_433), .B(n_382), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_413), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_416), .B(n_383), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_432), .B(n_382), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_417), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_415), .B(n_384), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_420), .B(n_398), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_420), .B(n_385), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_424), .B(n_385), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_427), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_424), .B(n_404), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_428), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_429), .B(n_404), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_425), .A2(n_387), .B1(n_407), .B2(n_401), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_436), .A2(n_408), .B(n_395), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_414), .A2(n_408), .B(n_151), .C(n_156), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_445), .B(n_431), .Y(n_457) );
NOR4xp25_ASAP7_75t_L g458 ( .A(n_442), .B(n_412), .C(n_435), .D(n_422), .Y(n_458) );
NAND3x1_ASAP7_75t_SL g459 ( .A(n_437), .B(n_423), .C(n_418), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_439), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_454), .A2(n_430), .B1(n_434), .B2(n_421), .Y(n_461) );
XNOR2x1_ASAP7_75t_L g462 ( .A(n_438), .B(n_423), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_456), .B(n_422), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_441), .B(n_450), .Y(n_464) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_460), .A2(n_453), .B1(n_451), .B2(n_444), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_463), .A2(n_447), .B1(n_451), .B2(n_452), .C1(n_449), .C2(n_448), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_457), .Y(n_467) );
NOR2xp33_ASAP7_75t_R g468 ( .A(n_459), .B(n_443), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_464), .Y(n_469) );
NOR2xp33_ASAP7_75t_R g470 ( .A(n_458), .B(n_440), .Y(n_470) );
NAND4xp75_ASAP7_75t_L g471 ( .A(n_458), .B(n_455), .C(n_448), .D(n_449), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_462), .A2(n_446), .B1(n_455), .B2(n_172), .Y(n_472) );
OA22x2_ASAP7_75t_L g473 ( .A1(n_460), .A2(n_442), .B1(n_438), .B2(n_461), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_473), .A2(n_471), .B1(n_465), .B2(n_469), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_470), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_467), .B(n_466), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_468), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_475), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_476), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_478), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_479), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_480), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_482), .A2(n_474), .B1(n_479), .B2(n_481), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_483), .A2(n_477), .B(n_472), .Y(n_484) );
endmodule