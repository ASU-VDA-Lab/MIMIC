module fake_netlist_1_1263_n_688 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_688);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_688;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g77 ( .A(n_66), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_56), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_31), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_45), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_6), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_40), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_53), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_26), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_74), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_33), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_55), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_27), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_36), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_38), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_64), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_57), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_52), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_70), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_42), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_19), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_17), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_2), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_23), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_21), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_28), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_54), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_43), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_32), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_7), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_68), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_12), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_10), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_47), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_46), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_119), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_109), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_109), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_77), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_105), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_105), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_116), .Y(n_134) );
NOR2xp33_ASAP7_75t_R g135 ( .A(n_96), .B(n_76), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_80), .B(n_75), .Y(n_136) );
INVx5_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_120), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
NOR2xp33_ASAP7_75t_R g140 ( .A(n_80), .B(n_73), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_77), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_107), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_83), .B(n_0), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_115), .B(n_1), .Y(n_146) );
NOR2xp33_ASAP7_75t_R g147 ( .A(n_84), .B(n_72), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_110), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_79), .B(n_1), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_83), .B(n_2), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_123), .Y(n_156) );
NOR2xp67_ASAP7_75t_L g157 ( .A(n_118), .B(n_3), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_85), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_118), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_114), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_106), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_118), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_84), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_118), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_97), .B(n_3), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_118), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_160), .B(n_117), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_128), .B(n_97), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_127), .B(n_121), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_164), .Y(n_173) );
INVx3_ASAP7_75t_R g174 ( .A(n_166), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_127), .A2(n_118), .B1(n_78), .B2(n_82), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_133), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_146), .B(n_121), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_161), .B(n_124), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_163), .B(n_122), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_160), .B(n_122), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_126), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_153), .B(n_98), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_129), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_158), .B(n_124), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_136), .B(n_113), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_163), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_130), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_142), .A2(n_113), .B1(n_112), .B2(n_111), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_142), .A2(n_112), .B1(n_111), .B2(n_104), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
AND2x6_ASAP7_75t_L g213 ( .A(n_152), .B(n_94), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_140), .B(n_104), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_151), .A2(n_103), .B1(n_102), .B2(n_101), .Y(n_215) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_152), .B(n_103), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_134), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_125), .B(n_102), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_139), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_143), .B(n_101), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_148), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g224 ( .A1(n_151), .A2(n_100), .B1(n_99), .B2(n_98), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_134), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_144), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_134), .B(n_100), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_145), .B(n_99), .Y(n_228) );
INVx4_ASAP7_75t_L g229 ( .A(n_145), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_225), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_226), .B(n_165), .Y(n_233) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_182), .A2(n_147), .B(n_155), .Y(n_234) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_213), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_198), .B(n_145), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_196), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_173), .Y(n_238) );
NOR2xp33_ASAP7_75t_R g239 ( .A(n_180), .B(n_162), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_219), .B(n_162), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_198), .B(n_159), .Y(n_242) );
AND3x1_ASAP7_75t_SL g243 ( .A(n_180), .B(n_133), .C(n_87), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_200), .B(n_135), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_191), .A2(n_219), .B1(n_222), .B2(n_185), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_189), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_224), .B(n_86), .C(n_87), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_212), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_168), .Y(n_253) );
NAND2xp33_ASAP7_75t_SL g254 ( .A(n_200), .B(n_159), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_172), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_219), .B(n_157), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_222), .B(n_92), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_188), .B(n_92), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_179), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_183), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_210), .B(n_86), .C(n_88), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_187), .B(n_88), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_179), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_181), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_215), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_216), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_175), .A2(n_93), .B(n_90), .C(n_95), .Y(n_267) );
CKINVDCx14_ASAP7_75t_R g268 ( .A(n_209), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_216), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_172), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_167), .Y(n_271) );
INVx6_ASAP7_75t_L g272 ( .A(n_225), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_178), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
NOR3xp33_ASAP7_75t_SL g277 ( .A(n_195), .B(n_90), .C(n_91), .Y(n_277) );
NOR2xp33_ASAP7_75t_R g278 ( .A(n_167), .B(n_91), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_195), .B(n_177), .C(n_171), .Y(n_280) );
NAND2xp33_ASAP7_75t_SL g281 ( .A(n_200), .B(n_95), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_206), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_194), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_225), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_194), .Y(n_286) );
NOR2xp33_ASAP7_75t_R g287 ( .A(n_197), .B(n_93), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_229), .B(n_94), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g289 ( .A(n_191), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_201), .B(n_169), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_191), .A2(n_89), .B1(n_149), .B2(n_150), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_223), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_193), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_193), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_229), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_233), .A2(n_201), .B(n_182), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_239), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_268), .A2(n_190), .B1(n_186), .B2(n_184), .C(n_187), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_266), .B(n_229), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_230), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_232), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_290), .A2(n_214), .B(n_227), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_262), .B(n_191), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
BUFx4_ASAP7_75t_SL g306 ( .A(n_250), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_262), .B(n_191), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_232), .Y(n_308) );
BUFx4f_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_236), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_231), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_269), .B(n_218), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_236), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_262), .B(n_191), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_237), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_267), .A2(n_214), .B(n_218), .C(n_228), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_255), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_272), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_248), .B(n_228), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_236), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_289), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_249), .B(n_218), .Y(n_325) );
INVx3_ASAP7_75t_SL g326 ( .A(n_250), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_238), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_241), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_265), .A2(n_228), .B1(n_213), .B2(n_197), .C1(n_89), .C2(n_221), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_271), .A2(n_197), .B1(n_213), .B2(n_221), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_244), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_230), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_242), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_249), .B(n_213), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_242), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_271), .A2(n_197), .B1(n_213), .B2(n_199), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_245), .B(n_197), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_242), .B(n_89), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_265), .A2(n_197), .B1(n_213), .B2(n_199), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_252), .B(n_211), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_252), .B(n_207), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_244), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_260), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_281), .A2(n_211), .B(n_207), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_241), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_240), .A2(n_207), .B1(n_150), .B2(n_6), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_332), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_338), .A2(n_278), .B(n_251), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_311), .B(n_283), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_313), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_311), .B(n_283), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_298), .A2(n_280), .B1(n_261), .B2(n_260), .C(n_257), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_312), .B(n_292), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_292), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_235), .B1(n_258), .B2(n_247), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_308), .A2(n_277), .B1(n_256), .B2(n_247), .C(n_288), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_317), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_308), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_317), .Y(n_362) );
NAND2x1_ASAP7_75t_L g363 ( .A(n_332), .B(n_272), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
INVx4_ASAP7_75t_L g365 ( .A(n_309), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_343), .A2(n_254), .B1(n_243), .B2(n_295), .C(n_279), .Y(n_366) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_310), .B(n_287), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_322), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_309), .A2(n_235), .B1(n_291), .B2(n_256), .Y(n_370) );
NAND3xp33_ASAP7_75t_SL g371 ( .A(n_318), .B(n_282), .C(n_279), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_319), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
NAND3xp33_ASAP7_75t_SL g374 ( .A(n_301), .B(n_282), .C(n_276), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_297), .A2(n_256), .B1(n_235), .B2(n_234), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_328), .B(n_285), .Y(n_376) );
AOI21xp5_ASAP7_75t_SL g377 ( .A1(n_338), .A2(n_255), .B(n_270), .Y(n_377) );
NOR2x1_ASAP7_75t_SL g378 ( .A(n_338), .B(n_274), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_349), .B(n_328), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_354), .A2(n_345), .B(n_303), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_349), .B(n_345), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_333), .B1(n_335), .B2(n_346), .C(n_321), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_350), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_338), .B1(n_315), .B2(n_310), .Y(n_384) );
AO21x2_ASAP7_75t_L g385 ( .A1(n_371), .A2(n_296), .B(n_307), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_361), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_329), .B(n_234), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_352), .B(n_325), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_359), .A2(n_304), .B(n_316), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_357), .A2(n_339), .B(n_336), .C(n_330), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_352), .B(n_325), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_348), .A2(n_315), .B1(n_323), .B2(n_234), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_362), .A2(n_323), .B1(n_297), .B2(n_334), .Y(n_395) );
BUFx4f_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_366), .B(n_314), .C(n_341), .D(n_324), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_362), .A2(n_342), .B(n_327), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_334), .B1(n_342), .B2(n_331), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_331), .B1(n_299), .B2(n_324), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_369), .A2(n_299), .B1(n_324), .B2(n_340), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_355), .A2(n_299), .B1(n_305), .B2(n_300), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_375), .A2(n_326), .B1(n_314), .B2(n_341), .C(n_300), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_347), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_355), .A2(n_326), .B1(n_300), .B2(n_305), .Y(n_406) );
CKINVDCx11_ASAP7_75t_R g407 ( .A(n_386), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_404), .A2(n_365), .B1(n_373), .B2(n_378), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_395), .A2(n_306), .B(n_377), .C(n_360), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_404), .A2(n_365), .B1(n_373), .B2(n_347), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_405), .Y(n_411) );
NOR2xp33_ASAP7_75t_R g412 ( .A(n_383), .B(n_367), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_379), .B(n_351), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_382), .A2(n_356), .B1(n_374), .B2(n_370), .C(n_373), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_373), .B1(n_365), .B2(n_370), .C(n_347), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_394), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_405), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_384), .A2(n_365), .B1(n_377), .B2(n_358), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
NOR2xp33_ASAP7_75t_R g420 ( .A(n_396), .B(n_360), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_402), .A2(n_376), .B(n_344), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_379), .B(n_351), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_384), .A2(n_358), .B1(n_364), .B2(n_351), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
AOI211xp5_ASAP7_75t_SL g425 ( .A1(n_400), .A2(n_360), .B(n_376), .C(n_364), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_379), .B(n_364), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_381), .B(n_358), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_394), .B(n_372), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_397), .B(n_337), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_400), .A2(n_363), .B1(n_305), .B2(n_372), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_402), .A2(n_378), .B(n_363), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_381), .B(n_372), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_393), .B(n_150), .C(n_319), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_381), .B(n_337), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_396), .B(n_319), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_389), .A2(n_320), .B1(n_337), .B2(n_276), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_398), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_397), .A2(n_320), .B1(n_319), .B2(n_295), .Y(n_442) );
OAI21x1_ASAP7_75t_L g443 ( .A1(n_434), .A2(n_393), .B(n_398), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_419), .B(n_401), .Y(n_444) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_420), .A2(n_388), .B(n_406), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_426), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_426), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_419), .B(n_401), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_441), .B(n_396), .Y(n_449) );
AOI33xp33_ASAP7_75t_L g450 ( .A1(n_424), .A2(n_395), .A3(n_406), .B1(n_392), .B2(n_399), .B3(n_9), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_441), .Y(n_451) );
OAI31xp33_ASAP7_75t_L g452 ( .A1(n_409), .A2(n_403), .A3(n_391), .B(n_392), .Y(n_452) );
AND2x4_ASAP7_75t_SL g453 ( .A(n_413), .B(n_392), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_440), .A2(n_403), .B1(n_398), .B2(n_399), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_436), .A2(n_388), .B1(n_391), .B2(n_390), .C(n_396), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_398), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_417), .Y(n_457) );
NAND3xp33_ASAP7_75t_SL g458 ( .A(n_412), .B(n_4), .C(n_5), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_415), .A2(n_390), .B1(n_150), .B2(n_385), .C(n_294), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_413), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_417), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_422), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_438), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_427), .B(n_380), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_438), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_430), .A2(n_414), .B1(n_442), .B2(n_423), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_433), .B(n_390), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_390), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_434), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_428), .B(n_380), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_429), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_429), .B(n_380), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_411), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_411), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_408), .A2(n_380), .B1(n_285), .B2(n_293), .C(n_294), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_418), .B(n_380), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_425), .B(n_385), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_425), .B(n_385), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_435), .B(n_385), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_410), .B(n_246), .C(n_293), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_432), .B(n_319), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_421), .B(n_439), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_439), .B(n_150), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_407), .Y(n_488) );
OAI222xp33_ASAP7_75t_L g489 ( .A1(n_431), .A2(n_4), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_10), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_426), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_426), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_460), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_456), .B(n_8), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_460), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_466), .B(n_11), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_466), .B(n_12), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_464), .B(n_13), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_464), .B(n_13), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_466), .B(n_14), .Y(n_504) );
NOR4xp25_ASAP7_75t_SL g505 ( .A(n_478), .B(n_14), .C(n_15), .D(n_16), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_448), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_446), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_446), .Y(n_508) );
AOI21xp33_ASAP7_75t_SL g509 ( .A1(n_449), .A2(n_15), .B(n_16), .Y(n_509) );
OAI21xp33_ASAP7_75t_SL g510 ( .A1(n_449), .A2(n_18), .B(n_19), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_453), .B(n_18), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_461), .B(n_69), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_447), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_20), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_482), .B(n_20), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_492), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_492), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_447), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_461), .B(n_37), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_473), .B(n_21), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_467), .B(n_264), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g524 ( .A1(n_458), .A2(n_285), .B(n_24), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_474), .B(n_22), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_453), .B(n_29), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_474), .B(n_30), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_469), .A2(n_272), .B1(n_259), .B2(n_263), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_447), .Y(n_529) );
NAND2xp33_ASAP7_75t_SL g530 ( .A(n_467), .B(n_34), .Y(n_530) );
NOR2xp67_ASAP7_75t_SL g531 ( .A(n_478), .B(n_272), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_467), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_490), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_461), .B(n_35), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_451), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_473), .B(n_470), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_491), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_486), .A2(n_264), .B1(n_263), .B2(n_259), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_451), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
NAND2xp33_ASAP7_75t_R g543 ( .A(n_493), .B(n_39), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_470), .B(n_44), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_471), .B(n_49), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_462), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_471), .B(n_51), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_462), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_451), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_468), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_468), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_537), .B(n_538), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_497), .B(n_474), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_524), .A2(n_453), .B1(n_449), .B2(n_469), .Y(n_554) );
AOI222xp33_ASAP7_75t_L g555 ( .A1(n_510), .A2(n_458), .B1(n_489), .B2(n_488), .C1(n_486), .C2(n_455), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_509), .A2(n_489), .B(n_488), .C(n_445), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_513), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_511), .A2(n_454), .B(n_457), .C(n_445), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_542), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_537), .B(n_475), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_507), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_507), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_497), .B(n_468), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_530), .A2(n_450), .B(n_487), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_543), .A2(n_454), .B1(n_463), .B2(n_465), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_513), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_498), .B(n_463), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_502), .B(n_457), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_495), .A2(n_463), .B1(n_465), .B2(n_457), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g571 ( .A1(n_498), .A2(n_481), .B(n_480), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_504), .B(n_465), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_519), .Y(n_573) );
AOI322xp5_ASAP7_75t_L g574 ( .A1(n_504), .A2(n_455), .A3(n_459), .B1(n_487), .B2(n_472), .C1(n_475), .C2(n_481), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_503), .A2(n_487), .B1(n_459), .B2(n_452), .C(n_480), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_530), .B(n_514), .C(n_515), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_533), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_514), .B(n_457), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_515), .A2(n_476), .B1(n_484), .B2(n_477), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_521), .B(n_477), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_521), .B(n_477), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_508), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_495), .A2(n_452), .B(n_472), .C(n_485), .Y(n_585) );
AOI221xp5_ASAP7_75t_SL g586 ( .A1(n_522), .A2(n_479), .B1(n_485), .B2(n_484), .C(n_476), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_523), .A2(n_526), .B(n_544), .C(n_547), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_516), .Y(n_588) );
OAI22x1_ASAP7_75t_L g589 ( .A1(n_539), .A2(n_476), .B1(n_479), .B2(n_484), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_517), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_512), .A2(n_443), .B(n_476), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_512), .A2(n_443), .B(n_483), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_518), .B(n_443), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_517), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_544), .A2(n_483), .B1(n_273), .B2(n_176), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_518), .B(n_59), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_500), .B(n_61), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g598 ( .A1(n_501), .A2(n_273), .A3(n_62), .B1(n_204), .B2(n_205), .C1(n_217), .C2(n_176), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_506), .B(n_204), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_494), .Y(n_600) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_505), .B(n_536), .C(n_539), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_578), .B(n_548), .Y(n_602) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_577), .B(n_547), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_552), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_554), .A2(n_520), .B(n_512), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_560), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_560), .B(n_546), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g608 ( .A1(n_566), .A2(n_531), .B(n_545), .C(n_534), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_562), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g610 ( .A(n_557), .B(n_531), .C(n_494), .Y(n_610) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_566), .B(n_520), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_558), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_561), .B(n_564), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_563), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_575), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_565), .A2(n_520), .B1(n_534), .B2(n_527), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_583), .Y(n_617) );
NOR2xp33_ASAP7_75t_R g618 ( .A(n_595), .B(n_525), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_553), .B(n_551), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_584), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_570), .B(n_534), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_556), .B(n_601), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_555), .B(n_540), .C(n_528), .D(n_550), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_568), .B(n_551), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_570), .B(n_525), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_569), .B(n_550), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_590), .B(n_496), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_594), .B(n_499), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_582), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_579), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_558), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_587), .A2(n_527), .B(n_541), .C(n_549), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
NOR3x1_ASAP7_75t_L g637 ( .A(n_593), .B(n_549), .C(n_541), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_622), .B(n_569), .Y(n_638) );
XOR2xp5_ASAP7_75t_L g639 ( .A(n_603), .B(n_572), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_613), .B(n_581), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_611), .A2(n_559), .B(n_589), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_606), .Y(n_642) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_637), .A2(n_559), .B1(n_586), .B2(n_599), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_622), .A2(n_585), .B(n_595), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_632), .B(n_574), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_610), .A2(n_592), .B(n_571), .Y(n_646) );
XNOR2xp5_ASAP7_75t_L g647 ( .A(n_604), .B(n_580), .Y(n_647) );
AOI221xp5_ASAP7_75t_SL g648 ( .A1(n_624), .A2(n_576), .B1(n_591), .B2(n_599), .C(n_597), .Y(n_648) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_608), .A2(n_596), .B(n_573), .Y(n_649) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_605), .B(n_598), .C(n_535), .D(n_529), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_607), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_625), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_602), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_630), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_619), .Y(n_655) );
O2A1O1Ixp5_ASAP7_75t_L g656 ( .A1(n_621), .A2(n_529), .B(n_519), .C(n_217), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_634), .A2(n_286), .B(n_270), .C(n_217), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_612), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_651), .Y(n_659) );
NAND3x1_ASAP7_75t_SL g660 ( .A(n_644), .B(n_626), .C(n_616), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_638), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_641), .A2(n_627), .B(n_616), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_645), .B(n_631), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_638), .A2(n_617), .B1(n_623), .B2(n_620), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_639), .B(n_614), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_654), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_656), .A2(n_615), .B(n_609), .C(n_628), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_642), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_658), .Y(n_669) );
AOI21xp33_ASAP7_75t_SL g670 ( .A1(n_643), .A2(n_618), .B(n_629), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_648), .A2(n_636), .B1(n_635), .B2(n_633), .C(n_618), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_652), .A2(n_205), .B1(n_274), .B2(n_275), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_275), .B(n_284), .C(n_286), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_655), .B(n_653), .Y(n_674) );
OA22x2_ASAP7_75t_L g675 ( .A1(n_647), .A2(n_275), .B1(n_284), .B2(n_658), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_649), .A2(n_284), .B1(n_650), .B2(n_640), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_670), .A2(n_662), .B1(n_676), .B2(n_675), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_661), .B(n_671), .Y(n_678) );
OR3x2_ASAP7_75t_L g679 ( .A(n_660), .B(n_659), .C(n_666), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_674), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_677), .B(n_663), .C(n_656), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_679), .A2(n_663), .B1(n_665), .B2(n_668), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_680), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_683), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_681), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_682), .B1(n_677), .B2(n_678), .C(n_667), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_684), .B1(n_685), .B2(n_664), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_672), .B1(n_673), .B2(n_657), .C(n_669), .Y(n_688) );
endmodule