module real_jpeg_17136_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI32xp33_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_22),
.A3(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_21)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_0),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_0),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_0),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_0),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_0),
.A2(n_181),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_89),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_2),
.A2(n_89),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_2),
.A2(n_89),
.B1(n_235),
.B2(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_3),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_3),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_4),
.A2(n_130),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_4),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_5),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_5),
.Y(n_302)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_6),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_8),
.Y(n_209)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_8),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_320),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_267),
.B(n_315),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_214),
.B(n_266),
.Y(n_15)
);

AOI21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_190),
.B(n_213),
.Y(n_16)
);

OAI21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_138),
.B(n_189),
.Y(n_17)
);

NOR2xp67_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_19),
.B(n_124),
.Y(n_189)
);

XOR2x2_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_61),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_20),
.B(n_93),
.C(n_122),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_21),
.B(n_40),
.Y(n_193)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_29),
.A2(n_285),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_34),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_72)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_41),
.A2(n_128),
.B1(n_129),
.B2(n_134),
.Y(n_127)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_42),
.B(n_50),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_43),
.A2(n_95),
.B(n_98),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_45),
.A2(n_107),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_45),
.Y(n_170)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_45),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_48),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_49),
.B(n_299),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_53),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_57),
.A2(n_129),
.B(n_177),
.Y(n_176)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_60),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_93),
.B1(n_122),
.B2(n_123),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_62),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_62),
.A2(n_122),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_62),
.A2(n_122),
.B1(n_274),
.B2(n_275),
.Y(n_347)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_72),
.B1(n_78),
.B2(n_85),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_63),
.A2(n_72),
.B1(n_78),
.B2(n_85),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_63),
.A2(n_72),
.B(n_78),
.Y(n_313)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_70),
.Y(n_207)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_71),
.Y(n_260)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_92),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_93),
.A2(n_123),
.B1(n_141),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_93),
.A2(n_123),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_93),
.B(n_281),
.Y(n_310)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_101),
.B1(n_111),
.B2(n_116),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_101),
.B1(n_111),
.B2(n_116),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_94),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_94),
.B(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_142),
.A3(n_146),
.B1(n_148),
.B2(n_153),
.Y(n_141)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_101),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_101),
.Y(n_341)
);

NOR2x1p5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_105),
.Y(n_339)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_113),
.Y(n_305)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_122),
.B(n_220),
.C(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_136),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_126),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_125),
.B(n_193),
.C(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_125),
.A2(n_126),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_126),
.B(n_298),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_179),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_127),
.A2(n_160),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_128),
.A2(n_282),
.B1(n_299),
.B2(n_306),
.Y(n_298)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21x1_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_163),
.B(n_188),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_159),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_SL g188 ( 
.A(n_140),
.B(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_160),
.B(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_183),
.B(n_187),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_178),
.B(n_182),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_170),
.Y(n_284)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_184),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_197),
.C(n_201),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_177),
.A2(n_282),
.B(n_286),
.Y(n_281)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_181),
.B(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_212),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_212),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_211),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_210),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_197),
.A2(n_210),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_197),
.B(n_274),
.C(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_226),
.B1(n_233),
.B2(n_243),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_234),
.B(n_239),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_203),
.A2(n_226),
.B1(n_233),
.B2(n_243),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_216),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_247),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_248),
.C(n_249),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B(n_223),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_222),
.A2(n_334),
.B(n_340),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_224),
.A2(n_225),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_225),
.Y(n_328)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_292),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_271),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_279),
.C(n_289),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_274),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_289),
.B2(n_290),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_318),
.Y(n_317)
);

NAND2x1_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_314),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_314),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_309),
.C(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_309),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_312),
.C(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_348),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_325),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_345),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_342),
.B2(n_344),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_342),
.Y(n_344)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);


endmodule