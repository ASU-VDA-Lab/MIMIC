module real_jpeg_1645_n_22 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_22);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_22;

wire n_43;
wire n_57;
wire n_37;
wire n_54;
wire n_73;
wire n_65;
wire n_38;
wire n_33;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_69;
wire n_58;
wire n_52;
wire n_31;
wire n_67;
wire n_49;
wire n_63;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_51;
wire n_47;
wire n_45;
wire n_61;
wire n_25;
wire n_71;
wire n_42;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_70;
wire n_74;
wire n_27;
wire n_26;
wire n_41;
wire n_32;
wire n_30;
wire n_56;
wire n_48;

AOI221xp5_ASAP7_75t_L g25 ( 
.A1(n_0),
.A2(n_13),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_73),
.B2(n_74),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_1),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI321xp33_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_4),
.A3(n_41),
.B1(n_42),
.B2(n_43),
.C(n_45),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_3),
.B1(n_4),
.B2(n_18),
.Y(n_72)
);

AOI222xp33_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_7),
.B1(n_18),
.B2(n_37),
.C1(n_38),
.C2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_4),
.B(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_13),
.B(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_12),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_9),
.B1(n_39),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_9),
.A3(n_17),
.B1(n_21),
.B2(n_58),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

NAND5xp2_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_10),
.C(n_14),
.D(n_20),
.E(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

OAI211xp5_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_17),
.B(n_55),
.C(n_58),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

AOI31xp33_ASAP7_75t_L g60 ( 
.A1(n_12),
.A2(n_19),
.A3(n_61),
.B(n_68),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_19),
.A3(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_24),
.A3(n_40),
.B1(n_50),
.B2(n_53),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_15),
.A2(n_36),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

OAI321xp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_25),
.A3(n_31),
.B1(n_33),
.B2(n_35),
.C(n_36),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_32),
.B(n_34),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_19),
.A2(n_61),
.B(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_64),
.Y(n_63)
);

OAI221xp5_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.C(n_67),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_30),
.B(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_42),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_41),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_59),
.Y(n_58)
);

NAND4xp25_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.C(n_48),
.D(n_49),
.Y(n_45)
);

OAI322xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.A3(n_60),
.B1(n_69),
.B2(n_70),
.C1(n_71),
.C2(n_72),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);


endmodule