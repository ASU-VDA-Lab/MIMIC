module fake_netlist_6_3759_n_1072 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1072);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1072;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_923;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_843;
wire n_656;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_964;
wire n_982;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_1001;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g182 ( 
.A(n_34),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_107),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_87),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_41),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_145),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_78),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_73),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_45),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_19),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_104),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_61),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_58),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_49),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_128),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_40),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_132),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_64),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_171),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_175),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_56),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_16),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_57),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_131),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_20),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_137),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_72),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_25),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_105),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_154),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_179),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_42),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_52),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_125),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_90),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_172),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_115),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_170),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_25),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_62),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_92),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_75),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_103),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_109),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_178),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_27),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_9),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_196),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

BUFx2_ASAP7_75t_SL g273 ( 
.A(n_197),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_247),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_198),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_186),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_201),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_182),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_184),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_192),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_209),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_213),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_210),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_231),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_183),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_183),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_185),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_257),
.A2(n_188),
.B(n_187),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_255),
.A2(n_249),
.B1(n_207),
.B2(n_248),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_254),
.A2(n_232),
.B(n_190),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_284),
.A2(n_224),
.B1(n_246),
.B2(n_245),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_189),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_191),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_266),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_258),
.A2(n_195),
.B(n_194),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_266),
.B(n_199),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

AOI22x1_ASAP7_75t_SL g325 ( 
.A1(n_275),
.A2(n_287),
.B1(n_274),
.B2(n_299),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_293),
.A2(n_302),
.B1(n_299),
.B2(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_261),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_250),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_302),
.A2(n_263),
.B1(n_265),
.B2(n_282),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_267),
.Y(n_334)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_266),
.B(n_33),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_L g338 ( 
.A(n_281),
.B(n_200),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_202),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_284),
.A2(n_298),
.B1(n_256),
.B2(n_265),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_268),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_295),
.B(n_35),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_268),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

AOI22x1_ASAP7_75t_SL g348 ( 
.A1(n_274),
.A2(n_244),
.B1(n_242),
.B2(n_239),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_295),
.A2(n_204),
.B(n_203),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_278),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_211),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_279),
.A2(n_238),
.B1(n_236),
.B2(n_235),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_301),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_333),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_262),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_317),
.B(n_300),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_305),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_305),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_355),
.B(n_212),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_341),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_355),
.B(n_214),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_L g373 ( 
.A(n_310),
.B(n_338),
.C(n_339),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

NOR2x1p5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_300),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_348),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_356),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_215),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_314),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_223),
.C(n_220),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_304),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_320),
.B(n_226),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_229),
.C(n_228),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_328),
.B(n_278),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_230),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_325),
.B(n_273),
.Y(n_408)
);

BUFx6f_ASAP7_75t_SL g409 ( 
.A(n_331),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_L g411 ( 
.A(n_335),
.B(n_233),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_353),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_348),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_320),
.B(n_315),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_313),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_353),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_234),
.C(n_273),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_315),
.B(n_0),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_323),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_323),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_315),
.B(n_36),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_325),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_373),
.B(n_316),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_361),
.B(n_316),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_430),
.B(n_316),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_379),
.B(n_309),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_318),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_374),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

OR2x2_ASAP7_75t_SL g446 ( 
.A(n_422),
.B(n_309),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_425),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_377),
.B(n_312),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_R g450 ( 
.A(n_418),
.B(n_307),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_360),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_395),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g457 ( 
.A1(n_427),
.A2(n_318),
.B(n_307),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_386),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_318),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_401),
.B(n_362),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_409),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_367),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_374),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_384),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_362),
.B(n_352),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_401),
.B(n_352),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_363),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_363),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_359),
.B(n_352),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_411),
.A2(n_307),
.B(n_312),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_374),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_366),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_388),
.B(n_332),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_359),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_366),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_369),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_418),
.B(n_37),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_369),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_323),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_394),
.B(n_349),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_380),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_382),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_375),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_374),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

OR2x2_ASAP7_75t_SL g501 ( 
.A(n_399),
.B(n_336),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_409),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_411),
.A2(n_351),
.B(n_335),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_384),
.B(n_344),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_384),
.B(n_404),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_370),
.B(n_372),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_505),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_SL g516 ( 
.A(n_487),
.B(n_371),
.C(n_365),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_467),
.B(n_370),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_511),
.A2(n_335),
.B1(n_343),
.B2(n_407),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_489),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_456),
.Y(n_521)
);

AOI221x1_ASAP7_75t_L g522 ( 
.A1(n_483),
.A2(n_412),
.B1(n_415),
.B2(n_423),
.C(n_421),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_476),
.B(n_372),
.Y(n_524)
);

OR2x6_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_407),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_511),
.B(n_509),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_450),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_439),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_435),
.A2(n_335),
.B1(n_343),
.B2(n_407),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_474),
.B(n_406),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_407),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_482),
.B(n_406),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_436),
.B(n_410),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_436),
.B(n_364),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_512),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_477),
.B(n_378),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_502),
.B(n_364),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_497),
.B(n_413),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_450),
.A2(n_371),
.B1(n_428),
.B2(n_419),
.Y(n_540)
);

NOR3x1_ASAP7_75t_L g541 ( 
.A(n_433),
.B(n_350),
.C(n_349),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_461),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_489),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_SL g546 ( 
.A(n_502),
.B(n_347),
.C(n_346),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_435),
.A2(n_335),
.B1(n_463),
.B2(n_442),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_444),
.B(n_410),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_438),
.B(n_364),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_444),
.B(n_400),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_434),
.B(n_400),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_458),
.Y(n_552)
);

AND2x6_ASAP7_75t_SL g553 ( 
.A(n_432),
.B(n_0),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_508),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_L g556 ( 
.A(n_469),
.B(n_351),
.C(n_347),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_472),
.B(n_400),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_437),
.B(n_391),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_440),
.B(n_391),
.Y(n_559)
);

AOI221xp5_ASAP7_75t_SL g560 ( 
.A1(n_501),
.A2(n_452),
.B1(n_447),
.B2(n_445),
.C(n_441),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_453),
.B(n_391),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_508),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_472),
.B(n_420),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_464),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_465),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_466),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_484),
.B(n_426),
.Y(n_567)
);

BUFx6f_ASAP7_75t_SL g568 ( 
.A(n_449),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_484),
.B(n_426),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_499),
.B(n_429),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_486),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_499),
.B(n_429),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_SL g574 ( 
.A1(n_507),
.A2(n_431),
.B(n_346),
.C(n_337),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_481),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_468),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_471),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_438),
.A2(n_343),
.B1(n_431),
.B2(n_323),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_520),
.Y(n_579)
);

AND2x2_ASAP7_75t_SL g580 ( 
.A(n_532),
.B(n_492),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_525),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_555),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_527),
.B(n_493),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_525),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_517),
.B(n_454),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_528),
.B(n_493),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_520),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_526),
.B(n_475),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_544),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_526),
.B(n_478),
.Y(n_591)
);

OR2x2_ASAP7_75t_SL g592 ( 
.A(n_516),
.B(n_451),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_SL g593 ( 
.A(n_515),
.B(n_455),
.C(n_451),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_518),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_544),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_524),
.B(n_479),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_551),
.B(n_485),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_555),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_575),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_525),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_556),
.B(n_500),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_551),
.B(n_448),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_SL g603 ( 
.A(n_546),
.B(n_455),
.C(n_446),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_540),
.B(n_449),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_521),
.B(n_449),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_537),
.B(n_552),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_541),
.B(n_504),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_575),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_518),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_536),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_554),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_536),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_530),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_571),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_488),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_543),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_568),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_564),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_565),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_534),
.B(n_533),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_531),
.B(n_576),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_577),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_539),
.B(n_504),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_563),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_573),
.B(n_503),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_548),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_567),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_568),
.A2(n_491),
.B1(n_494),
.B2(n_495),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_569),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_558),
.Y(n_634)
);

BUFx4f_ASAP7_75t_SL g635 ( 
.A(n_538),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_558),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_623),
.A2(n_549),
.B(n_550),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_628),
.A2(n_457),
.B(n_522),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_604),
.A2(n_547),
.B1(n_535),
.B2(n_559),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_584),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_559),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_628),
.A2(n_618),
.B(n_547),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_602),
.A2(n_549),
.B(n_557),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_631),
.B(n_561),
.Y(n_645)
);

CKINVDCx6p67_ASAP7_75t_R g646 ( 
.A(n_611),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_606),
.A2(n_561),
.B1(n_529),
.B2(n_519),
.Y(n_647)
);

OAI21x1_ASAP7_75t_SL g648 ( 
.A1(n_600),
.A2(n_572),
.B(n_570),
.Y(n_648)
);

AOI21x1_ASAP7_75t_SL g649 ( 
.A1(n_597),
.A2(n_574),
.B(n_529),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_631),
.B(n_443),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_628),
.A2(n_578),
.B(n_513),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_625),
.B(n_470),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_580),
.A2(n_574),
.B(n_519),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_588),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_615),
.B(n_506),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_615),
.B(n_337),
.Y(n_656)
);

AOI21xp33_ASAP7_75t_L g657 ( 
.A1(n_604),
.A2(n_583),
.B(n_587),
.Y(n_657)
);

BUFx2_ASAP7_75t_R g658 ( 
.A(n_611),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_580),
.A2(n_578),
.B(n_391),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_607),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_633),
.B(n_514),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_614),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_603),
.B(n_345),
.Y(n_664)
);

AOI21x1_ASAP7_75t_L g665 ( 
.A1(n_596),
.A2(n_510),
.B(n_496),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_589),
.A2(n_343),
.B(n_345),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_633),
.A2(n_448),
.B(n_342),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_591),
.A2(n_448),
.B(n_343),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_624),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_613),
.A2(n_448),
.B(n_343),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_634),
.B(n_448),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_600),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_617),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_622),
.B(n_636),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_613),
.A2(n_448),
.B(n_43),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_617),
.B(n_342),
.Y(n_676)
);

AOI221x1_ASAP7_75t_L g677 ( 
.A1(n_630),
.A2(n_342),
.B1(n_553),
.B2(n_3),
.C(n_4),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_599),
.Y(n_678)
);

CKINVDCx6p67_ASAP7_75t_R g679 ( 
.A(n_620),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_613),
.A2(n_44),
.B(n_38),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_614),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_626),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_581),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_601),
.A2(n_47),
.B(n_46),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_626),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g686 ( 
.A1(n_605),
.A2(n_50),
.B(n_48),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_636),
.B(n_1),
.Y(n_687)
);

OAI21xp33_ASAP7_75t_L g688 ( 
.A1(n_624),
.A2(n_1),
.B(n_2),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_607),
.B(n_51),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_629),
.B(n_53),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_630),
.A2(n_55),
.B(n_54),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_677),
.B(n_632),
.C(n_593),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_637),
.A2(n_601),
.B(n_627),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_661),
.Y(n_694)
);

CKINVDCx11_ASAP7_75t_R g695 ( 
.A(n_646),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_640),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_641),
.A2(n_630),
.B(n_598),
.Y(n_697)
);

AOI31xp67_ASAP7_75t_L g698 ( 
.A1(n_647),
.A2(n_608),
.A3(n_622),
.B(n_607),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_669),
.B(n_581),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_639),
.A2(n_627),
.B(n_582),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_689),
.A2(n_627),
.B1(n_635),
.B2(n_605),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_674),
.B(n_645),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_658),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_621),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_660),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_684),
.A2(n_605),
.B(n_619),
.C(n_616),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_SL g707 ( 
.A(n_644),
.B(n_620),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_663),
.Y(n_708)
);

AO22x2_ASAP7_75t_L g709 ( 
.A1(n_648),
.A2(n_600),
.B1(n_619),
.B2(n_616),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_666),
.A2(n_630),
.B(n_619),
.Y(n_710)
);

AOI211x1_ASAP7_75t_L g711 ( 
.A1(n_657),
.A2(n_579),
.B(n_590),
.C(n_595),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_688),
.A2(n_616),
.B(n_608),
.C(n_594),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_673),
.B(n_620),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_667),
.A2(n_630),
.B(n_605),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_673),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_675),
.A2(n_590),
.B(n_579),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_659),
.A2(n_595),
.B(n_594),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_681),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_687),
.B(n_610),
.Y(n_719)
);

CKINVDCx6p67_ASAP7_75t_R g720 ( 
.A(n_679),
.Y(n_720)
);

OAI21x1_ASAP7_75t_SL g721 ( 
.A1(n_686),
.A2(n_612),
.B(n_610),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_682),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_685),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_660),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_653),
.A2(n_609),
.B(n_594),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_650),
.B(n_687),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_678),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_672),
.B(n_609),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_669),
.B(n_609),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_639),
.A2(n_585),
.B(n_581),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_655),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_683),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_690),
.A2(n_585),
.B1(n_581),
.B2(n_612),
.Y(n_733)
);

AOI21x1_ASAP7_75t_L g734 ( 
.A1(n_665),
.A2(n_592),
.B(n_585),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_678),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_664),
.B(n_592),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_652),
.A2(n_585),
.B(n_581),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_643),
.A2(n_671),
.B(n_691),
.Y(n_738)
);

AO32x2_ASAP7_75t_L g739 ( 
.A1(n_649),
.A2(n_585),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_689),
.B(n_2),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_689),
.B(n_5),
.Y(n_741)
);

CKINVDCx9p33_ASAP7_75t_R g742 ( 
.A(n_662),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_675),
.A2(n_60),
.B(n_59),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_683),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_642),
.Y(n_745)
);

AOI21x1_ASAP7_75t_L g746 ( 
.A1(n_643),
.A2(n_122),
.B(n_180),
.Y(n_746)
);

AND2x6_ASAP7_75t_SL g747 ( 
.A(n_676),
.B(n_6),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_638),
.A2(n_181),
.B(n_121),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_642),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_654),
.B(n_7),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_672),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_638),
.A2(n_651),
.B(n_668),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_668),
.A2(n_123),
.B(n_176),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_661),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_654),
.B(n_8),
.Y(n_755)
);

BUFx8_ASAP7_75t_L g756 ( 
.A(n_715),
.Y(n_756)
);

CKINVDCx11_ASAP7_75t_R g757 ( 
.A(n_695),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_708),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_702),
.B(n_651),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_732),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_692),
.A2(n_680),
.B1(n_661),
.B2(n_670),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_726),
.B(n_680),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_705),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_731),
.B(n_719),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_696),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_701),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_767)
);

BUFx10_ASAP7_75t_L g768 ( 
.A(n_747),
.Y(n_768)
);

INVx6_ASAP7_75t_L g769 ( 
.A(n_732),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_740),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_704),
.B(n_12),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_736),
.A2(n_670),
.B1(n_14),
.B2(n_15),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_732),
.Y(n_773)
);

INVx6_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_694),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_722),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_744),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_741),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_699),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_712),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_720),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_693),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_742),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_751),
.B(n_63),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_730),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_700),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_694),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_SL g788 ( 
.A1(n_709),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_707),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_729),
.B(n_30),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_755),
.B(n_66),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_723),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_737),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_794)
);

CKINVDCx11_ASAP7_75t_R g795 ( 
.A(n_703),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_750),
.B(n_31),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_714),
.A2(n_32),
.B1(n_68),
.B2(n_69),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_735),
.Y(n_798)
);

BUFx4f_ASAP7_75t_SL g799 ( 
.A(n_754),
.Y(n_799)
);

CKINVDCx11_ASAP7_75t_R g800 ( 
.A(n_724),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_SL g801 ( 
.A1(n_709),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_801)
);

BUFx12f_ASAP7_75t_L g802 ( 
.A(n_713),
.Y(n_802)
);

CKINVDCx11_ASAP7_75t_R g803 ( 
.A(n_745),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_749),
.Y(n_804)
);

CKINVDCx11_ASAP7_75t_R g805 ( 
.A(n_739),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_754),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_706),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_749),
.Y(n_808)
);

CKINVDCx11_ASAP7_75t_R g809 ( 
.A(n_739),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_711),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_749),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_738),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_765),
.B(n_697),
.Y(n_813)
);

AOI21xp33_ASAP7_75t_L g814 ( 
.A1(n_807),
.A2(n_733),
.B(n_721),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_806),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_804),
.Y(n_816)
);

INVx5_ASAP7_75t_L g817 ( 
.A(n_774),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_777),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_808),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_811),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_806),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_758),
.B(n_739),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_761),
.B(n_752),
.Y(n_823)
);

AOI21xp33_ASAP7_75t_L g824 ( 
.A1(n_807),
.A2(n_748),
.B(n_743),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_776),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_792),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_775),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_759),
.Y(n_828)
);

AO21x1_ASAP7_75t_SL g829 ( 
.A1(n_763),
.A2(n_698),
.B(n_734),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_805),
.B(n_716),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_759),
.B(n_746),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_764),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_793),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_756),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_798),
.Y(n_835)
);

AOI21xp33_ASAP7_75t_L g836 ( 
.A1(n_780),
.A2(n_753),
.B(n_725),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_809),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_775),
.B(n_710),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_810),
.Y(n_839)
);

OA21x2_ASAP7_75t_L g840 ( 
.A1(n_810),
.A2(n_717),
.B(n_728),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_788),
.B(n_728),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_774),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_790),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_780),
.A2(n_711),
.B(n_89),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_789),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_762),
.B(n_95),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_756),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_760),
.B(n_96),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_757),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_760),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_796),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_773),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_787),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_799),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_795),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_773),
.B(n_97),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_815),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_813),
.B(n_783),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_825),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_817),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_826),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_828),
.B(n_771),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_851),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_826),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_819),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_823),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_822),
.B(n_800),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_SL g868 ( 
.A1(n_840),
.A2(n_784),
.B(n_839),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_823),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_819),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_828),
.B(n_766),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_817),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_816),
.B(n_767),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_820),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_836),
.A2(n_767),
.B(n_770),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_824),
.A2(n_791),
.B(n_784),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_850),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_820),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_816),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_815),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_822),
.B(n_803),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_833),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_833),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_835),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_835),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_874),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_866),
.B(n_830),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_860),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_874),
.Y(n_889)
);

AO21x2_ASAP7_75t_L g890 ( 
.A1(n_868),
.A2(n_844),
.B(n_831),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_880),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_865),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_866),
.B(n_831),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_869),
.B(n_830),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_859),
.B(n_843),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_868),
.B(n_839),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_865),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_858),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_869),
.B(n_831),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_879),
.A2(n_844),
.B(n_831),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_870),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_877),
.B(n_843),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_867),
.B(n_837),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_870),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_862),
.B(n_851),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_860),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_860),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_903),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_888),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_902),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_886),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_896),
.A2(n_837),
.B1(n_873),
.B2(n_786),
.Y(n_912)
);

NOR2x1_ASAP7_75t_SL g913 ( 
.A(n_896),
.B(n_860),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_892),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_907),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_893),
.B(n_871),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_892),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_897),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_902),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_897),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_901),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_886),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_905),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_889),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_L g925 ( 
.A(n_907),
.B(n_849),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_889),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_917),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_909),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_908),
.B(n_903),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_909),
.B(n_887),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_923),
.B(n_887),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_915),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_915),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_913),
.B(n_894),
.Y(n_934)
);

AOI21xp33_ASAP7_75t_L g935 ( 
.A1(n_912),
.A2(n_875),
.B(n_890),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_913),
.B(n_894),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_915),
.B(n_906),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_916),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_927),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_938),
.B(n_910),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_937),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_927),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_929),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_930),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_928),
.B(n_916),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_931),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_946),
.B(n_932),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_942),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_941),
.A2(n_935),
.B1(n_936),
.B2(n_934),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_944),
.B(n_925),
.Y(n_950)
);

OAI221xp5_ASAP7_75t_L g951 ( 
.A1(n_943),
.A2(n_935),
.B1(n_933),
.B2(n_896),
.C(n_906),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_939),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_940),
.B(n_945),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_949),
.A2(n_768),
.B1(n_875),
.B2(n_890),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_948),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_951),
.A2(n_940),
.B1(n_942),
.B2(n_896),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_950),
.B(n_849),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_947),
.B(n_834),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_948),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_948),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_952),
.B(n_919),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_950),
.B(n_834),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_955),
.Y(n_963)
);

AO22x2_ASAP7_75t_L g964 ( 
.A1(n_959),
.A2(n_853),
.B1(n_847),
.B2(n_854),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_960),
.B(n_867),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_961),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_953),
.A2(n_890),
.B1(n_896),
.B2(n_907),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_957),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_958),
.B(n_881),
.Y(n_969)
);

AOI21xp33_ASAP7_75t_L g970 ( 
.A1(n_956),
.A2(n_875),
.B(n_853),
.Y(n_970)
);

AOI21xp33_ASAP7_75t_L g971 ( 
.A1(n_968),
.A2(n_962),
.B(n_954),
.Y(n_971)
);

NOR4xp25_ASAP7_75t_SL g972 ( 
.A(n_963),
.B(n_954),
.C(n_854),
.D(n_855),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_964),
.B(n_966),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_969),
.B(n_847),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_965),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_967),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_863),
.B1(n_845),
.B2(n_778),
.C(n_881),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_963),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_972),
.A2(n_898),
.B1(n_818),
.B2(n_888),
.Y(n_979)
);

AOI221xp5_ASAP7_75t_SL g980 ( 
.A1(n_973),
.A2(n_768),
.B1(n_782),
.B2(n_846),
.C(n_785),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_976),
.A2(n_975),
.B1(n_977),
.B2(n_971),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_SL g982 ( 
.A1(n_978),
.A2(n_781),
.B(n_856),
.Y(n_982)
);

AOI322xp5_ASAP7_75t_L g983 ( 
.A1(n_974),
.A2(n_779),
.A3(n_846),
.B1(n_841),
.B2(n_794),
.C1(n_888),
.C2(n_879),
.Y(n_983)
);

AOI222xp33_ASAP7_75t_L g984 ( 
.A1(n_973),
.A2(n_841),
.B1(n_797),
.B2(n_907),
.C1(n_772),
.C2(n_812),
.Y(n_984)
);

AOI322xp5_ASAP7_75t_L g985 ( 
.A1(n_973),
.A2(n_917),
.A3(n_921),
.B1(n_920),
.B2(n_895),
.C1(n_801),
.C2(n_918),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_982),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_981),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_979),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_984),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_980),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_983),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_985),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_982),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_981),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_981),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_L g996 ( 
.A(n_988),
.B(n_856),
.C(n_848),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_986),
.A2(n_926),
.B(n_924),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_987),
.Y(n_998)
);

NOR4xp25_ASAP7_75t_L g999 ( 
.A(n_994),
.B(n_920),
.C(n_921),
.D(n_914),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_986),
.B(n_860),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_995),
.A2(n_871),
.B1(n_924),
.B2(n_922),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_990),
.B(n_856),
.C(n_848),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_992),
.A2(n_991),
.B1(n_989),
.B2(n_993),
.Y(n_1003)
);

NOR2x1p5_ASAP7_75t_L g1004 ( 
.A(n_986),
.B(n_802),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_988),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_1005),
.B(n_911),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_1000),
.Y(n_1007)
);

OAI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_817),
.B(n_862),
.C(n_842),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_996),
.A2(n_891),
.B(n_922),
.C(n_911),
.Y(n_1009)
);

NOR5xp2_ASAP7_75t_L g1010 ( 
.A(n_1004),
.B(n_999),
.C(n_997),
.D(n_1002),
.E(n_1001),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1000),
.A2(n_926),
.B(n_856),
.Y(n_1011)
);

AOI211x1_ASAP7_75t_SL g1012 ( 
.A1(n_1000),
.A2(n_842),
.B(n_852),
.C(n_814),
.Y(n_1012)
);

AOI221xp5_ASAP7_75t_L g1013 ( 
.A1(n_1007),
.A2(n_848),
.B1(n_891),
.B2(n_900),
.C(n_773),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_L g1014 ( 
.A(n_1008),
.B(n_848),
.C(n_827),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1006),
.B(n_900),
.Y(n_1015)
);

OAI221xp5_ASAP7_75t_SL g1016 ( 
.A1(n_1009),
.A2(n_873),
.B1(n_872),
.B2(n_893),
.C(n_899),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_1011),
.B(n_769),
.Y(n_1017)
);

OAI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_1012),
.A2(n_872),
.B1(n_827),
.B2(n_817),
.C(n_769),
.Y(n_1018)
);

NOR5xp2_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_904),
.C(n_901),
.D(n_878),
.E(n_861),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1007),
.B(n_900),
.Y(n_1020)
);

OAI221xp5_ASAP7_75t_L g1021 ( 
.A1(n_1007),
.A2(n_827),
.B1(n_817),
.B2(n_838),
.C(n_899),
.Y(n_1021)
);

NOR4xp25_ASAP7_75t_L g1022 ( 
.A(n_1007),
.B(n_904),
.C(n_852),
.D(n_857),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_817),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_1020),
.B(n_876),
.Y(n_1024)
);

NAND4xp75_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_884),
.C(n_883),
.D(n_882),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_1016),
.B(n_857),
.C(n_821),
.Y(n_1026)
);

NAND4xp25_ASAP7_75t_SL g1027 ( 
.A(n_1014),
.B(n_1013),
.C(n_1021),
.D(n_1019),
.Y(n_1027)
);

OAI211xp5_ASAP7_75t_SL g1028 ( 
.A1(n_1018),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_1028)
);

NAND4xp25_ASAP7_75t_L g1029 ( 
.A(n_1022),
.B(n_815),
.C(n_821),
.D(n_857),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_SL g1030 ( 
.A1(n_1017),
.A2(n_880),
.B1(n_838),
.B2(n_840),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1015),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_1020),
.A2(n_876),
.B(n_838),
.C(n_882),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1023),
.B(n_876),
.Y(n_1033)
);

NOR4xp75_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_821),
.C(n_102),
.D(n_106),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_101),
.C(n_108),
.Y(n_1035)
);

NAND4xp75_ASAP7_75t_L g1036 ( 
.A(n_1024),
.B(n_111),
.C(n_112),
.D(n_113),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_883),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_1027),
.B(n_116),
.Y(n_1038)
);

AOI31xp33_ASAP7_75t_L g1039 ( 
.A1(n_1028),
.A2(n_884),
.A3(n_864),
.B(n_861),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1026),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_1030),
.B(n_117),
.C(n_120),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_1027),
.B(n_124),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_SL g1044 ( 
.A(n_1023),
.B(n_126),
.C(n_127),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1031),
.Y(n_1045)
);

AO22x1_ASAP7_75t_L g1046 ( 
.A1(n_1043),
.A2(n_864),
.B1(n_878),
.B2(n_885),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1036),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1038),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1045),
.B(n_885),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1040),
.A2(n_1035),
.B1(n_1042),
.B2(n_1044),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1041),
.A2(n_832),
.B1(n_840),
.B2(n_134),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_1037),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1039),
.B(n_832),
.Y(n_1053)
);

XOR2xp5_ASAP7_75t_L g1054 ( 
.A(n_1033),
.B(n_129),
.Y(n_1054)
);

AO22x1_ASAP7_75t_L g1055 ( 
.A1(n_1048),
.A2(n_1034),
.B1(n_135),
.B2(n_136),
.Y(n_1055)
);

AO22x2_ASAP7_75t_L g1056 ( 
.A1(n_1054),
.A2(n_133),
.B1(n_138),
.B2(n_141),
.Y(n_1056)
);

AO22x2_ASAP7_75t_L g1057 ( 
.A1(n_1047),
.A2(n_1049),
.B1(n_1053),
.B2(n_1052),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1050),
.A2(n_840),
.B1(n_143),
.B2(n_144),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1051),
.A2(n_829),
.B1(n_146),
.B2(n_147),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1046),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

XOR2xp5_ASAP7_75t_L g1062 ( 
.A(n_1057),
.B(n_142),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_1056),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1055),
.B(n_148),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_1062),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_1065),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1066),
.A2(n_1061),
.B1(n_1063),
.B2(n_1060),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_1067),
.A2(n_1064),
.B1(n_1058),
.B2(n_1059),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1068),
.B(n_150),
.Y(n_1069)
);

AOI311xp33_ASAP7_75t_L g1070 ( 
.A1(n_1069),
.A2(n_151),
.A3(n_153),
.B(n_156),
.C(n_157),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1070),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_1071)
);

AOI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_1071),
.A2(n_165),
.B(n_166),
.C(n_167),
.Y(n_1072)
);


endmodule