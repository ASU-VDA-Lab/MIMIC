module fake_jpeg_24667_n_137 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_11),
.Y(n_37)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_29),
.B1(n_30),
.B2(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_21),
.B1(n_12),
.B2(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_21),
.B1(n_19),
.B2(n_11),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_21),
.B1(n_13),
.B2(n_19),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_18),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_50),
.B1(n_51),
.B2(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_31),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_38),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_32),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_40),
.B(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_59),
.B1(n_11),
.B2(n_20),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_42),
.B(n_49),
.C(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_64),
.B1(n_19),
.B2(n_13),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_33),
.B1(n_34),
.B2(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_62),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_58),
.B(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_61),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_16),
.B1(n_14),
.B2(n_18),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_77),
.B(n_56),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_28),
.B1(n_27),
.B2(n_45),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_32),
.B1(n_19),
.B2(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_46),
.B1(n_60),
.B2(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_57),
.C(n_66),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_75),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_59),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_81),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_74),
.B(n_77),
.C(n_15),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_82),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_14),
.B(n_16),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_52),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_87),
.C(n_85),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.C(n_108),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_9),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_15),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_110),
.C(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_93),
.C(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_2),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_96),
.B1(n_98),
.B2(n_32),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_52),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_105),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_111),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_3),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_3),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_121),
.B(n_120),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_6),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_3),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_125),
.B(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_5),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_5),
.C(n_6),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);


endmodule