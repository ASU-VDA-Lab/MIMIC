module fake_jpeg_10701_n_400 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_400);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_400;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_74),
.Y(n_125)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_7),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_65),
.B(n_91),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_72),
.Y(n_132)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_17),
.B(n_5),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_77),
.B(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_25),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_88),
.Y(n_145)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_85),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_95),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_41),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_6),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_111),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_108),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_49),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_27),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_27),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_110),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_32),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_32),
.B(n_10),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_51),
.B(n_50),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_99),
.Y(n_182)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_39),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_122),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_124),
.B(n_126),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_39),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_24),
.B1(n_31),
.B2(n_29),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_127),
.A2(n_139),
.B1(n_150),
.B2(n_156),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_59),
.A2(n_31),
.B1(n_50),
.B2(n_42),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_80),
.A2(n_40),
.B(n_47),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_161),
.C(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_40),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_143),
.B(n_176),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_41),
.B1(n_47),
.B2(n_45),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_149),
.B1(n_154),
.B2(n_158),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g147 ( 
.A(n_92),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_147),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_97),
.A2(n_37),
.B1(n_51),
.B2(n_42),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_71),
.A2(n_37),
.B1(n_53),
.B2(n_36),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_98),
.A2(n_36),
.B(n_45),
.C(n_53),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_93),
.B1(n_57),
.B2(n_104),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_11),
.B1(n_16),
.B2(n_1),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_11),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_94),
.A2(n_11),
.B1(n_16),
.B2(n_3),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_3),
.B1(n_16),
.B2(n_106),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_153),
.B1(n_131),
.B2(n_141),
.Y(n_205)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_78),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_182),
.B(n_188),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_3),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_186),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_101),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_93),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_189),
.B(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_73),
.B1(n_86),
.B2(n_104),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_190),
.A2(n_200),
.B1(n_203),
.B2(n_205),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_201),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_131),
.A2(n_112),
.B1(n_119),
.B2(n_159),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_169),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_232),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

INVx2_ASAP7_75t_R g198 ( 
.A(n_115),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_202),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_137),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_139),
.A2(n_112),
.B1(n_149),
.B2(n_162),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

NAND2x1_ASAP7_75t_SL g202 ( 
.A(n_136),
.B(n_141),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_156),
.A2(n_127),
.B1(n_134),
.B2(n_116),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_145),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_214),
.C(n_182),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_138),
.A2(n_117),
.B1(n_170),
.B2(n_129),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_224),
.B1(n_236),
.B2(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_217),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_168),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

OR2x2_ASAP7_75t_SL g217 ( 
.A(n_171),
.B(n_120),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_160),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_220),
.B(n_230),
.Y(n_273)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_222),
.B(n_226),
.Y(n_267)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_128),
.A2(n_165),
.B1(n_129),
.B2(n_170),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_123),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_130),
.A2(n_155),
.B1(n_167),
.B2(n_165),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_227),
.A2(n_231),
.B1(n_228),
.B2(n_232),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_130),
.B(n_155),
.CI(n_167),
.CON(n_228),
.SN(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_233),
.Y(n_253)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_123),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_175),
.A2(n_150),
.B1(n_139),
.B2(n_125),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_175),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_125),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_235),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_132),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_124),
.A2(n_158),
.B1(n_139),
.B2(n_57),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_124),
.B(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_195),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_241),
.A2(n_194),
.B1(n_225),
.B2(n_210),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_186),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_182),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_262),
.Y(n_289)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_183),
.B(n_228),
.C(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_207),
.C(n_181),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_185),
.C(n_206),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_204),
.C(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_191),
.B(n_187),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_191),
.B(n_214),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_203),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_213),
.A2(n_188),
.B1(n_223),
.B2(n_224),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_268),
.B1(n_251),
.B2(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_197),
.B(n_209),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_266),
.B(n_271),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_201),
.B(n_215),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_216),
.Y(n_275)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_277),
.Y(n_331)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_219),
.B(n_202),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_296),
.B(n_293),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_185),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_303),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_300),
.B(n_308),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_284),
.A2(n_259),
.B1(n_270),
.B2(n_257),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_229),
.B1(n_196),
.B2(n_221),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_241),
.B1(n_304),
.B2(n_286),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_292),
.Y(n_310)
);

XOR2x2_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_206),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_291),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_240),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_294),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_240),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_238),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_306),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_301),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_264),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_307),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_253),
.A2(n_238),
.B(n_248),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_239),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_304),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_252),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_242),
.B(n_246),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_242),
.B(n_249),
.C(n_263),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_261),
.B(n_265),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_313),
.A2(n_322),
.B1(n_294),
.B2(n_288),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_289),
.A2(n_257),
.B1(n_276),
.B2(n_271),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_320),
.B1(n_290),
.B2(n_305),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_321),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_276),
.B(n_274),
.C(n_259),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_318),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_282),
.A2(n_299),
.B1(n_308),
.B2(n_306),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_299),
.A2(n_287),
.B1(n_278),
.B2(n_298),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_307),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_279),
.Y(n_340)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_303),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_338),
.C(n_339),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_335),
.B(n_345),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_279),
.B1(n_300),
.B2(n_290),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_337),
.B1(n_342),
.B2(n_330),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_283),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_283),
.Y(n_339)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_326),
.A2(n_321),
.B(n_283),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_341),
.A2(n_311),
.B(n_327),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_302),
.B1(n_295),
.B2(n_285),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_298),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_347),
.C(n_330),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_295),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_344),
.B(n_348),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_327),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_280),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_324),
.B(n_291),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_310),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_310),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_335),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_320),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_353),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_317),
.B1(n_328),
.B2(n_315),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_356),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_346),
.A2(n_317),
.B1(n_329),
.B2(n_318),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_359),
.B(n_324),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_329),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_334),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_361),
.A2(n_311),
.B(n_331),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_332),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_314),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_351),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_361),
.B(n_346),
.C(n_356),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_370),
.Y(n_380)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

XOR2x2_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_369),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_363),
.A2(n_336),
.B(n_341),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_373),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_343),
.C(n_347),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_352),
.C(n_350),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_376),
.B(n_377),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_360),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_378),
.B(n_364),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_367),
.A2(n_355),
.B1(n_354),
.B2(n_313),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_382),
.A2(n_372),
.B(n_371),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_369),
.B(n_366),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_384),
.A2(n_379),
.B(n_368),
.Y(n_392)
);

AOI21x1_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_353),
.B(n_374),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_376),
.C(n_378),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_386),
.B(n_388),
.Y(n_391)
);

AOI31xp67_ASAP7_75t_SL g388 ( 
.A1(n_375),
.A2(n_316),
.A3(n_331),
.B(n_358),
.Y(n_388)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_387),
.A2(n_377),
.B(n_379),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_389),
.A2(n_390),
.B(n_392),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_365),
.B(n_319),
.C(n_316),
.Y(n_394)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_323),
.B1(n_256),
.B2(n_260),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_323),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_396),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_399),
.B(n_398),
.Y(n_400)
);


endmodule