module fake_jpeg_10654_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_30),
.Y(n_67)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_49),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_24),
.B(n_33),
.C(n_17),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_56),
.B(n_70),
.C(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_59),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_26),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_34),
.B1(n_26),
.B2(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_26),
.Y(n_70)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_70),
.B1(n_51),
.B2(n_44),
.Y(n_72)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_44),
.B1(n_58),
.B2(n_35),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_80),
.B1(n_89),
.B2(n_94),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_34),
.B(n_19),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_42),
.B1(n_41),
.B2(n_31),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_86),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_45),
.B1(n_35),
.B2(n_38),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_57),
.B1(n_49),
.B2(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_31),
.B1(n_45),
.B2(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_50),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_47),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_52),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_122),
.B1(n_78),
.B2(n_71),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_56),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_109),
.B(n_72),
.Y(n_147)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_45),
.B1(n_38),
.B2(n_54),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_45),
.B1(n_38),
.B2(n_63),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_22),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_124),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_68),
.B1(n_46),
.B2(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_50),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_145),
.B1(n_104),
.B2(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_124),
.B1(n_108),
.B2(n_115),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_72),
.B(n_89),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_101),
.B(n_99),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_73),
.B1(n_78),
.B2(n_63),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_153),
.B1(n_104),
.B2(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_112),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_109),
.B1(n_108),
.B2(n_113),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_157),
.B(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_180),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_107),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_170),
.B1(n_135),
.B2(n_133),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_103),
.A3(n_116),
.B1(n_107),
.B2(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_165),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_107),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_28),
.B(n_20),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_176),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_111),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_169),
.C(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_98),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_86),
.B1(n_75),
.B2(n_81),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_81),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_33),
.B(n_22),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_139),
.B(n_28),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_106),
.C(n_86),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_106),
.C(n_50),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_19),
.C(n_25),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_23),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_181),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_23),
.B(n_18),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_152),
.B(n_136),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_138),
.B(n_137),
.C(n_141),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_23),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_33),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_191),
.B1(n_176),
.B2(n_165),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_186),
.B(n_194),
.Y(n_234)
);

OR2x6_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_153),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_181),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_126),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_193),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_145),
.B1(n_127),
.B2(n_28),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_162),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_127),
.B(n_87),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_19),
.B(n_25),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_206),
.B1(n_32),
.B2(n_20),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_198),
.B(n_202),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_32),
.B(n_18),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_44),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_174),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_169),
.Y(n_225)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_219),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_157),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_164),
.B1(n_155),
.B2(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_163),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_225),
.C(n_229),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_170),
.B1(n_172),
.B2(n_158),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_231),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_232),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_171),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_19),
.C(n_10),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_29),
.B1(n_8),
.B2(n_10),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_17),
.C(n_22),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_9),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_189),
.C(n_207),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_186),
.B1(n_199),
.B2(n_203),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_243),
.B1(n_245),
.B2(n_251),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_186),
.B1(n_201),
.B2(n_192),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_187),
.B1(n_183),
.B2(n_198),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_17),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_0),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_212),
.B(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_29),
.C(n_1),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_0),
.C(n_1),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_212),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_211),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_244),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_269),
.B(n_271),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_248),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_251),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_210),
.B(n_222),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_241),
.C(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_SL g275 ( 
.A(n_269),
.B(n_253),
.C(n_256),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_268),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_237),
.B(n_245),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_283),
.B(n_5),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_0),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_235),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_288),
.C(n_5),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_254),
.B1(n_253),
.B2(n_242),
.Y(n_281)
);

AOI22x1_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_262),
.B1(n_258),
.B2(n_260),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_249),
.B(n_225),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_7),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_6),
.C(n_15),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_291),
.B(n_293),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_292),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_281),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_272),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_279),
.B(n_275),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_296),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_11),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.C(n_300),
.Y(n_304)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_279),
.B1(n_277),
.B2(n_2),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_305),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_311),
.Y(n_312)
);

NAND4xp25_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_299),
.C(n_301),
.D(n_290),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_300),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_4),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_317),
.B(n_318),
.Y(n_321)
);

AOI21x1_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_3),
.B(n_12),
.Y(n_316)
);

AO21x2_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_16),
.B(n_1),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_3),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_13),
.C(n_16),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_13),
.C(n_16),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_0),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_303),
.C(n_310),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_322),
.C(n_323),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_305),
.B(n_13),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_312),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_312),
.B(n_321),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_2),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_2),
.Y(n_329)
);


endmodule