module real_aes_17250_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_269;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1280;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g687 ( .A(n_0), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_0), .A2(n_214), .B1(n_1296), .B2(n_1311), .Y(n_1323) );
INVx1_ASAP7_75t_L g554 ( .A(n_1), .Y(n_554) );
AOI221x1_ASAP7_75t_SL g585 ( .A1(n_1), .A2(n_2), .B1(n_586), .B2(n_588), .C(n_590), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_2), .A2(n_23), .B1(n_560), .B2(n_562), .Y(n_570) );
INVx1_ASAP7_75t_L g1525 ( .A(n_3), .Y(n_1525) );
OAI211xp5_ASAP7_75t_L g1221 ( .A1(n_4), .A2(n_418), .B(n_1217), .C(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1238 ( .A(n_4), .Y(n_1238) );
AOI221x1_ASAP7_75t_SL g700 ( .A1(n_5), .A2(n_255), .B1(n_701), .B2(n_705), .C(n_707), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g774 ( .A1(n_5), .A2(n_599), .B(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_6), .A2(n_54), .B1(n_1296), .B2(n_1311), .Y(n_1319) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_7), .Y(n_924) );
INVx1_ASAP7_75t_L g616 ( .A(n_8), .Y(n_616) );
OAI211xp5_ASAP7_75t_L g671 ( .A1(n_8), .A2(n_645), .B(n_672), .C(n_673), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_9), .A2(n_218), .B1(n_1042), .B2(n_1043), .C(n_1046), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_9), .A2(n_218), .B1(n_522), .B2(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g319 ( .A(n_10), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_11), .A2(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g602 ( .A(n_11), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_12), .A2(n_252), .B1(n_967), .B2(n_1031), .C(n_1032), .Y(n_1030) );
AOI222xp33_ASAP7_75t_L g1069 ( .A1(n_12), .A2(n_64), .B1(n_147), .B2(n_342), .C1(n_361), .C2(n_921), .Y(n_1069) );
INVx1_ASAP7_75t_L g1039 ( .A(n_13), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_13), .A2(n_257), .B1(n_496), .B2(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g283 ( .A(n_14), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_14), .B(n_293), .Y(n_369) );
AND2x2_ASAP7_75t_L g493 ( .A(n_14), .B(n_447), .Y(n_493) );
AND2x2_ASAP7_75t_L g552 ( .A(n_14), .B(n_232), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_15), .A2(n_111), .B1(n_706), .B2(n_1032), .C(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1158 ( .A(n_15), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_16), .A2(n_187), .B1(n_798), .B2(n_918), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_16), .A2(n_88), .B1(n_543), .B2(n_819), .C(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g1253 ( .A(n_17), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g1283 ( .A1(n_17), .A2(n_125), .B1(n_1059), .B2(n_1284), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1256 ( .A1(n_18), .A2(n_256), .B1(n_1042), .B2(n_1043), .C(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1280 ( .A(n_18), .Y(n_1280) );
INVx1_ASAP7_75t_L g359 ( .A(n_19), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_20), .A2(n_265), .B1(n_1057), .B2(n_1527), .Y(n_1526) );
OAI211xp5_ASAP7_75t_L g1529 ( .A1(n_20), .A2(n_1027), .B(n_1530), .C(n_1534), .Y(n_1529) );
INVx1_ASAP7_75t_L g911 ( .A(n_21), .Y(n_911) );
INVx2_ASAP7_75t_L g1299 ( .A(n_22), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_22), .B(n_103), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_22), .B(n_1305), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_23), .A2(n_185), .B1(n_588), .B2(n_597), .C(n_600), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g1336 ( .A1(n_24), .A2(n_35), .B1(n_1303), .B2(n_1306), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_25), .A2(n_144), .B1(n_730), .B2(n_733), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_25), .A2(n_236), .B1(n_740), .B2(n_742), .C(n_744), .Y(n_739) );
INVx1_ASAP7_75t_L g1522 ( .A(n_26), .Y(n_1522) );
OAI221xp5_ASAP7_75t_L g1539 ( .A1(n_26), .A2(n_164), .B1(n_1540), .B2(n_1541), .C(n_1542), .Y(n_1539) );
AOI22xp5_ASAP7_75t_L g1322 ( .A1(n_27), .A2(n_123), .B1(n_1303), .B2(n_1306), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_28), .A2(n_201), .B1(n_796), .B2(n_918), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_28), .A2(n_128), .B1(n_990), .B2(n_1005), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_29), .A2(n_212), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI221xp5_ASAP7_75t_L g929 ( .A1(n_29), .A2(n_60), .B1(n_542), .B2(n_930), .C(n_932), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_30), .A2(n_128), .B1(n_796), .B2(n_918), .Y(n_1107) );
AOI22xp33_ASAP7_75t_SL g1118 ( .A1(n_30), .A2(n_201), .B1(n_1000), .B2(n_1119), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_31), .A2(n_70), .B1(n_562), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1162 ( .A(n_31), .Y(n_1162) );
OAI22xp33_ASAP7_75t_L g1219 ( .A1(n_32), .A2(n_189), .B1(n_410), .B2(n_1220), .Y(n_1219) );
OAI22xp33_ASAP7_75t_L g1230 ( .A1(n_32), .A2(n_189), .B1(n_285), .B2(n_1231), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_33), .A2(n_118), .B1(n_619), .B2(n_972), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_33), .A2(n_266), .B1(n_976), .B2(n_977), .Y(n_975) );
INVx1_ASAP7_75t_L g639 ( .A(n_34), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_36), .A2(n_101), .B1(n_796), .B2(n_891), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_36), .A2(n_245), .B1(n_542), .B2(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g845 ( .A(n_37), .Y(n_845) );
INVx1_ASAP7_75t_L g968 ( .A(n_38), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_39), .A2(n_96), .B1(n_1296), .B2(n_1300), .Y(n_1295) );
INVx1_ASAP7_75t_L g615 ( .A(n_40), .Y(n_615) );
INVx1_ASAP7_75t_L g1197 ( .A(n_41), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_42), .A2(n_229), .B1(n_819), .B2(n_1034), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_42), .A2(n_111), .B1(n_881), .B2(n_1164), .Y(n_1163) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_43), .A2(n_91), .B1(n_1296), .B2(n_1332), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_44), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_45), .A2(n_72), .B1(n_757), .B2(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g837 ( .A(n_45), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_46), .A2(n_166), .B1(n_618), .B2(n_619), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_46), .A2(n_166), .B1(n_668), .B2(n_670), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_47), .A2(n_140), .B1(n_967), .B2(n_1032), .C(n_1250), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_47), .A2(n_74), .B1(n_802), .B2(n_908), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_48), .A2(n_177), .B1(n_574), .B2(n_723), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_48), .A2(n_102), .B1(n_586), .B2(n_800), .Y(n_1277) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_49), .A2(n_186), .B1(n_535), .B2(n_537), .Y(n_534) );
INVx1_ASAP7_75t_L g541 ( .A(n_49), .Y(n_541) );
INVx1_ASAP7_75t_L g427 ( .A(n_50), .Y(n_427) );
INVx1_ASAP7_75t_L g318 ( .A(n_51), .Y(n_318) );
INVx1_ASAP7_75t_L g324 ( .A(n_51), .Y(n_324) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_52), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_52), .A2(n_252), .B1(n_748), .B2(n_794), .Y(n_1074) );
INVx1_ASAP7_75t_L g1187 ( .A(n_53), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g1345 ( .A1(n_55), .A2(n_138), .B1(n_1296), .B2(n_1332), .Y(n_1345) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_56), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_57), .A2(n_230), .B1(n_1303), .B2(n_1306), .Y(n_1302) );
INVx1_ASAP7_75t_L g966 ( .A(n_58), .Y(n_966) );
INVx1_ASAP7_75t_L g1146 ( .A(n_59), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_60), .A2(n_191), .B1(n_794), .B2(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g276 ( .A(n_61), .Y(n_276) );
INVx2_ASAP7_75t_L g310 ( .A(n_62), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_63), .A2(n_216), .B1(n_990), .B2(n_991), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_63), .A2(n_87), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_64), .A2(n_160), .B1(n_1005), .B2(n_1034), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_65), .A2(n_227), .B1(n_512), .B2(n_1128), .Y(n_1269) );
INVx1_ASAP7_75t_L g1268 ( .A(n_66), .Y(n_1268) );
INVx1_ASAP7_75t_L g312 ( .A(n_67), .Y(n_312) );
XNOR2xp5_ASAP7_75t_L g1557 ( .A(n_68), .B(n_1558), .Y(n_1557) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_69), .A2(n_107), .B1(n_556), .B2(n_706), .C(n_864), .Y(n_1140) );
INVxp67_ASAP7_75t_SL g1150 ( .A(n_69), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g1152 ( .A(n_70), .Y(n_1152) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_71), .A2(n_387), .B(n_472), .C(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g677 ( .A(n_71), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_72), .A2(n_127), .B1(n_817), .B2(n_819), .C(n_820), .Y(n_816) );
INVx1_ASAP7_75t_L g327 ( .A(n_73), .Y(n_327) );
INVxp67_ASAP7_75t_SL g1260 ( .A(n_74), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_75), .A2(n_85), .B1(n_408), .B2(n_411), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g443 ( .A1(n_75), .A2(n_116), .B1(n_285), .B2(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_76), .A2(n_180), .B1(n_709), .B2(n_711), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_76), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g915 ( .A(n_77), .Y(n_915) );
INVx1_ASAP7_75t_L g1076 ( .A(n_78), .Y(n_1076) );
INVx1_ASAP7_75t_L g1224 ( .A(n_79), .Y(n_1224) );
OAI211xp5_ASAP7_75t_L g1232 ( .A1(n_79), .A2(n_545), .B(n_1233), .C(n_1235), .Y(n_1232) );
AOI22xp5_ASAP7_75t_L g1312 ( .A1(n_80), .A2(n_124), .B1(n_1303), .B2(n_1306), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_81), .A2(n_108), .B1(n_1296), .B2(n_1311), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_82), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g1520 ( .A1(n_83), .A2(n_243), .B1(n_777), .B2(n_886), .Y(n_1520) );
AOI221xp5_ASAP7_75t_L g1535 ( .A1(n_83), .A2(n_129), .B1(n_967), .B2(n_1032), .C(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g565 ( .A(n_84), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_85), .A2(n_182), .B1(n_451), .B2(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g1199 ( .A(n_86), .Y(n_1199) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_87), .A2(n_208), .B1(n_990), .B2(n_1005), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_88), .A2(n_130), .B1(n_586), .B2(n_800), .Y(n_906) );
INVx1_ASAP7_75t_L g1092 ( .A(n_89), .Y(n_1092) );
INVx1_ASAP7_75t_L g1200 ( .A(n_90), .Y(n_1200) );
OA222x2_ASAP7_75t_L g689 ( .A1(n_92), .A2(n_213), .B1(n_236), .B2(n_690), .C1(n_694), .C2(n_698), .Y(n_689) );
INVx1_ASAP7_75t_L g755 ( .A(n_92), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_93), .A2(n_610), .B1(n_611), .B2(n_680), .Y(n_609) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_93), .Y(n_680) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_94), .Y(n_278) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_94), .B(n_276), .Y(n_1297) );
OAI211xp5_ASAP7_75t_SL g1026 ( .A1(n_95), .A2(n_1027), .B(n_1029), .C(n_1036), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_95), .A2(n_219), .B1(n_512), .B2(n_1057), .Y(n_1056) );
XNOR2xp5_ASAP7_75t_L g1024 ( .A(n_96), .B(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1095 ( .A(n_97), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_97), .A2(n_253), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
INVx1_ASAP7_75t_L g1174 ( .A(n_98), .Y(n_1174) );
INVx1_ASAP7_75t_L g363 ( .A(n_99), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_100), .Y(n_807) );
INVxp67_ASAP7_75t_SL g1543 ( .A(n_101), .Y(n_1543) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_102), .A2(n_162), .B1(n_703), .B2(n_1262), .C(n_1264), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_103), .B(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1305 ( .A(n_103), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_104), .A2(n_199), .B1(n_543), .B2(n_860), .Y(n_859) );
INVxp67_ASAP7_75t_SL g879 ( .A(n_104), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_105), .A2(n_137), .B1(n_987), .B2(n_988), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_105), .A2(n_172), .B1(n_1008), .B2(n_1010), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_106), .A2(n_115), .B1(n_588), .B2(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g839 ( .A(n_106), .Y(n_839) );
INVx1_ASAP7_75t_L g1160 ( .A(n_107), .Y(n_1160) );
INVx1_ASAP7_75t_L g1096 ( .A(n_109), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g1049 ( .A(n_110), .Y(n_1049) );
INVx1_ASAP7_75t_L g789 ( .A(n_112), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_112), .A2(n_241), .B1(n_378), .B2(n_710), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g1344 ( .A1(n_113), .A2(n_174), .B1(n_1303), .B2(n_1306), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_114), .A2(n_245), .B1(n_796), .B2(n_1518), .Y(n_1517) );
AOI21xp33_ASAP7_75t_L g1545 ( .A1(n_114), .A2(n_1031), .B(n_1264), .Y(n_1545) );
INVx1_ASAP7_75t_L g822 ( .A(n_115), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_116), .A2(n_182), .B1(n_432), .B2(n_435), .Y(n_431) );
INVx2_ASAP7_75t_L g309 ( .A(n_117), .Y(n_309) );
INVx1_ASAP7_75t_L g356 ( .A(n_117), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_117), .B(n_310), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_118), .A2(n_260), .B1(n_408), .B2(n_982), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g1225 ( .A1(n_119), .A2(n_244), .B1(n_982), .B2(n_1226), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_119), .A2(n_244), .B1(n_1240), .B2(n_1241), .Y(n_1239) );
INVx1_ASAP7_75t_L g1089 ( .A(n_120), .Y(n_1089) );
INVx1_ASAP7_75t_L g627 ( .A(n_121), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g1106 ( .A1(n_122), .A2(n_151), .B1(n_921), .B2(n_1067), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g1120 ( .A1(n_122), .A2(n_226), .B1(n_991), .B2(n_1119), .Y(n_1120) );
INVx1_ASAP7_75t_L g1254 ( .A(n_125), .Y(n_1254) );
OAI22xp33_ASAP7_75t_L g1511 ( .A1(n_126), .A2(n_211), .B1(n_496), .B2(n_1059), .Y(n_1511) );
INVx1_ASAP7_75t_L g1532 ( .A(n_126), .Y(n_1532) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_127), .A2(n_167), .B1(n_794), .B2(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_129), .A2(n_193), .B1(n_921), .B2(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g934 ( .A(n_130), .Y(n_934) );
INVxp67_ASAP7_75t_SL g914 ( .A(n_131), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_131), .A2(n_237), .B1(n_710), .B2(n_938), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_132), .A2(n_254), .B1(n_574), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_132), .A2(n_239), .B1(n_589), .B2(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_133), .A2(n_246), .B1(n_1303), .B2(n_1306), .Y(n_1329) );
NOR2xp33_ASAP7_75t_L g1143 ( .A(n_134), .B(n_1044), .Y(n_1143) );
INVxp67_ASAP7_75t_SL g1170 ( .A(n_134), .Y(n_1170) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_135), .A2(n_136), .B1(n_1296), .B2(n_1311), .Y(n_1310) );
XNOR2xp5_ASAP7_75t_L g1508 ( .A(n_135), .B(n_1509), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_135), .A2(n_1551), .B1(n_1556), .B2(n_1559), .Y(n_1550) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_137), .A2(n_231), .B1(n_881), .B2(n_1012), .Y(n_1017) );
INVx1_ASAP7_75t_L g634 ( .A(n_139), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_140), .A2(n_184), .B1(n_921), .B2(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g868 ( .A(n_141), .Y(n_868) );
INVx1_ASAP7_75t_L g484 ( .A(n_142), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_143), .A2(n_153), .B1(n_1303), .B2(n_1306), .Y(n_1318) );
INVx1_ASAP7_75t_L g756 ( .A(n_144), .Y(n_756) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_145), .Y(n_721) );
INVx1_ASAP7_75t_L g925 ( .A(n_146), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_147), .A2(n_225), .B1(n_556), .B2(n_864), .C(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g344 ( .A(n_148), .Y(n_344) );
INVx1_ASAP7_75t_L g1142 ( .A(n_149), .Y(n_1142) );
INVx1_ASAP7_75t_L g1189 ( .A(n_150), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_151), .A2(n_261), .B1(n_990), .B2(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1191 ( .A(n_152), .Y(n_1191) );
INVx1_ASAP7_75t_L g1145 ( .A(n_154), .Y(n_1145) );
OAI322xp33_ASAP7_75t_L g1148 ( .A1(n_154), .A2(n_302), .A3(n_350), .B1(n_505), .B2(n_1149), .C1(n_1153), .C2(n_1159), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_155), .A2(n_952), .B1(n_1018), .B2(n_1019), .Y(n_951) );
INVxp67_ASAP7_75t_SL g1019 ( .A(n_155), .Y(n_1019) );
BUFx3_ASAP7_75t_L g316 ( .A(n_156), .Y(n_316) );
INVx1_ASAP7_75t_L g638 ( .A(n_157), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g865 ( .A1(n_158), .A2(n_264), .B1(n_543), .B2(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_158), .A2(n_200), .B1(n_746), .B2(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1129 ( .A(n_159), .Y(n_1129) );
INVx1_ASAP7_75t_L g1073 ( .A(n_160), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_161), .A2(n_163), .B1(n_1303), .B2(n_1306), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_162), .A2(n_177), .B1(n_796), .B2(n_918), .Y(n_1276) );
INVx1_ASAP7_75t_L g1523 ( .A(n_164), .Y(n_1523) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_165), .A2(n_233), .B1(n_1296), .B2(n_1311), .Y(n_1337) );
AOI211xp5_ASAP7_75t_SL g834 ( .A1(n_167), .A2(n_835), .B(n_836), .C(n_838), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_168), .Y(n_913) );
INVx1_ASAP7_75t_L g948 ( .A(n_169), .Y(n_948) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_170), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_171), .A2(n_202), .B1(n_798), .B2(n_800), .Y(n_797) );
INVx1_ASAP7_75t_L g821 ( .A(n_171), .Y(n_821) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_172), .A2(n_231), .B1(n_999), .B2(n_1000), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g869 ( .A1(n_173), .A2(n_204), .B1(n_870), .B2(n_873), .C(n_874), .Y(n_869) );
INVx1_ASAP7_75t_L g892 ( .A(n_173), .Y(n_892) );
OAI22xp33_ASAP7_75t_SL g855 ( .A1(n_175), .A2(n_217), .B1(n_393), .B2(n_720), .Y(n_855) );
INVx1_ASAP7_75t_L g895 ( .A(n_175), .Y(n_895) );
AOI21xp5_ASAP7_75t_SL g863 ( .A1(n_176), .A2(n_568), .B(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g878 ( .A(n_176), .Y(n_878) );
INVx1_ASAP7_75t_L g857 ( .A(n_178), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_178), .A2(n_264), .B1(n_746), .B2(n_886), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_179), .Y(n_862) );
INVx1_ASAP7_75t_L g894 ( .A(n_180), .Y(n_894) );
INVx1_ASAP7_75t_L g963 ( .A(n_181), .Y(n_963) );
OAI211xp5_ASAP7_75t_L g979 ( .A1(n_181), .A2(n_416), .B(n_672), .C(n_980), .Y(n_979) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_183), .A2(n_416), .B(n_418), .C(n_422), .Y(n_415) );
INVx1_ASAP7_75t_L g471 ( .A(n_183), .Y(n_471) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_184), .Y(n_1258) );
AOI21xp33_ASAP7_75t_L g555 ( .A1(n_185), .A2(n_556), .B(n_557), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_186), .Y(n_548) );
INVx1_ASAP7_75t_L g933 ( .A(n_187), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_188), .Y(n_1167) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_190), .Y(n_785) );
INVx1_ASAP7_75t_L g946 ( .A(n_191), .Y(n_946) );
XOR2x2_ASAP7_75t_L g1243 ( .A(n_192), .B(n_1244), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_193), .A2(n_243), .B1(n_542), .B2(n_819), .Y(n_1546) );
INVx1_ASAP7_75t_L g1138 ( .A(n_194), .Y(n_1138) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_195), .A2(n_234), .B1(n_248), .B2(n_487), .C1(n_503), .C2(n_512), .Y(n_486) );
INVx1_ASAP7_75t_L g1184 ( .A(n_196), .Y(n_1184) );
XOR2x2_ASAP7_75t_L g1179 ( .A(n_197), .B(n_1180), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_198), .A2(n_263), .B1(n_560), .B2(n_562), .Y(n_559) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_198), .Y(n_601) );
INVxp67_ASAP7_75t_L g884 ( .A(n_199), .Y(n_884) );
AOI21xp33_ASAP7_75t_L g858 ( .A1(n_200), .A2(n_568), .B(n_569), .Y(n_858) );
INVx1_ASAP7_75t_L g841 ( .A(n_202), .Y(n_841) );
INVx1_ASAP7_75t_L g1223 ( .A(n_203), .Y(n_1223) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_204), .Y(n_897) );
INVx1_ASAP7_75t_L g335 ( .A(n_205), .Y(n_335) );
INVx1_ASAP7_75t_L g632 ( .A(n_206), .Y(n_632) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_208), .A2(n_216), .B1(n_918), .B2(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g630 ( .A(n_209), .Y(n_630) );
INVx1_ASAP7_75t_L g647 ( .A(n_210), .Y(n_647) );
INVx1_ASAP7_75t_L g1531 ( .A(n_211), .Y(n_1531) );
INVx1_ASAP7_75t_L g947 ( .A(n_212), .Y(n_947) );
INVx1_ASAP7_75t_L g745 ( .A(n_213), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_215), .Y(n_736) );
INVx1_ASAP7_75t_L g898 ( .A(n_217), .Y(n_898) );
INVx1_ASAP7_75t_L g349 ( .A(n_220), .Y(n_349) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_221), .A2(n_235), .B1(n_621), .B2(n_622), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_221), .A2(n_235), .B1(n_435), .B2(n_679), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g1083 ( .A(n_222), .B(n_1084), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_223), .Y(n_527) );
INVx1_ASAP7_75t_L g1194 ( .A(n_224), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_225), .Y(n_1072) );
AOI22xp33_ASAP7_75t_SL g1110 ( .A1(n_226), .A2(n_261), .B1(n_794), .B2(n_1010), .Y(n_1110) );
OAI211xp5_ASAP7_75t_L g1246 ( .A1(n_227), .A2(n_1247), .B(n_1248), .C(n_1252), .Y(n_1246) );
INVx1_ASAP7_75t_L g1088 ( .A(n_228), .Y(n_1088) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_229), .Y(n_1154) );
BUFx3_ASAP7_75t_L g293 ( .A(n_232), .Y(n_293) );
INVx1_ASAP7_75t_L g447 ( .A(n_232), .Y(n_447) );
INVxp67_ASAP7_75t_SL g927 ( .A(n_237), .Y(n_927) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_238), .Y(n_717) );
INVx1_ASAP7_75t_L g708 ( .A(n_239), .Y(n_708) );
INVx1_ASAP7_75t_L g430 ( .A(n_240), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_240), .A2(n_460), .B(n_463), .C(n_472), .Y(n_459) );
INVx1_ASAP7_75t_L g843 ( .A(n_241), .Y(n_843) );
INVx1_ASAP7_75t_L g644 ( .A(n_242), .Y(n_644) );
INVx1_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
INVx1_ASAP7_75t_L g355 ( .A(n_247), .Y(n_355) );
INVx2_ASAP7_75t_L g368 ( .A(n_247), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_248), .A2(n_250), .B1(n_572), .B2(n_576), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_249), .Y(n_737) );
INVx1_ASAP7_75t_L g533 ( .A(n_250), .Y(n_533) );
INVx1_ASAP7_75t_L g848 ( .A(n_251), .Y(n_848) );
INVx1_ASAP7_75t_L g1094 ( .A(n_253), .Y(n_1094) );
INVx1_ASAP7_75t_L g772 ( .A(n_254), .Y(n_772) );
INVx1_ASAP7_75t_L g770 ( .A(n_255), .Y(n_770) );
INVx1_ASAP7_75t_L g1282 ( .A(n_256), .Y(n_1282) );
INVx1_ASAP7_75t_L g1037 ( .A(n_257), .Y(n_1037) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_258), .Y(n_791) );
INVx1_ASAP7_75t_L g1091 ( .A(n_259), .Y(n_1091) );
INVx1_ASAP7_75t_L g961 ( .A(n_260), .Y(n_961) );
XOR2x2_ASAP7_75t_L g298 ( .A(n_262), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g591 ( .A(n_263), .Y(n_591) );
INVx1_ASAP7_75t_L g957 ( .A(n_266), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_294), .B(n_1289), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx4f_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_279), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_273), .B(n_282), .Y(n_1549) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_275), .B(n_278), .Y(n_1555) );
INVx1_ASAP7_75t_L g1562 ( .A(n_275), .Y(n_1562) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_278), .B(n_1562), .Y(n_1564) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g478 ( .A(n_282), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g403 ( .A(n_283), .B(n_293), .Y(n_403) );
AND2x4_ASAP7_75t_L g558 ( .A(n_283), .B(n_292), .Y(n_558) );
INVx1_ASAP7_75t_L g618 ( .A(n_284), .Y(n_618) );
INVxp67_ASAP7_75t_SL g972 ( .A(n_284), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_284), .A2(n_445), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
AND2x4_ASAP7_75t_SL g1548 ( .A(n_284), .B(n_1549), .Y(n_1548) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x6_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
INVx1_ASAP7_75t_L g398 ( .A(n_286), .Y(n_398) );
OR2x6_ASAP7_75t_L g453 ( .A(n_286), .B(n_446), .Y(n_453) );
INVxp67_ASAP7_75t_L g1186 ( .A(n_286), .Y(n_1186) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx4f_ASAP7_75t_L g373 ( .A(n_287), .Y(n_373) );
INVx3_ASAP7_75t_L g710 ( .A(n_287), .Y(n_710) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx2_ASAP7_75t_L g380 ( .A(n_289), .Y(n_380) );
INVx2_ASAP7_75t_L g386 ( .A(n_289), .Y(n_386) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_289), .B(n_290), .Y(n_389) );
AND2x2_ASAP7_75t_L g448 ( .A(n_289), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g470 ( .A(n_289), .Y(n_470) );
AND2x2_ASAP7_75t_L g476 ( .A(n_289), .B(n_290), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_290), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g385 ( .A(n_290), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g449 ( .A(n_290), .Y(n_449) );
BUFx2_ASAP7_75t_L g466 ( .A(n_290), .Y(n_466) );
INVx1_ASAP7_75t_L g495 ( .A(n_290), .Y(n_495) );
AND2x2_ASAP7_75t_L g563 ( .A(n_290), .B(n_380), .Y(n_563) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g474 ( .A(n_292), .Y(n_474) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g458 ( .A(n_293), .Y(n_458) );
AND2x4_ASAP7_75t_L g468 ( .A(n_293), .B(n_469), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_1020), .B1(n_1021), .B2(n_1288), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g1288 ( .A(n_296), .Y(n_1288) );
XNOR2x1_ASAP7_75t_L g296 ( .A(n_297), .B(n_682), .Y(n_296) );
XNOR2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_481), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_406), .C(n_442), .Y(n_299) );
NOR2xp33_ASAP7_75t_SL g300 ( .A(n_301), .B(n_364), .Y(n_300) );
OAI33xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_311), .A3(n_326), .B1(n_340), .B2(n_350), .B3(n_357), .Y(n_301) );
OAI33xp33_ASAP7_75t_L g625 ( .A1(n_302), .A2(n_626), .A3(n_631), .B1(n_636), .B2(n_640), .B3(n_643), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_302), .A2(n_876), .B1(n_882), .B2(n_887), .Y(n_875) );
BUFx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_304), .Y(n_1064) );
BUFx8_ASAP7_75t_L g1204 ( .A(n_304), .Y(n_1204) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
INVx1_ASAP7_75t_L g405 ( .A(n_305), .Y(n_405) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_305), .Y(n_441) );
OR2x2_ASAP7_75t_L g501 ( .A(n_305), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g480 ( .A(n_306), .Y(n_480) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g775 ( .A(n_308), .Y(n_775) );
NAND2xp33_ASAP7_75t_SL g308 ( .A(n_309), .B(n_310), .Y(n_308) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_309), .Y(n_439) );
INVx1_ASAP7_75t_L g517 ( .A(n_309), .Y(n_517) );
AND3x4_ASAP7_75t_L g605 ( .A(n_309), .B(n_425), .C(n_583), .Y(n_605) );
INVx3_ASAP7_75t_L g353 ( .A(n_310), .Y(n_353) );
BUFx3_ASAP7_75t_L g425 ( .A(n_310), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_319), .B2(n_320), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_312), .A2(n_359), .B1(n_371), .B2(n_374), .Y(n_370) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_314), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_314), .A2(n_601), .B1(n_602), .B2(n_603), .Y(n_600) );
BUFx4f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x4_ASAP7_75t_L g410 ( .A(n_315), .B(n_353), .Y(n_410) );
OR2x4_ASAP7_75t_L g413 ( .A(n_315), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g498 ( .A(n_315), .Y(n_498) );
BUFx3_ASAP7_75t_L g764 ( .A(n_315), .Y(n_764) );
BUFx3_ASAP7_75t_L g1157 ( .A(n_315), .Y(n_1157) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_316), .Y(n_325) );
INVx2_ASAP7_75t_L g334 ( .A(n_316), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_316), .B(n_324), .Y(n_339) );
AND2x4_ASAP7_75t_L g420 ( .A(n_316), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g515 ( .A(n_317), .Y(n_515) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVxp67_ASAP7_75t_L g333 ( .A(n_318), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_319), .A2(n_363), .B1(n_374), .B2(n_391), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_320), .A2(n_1154), .B1(n_1155), .B2(n_1158), .Y(n_1153) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g646 ( .A(n_321), .Y(n_646) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
BUFx2_ASAP7_75t_L g1210 ( .A(n_322), .Y(n_1210) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
BUFx2_ASAP7_75t_L g429 ( .A(n_323), .Y(n_429) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g421 ( .A(n_324), .Y(n_421) );
BUFx2_ASAP7_75t_L g426 ( .A(n_325), .Y(n_426) );
INVx2_ASAP7_75t_L g524 ( .A(n_325), .Y(n_524) );
AND2x4_ASAP7_75t_L g589 ( .A(n_325), .B(n_532), .Y(n_589) );
OAI22xp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_328), .B1(n_335), .B2(n_336), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_327), .A2(n_344), .B1(n_382), .B2(n_387), .Y(n_381) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_329), .A2(n_736), .B1(n_737), .B2(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx5_ASAP7_75t_L g587 ( .A(n_331), .Y(n_587) );
INVx2_ASAP7_75t_SL g799 ( .A(n_331), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_331), .A2(n_794), .B1(n_894), .B2(n_895), .Y(n_893) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g343 ( .A(n_332), .Y(n_343) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_332), .Y(n_434) );
BUFx8_ASAP7_75t_L g599 ( .A(n_332), .Y(n_599) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x4_ASAP7_75t_L g514 ( .A(n_334), .B(n_515), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_335), .A2(n_349), .B1(n_395), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_337), .Y(n_1215) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x6_ASAP7_75t_L g436 ( .A(n_338), .B(n_353), .Y(n_436) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_345), .B2(n_349), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g1071 ( .A(n_342), .Y(n_1071) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g507 ( .A(n_343), .Y(n_507) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_343), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_345), .A2(n_627), .B1(n_628), .B2(n_630), .Y(n_626) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g417 ( .A(n_348), .Y(n_417) );
OR2x2_ASAP7_75t_L g537 ( .A(n_348), .B(n_501), .Y(n_537) );
INVx4_ASAP7_75t_L g595 ( .A(n_348), .Y(n_595) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_351), .A2(n_585), .B1(n_596), .B2(n_604), .C(n_606), .Y(n_584) );
INVx2_ASAP7_75t_L g887 ( .A(n_351), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_351), .B(n_1014), .C(n_1017), .Y(n_1013) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g642 ( .A(n_352), .Y(n_642) );
OAI33xp33_ASAP7_75t_L g1203 ( .A1(n_352), .A2(n_1204), .A3(n_1205), .B1(n_1211), .B2(n_1212), .B3(n_1216), .Y(n_1203) );
NAND3x1_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .C(n_356), .Y(n_352) );
INVx1_ASAP7_75t_L g414 ( .A(n_353), .Y(n_414) );
AND2x4_ASAP7_75t_L g419 ( .A(n_353), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g516 ( .A(n_353), .B(n_517), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g766 ( .A(n_353), .B(n_356), .Y(n_766) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g526 ( .A(n_355), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_355), .B(n_493), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_360), .B2(n_363), .Y(n_357) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g635 ( .A(n_361), .Y(n_635) );
CKINVDCx8_ASAP7_75t_R g771 ( .A(n_361), .Y(n_771) );
INVx1_ASAP7_75t_L g1161 ( .A(n_361), .Y(n_1161) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g536 ( .A(n_362), .Y(n_536) );
OAI33xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_370), .A3(n_381), .B1(n_390), .B2(n_394), .B3(n_401), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g649 ( .A(n_366), .Y(n_649) );
INVx4_ASAP7_75t_L g996 ( .A(n_366), .Y(n_996) );
INVx2_ASAP7_75t_L g1114 ( .A(n_366), .Y(n_1114) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g779 ( .A(n_367), .Y(n_779) );
OR2x6_ASAP7_75t_L g805 ( .A(n_367), .B(n_766), .Y(n_805) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g583 ( .A(n_368), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_368), .B(n_552), .Y(n_728) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx3_ASAP7_75t_L g653 ( .A(n_373), .Y(n_653) );
INVx4_ASAP7_75t_L g840 ( .A(n_373), .Y(n_840) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g1183 ( .A1(n_376), .A2(n_1184), .B1(n_1185), .B2(n_1187), .Y(n_1183) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx4_ASAP7_75t_L g656 ( .A(n_377), .Y(n_656) );
INVx2_ASAP7_75t_L g712 ( .A(n_377), .Y(n_712) );
INVx2_ASAP7_75t_L g938 ( .A(n_377), .Y(n_938) );
BUFx6f_ASAP7_75t_L g1202 ( .A(n_377), .Y(n_1202) );
INVx8_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g457 ( .A(n_378), .B(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g1259 ( .A(n_378), .Y(n_1259) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g1190 ( .A(n_383), .Y(n_1190) );
INVx4_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g393 ( .A(n_385), .Y(n_393) );
INVx2_ASAP7_75t_L g659 ( .A(n_385), .Y(n_659) );
INVx1_ASAP7_75t_L g719 ( .A(n_385), .Y(n_719) );
AND2x2_ASAP7_75t_L g494 ( .A(n_386), .B(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_386), .Y(n_550) );
BUFx4f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx4_ASAP7_75t_L g400 ( .A(n_388), .Y(n_400) );
BUFx4f_ASAP7_75t_L g660 ( .A(n_388), .Y(n_660) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_388), .Y(n_720) );
OR2x6_ASAP7_75t_L g725 ( .A(n_388), .B(n_726), .Y(n_725) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_388), .Y(n_874) );
OAI221xp5_ASAP7_75t_L g945 ( .A1(n_388), .A2(n_393), .B1(n_403), .B2(n_946), .C(n_947), .Y(n_945) );
BUFx4f_ASAP7_75t_L g1192 ( .A(n_388), .Y(n_1192) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g462 ( .A(n_389), .Y(n_462) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g836 ( .A1(n_393), .A2(n_403), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g553 ( .A1(n_399), .A2(n_554), .B(n_555), .C(n_559), .Y(n_553) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g545 ( .A(n_400), .Y(n_545) );
INVx2_ASAP7_75t_L g566 ( .A(n_400), .Y(n_566) );
INVx2_ASAP7_75t_L g1544 ( .A(n_400), .Y(n_1544) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_402), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g997 ( .A(n_402), .B(n_998), .C(n_1004), .Y(n_997) );
AOI33xp33_ASAP7_75t_L g1111 ( .A1(n_402), .A2(n_1112), .A3(n_1115), .B1(n_1118), .B2(n_1120), .B3(n_1121), .Y(n_1111) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx4_ASAP7_75t_L g569 ( .A(n_403), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_403), .B(n_404), .Y(n_664) );
INVx1_ASAP7_75t_SL g1032 ( .A(n_403), .Y(n_1032) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI31xp33_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_415), .A3(n_431), .B(n_437), .Y(n_406) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_409), .A2(n_433), .B1(n_1091), .B2(n_1092), .Y(n_1104) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g669 ( .A(n_410), .Y(n_669) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g679 ( .A(n_412), .Y(n_679) );
INVx2_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g900 ( .A(n_413), .Y(n_900) );
BUFx3_ASAP7_75t_L g982 ( .A(n_413), .Y(n_982) );
AND2x4_ASAP7_75t_L g433 ( .A(n_414), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g603 ( .A(n_417), .Y(n_603) );
CKINVDCx8_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
CKINVDCx8_ASAP7_75t_R g672 ( .A(n_419), .Y(n_672) );
OAI31xp33_ASAP7_75t_L g888 ( .A1(n_419), .A2(n_889), .A3(n_899), .B(n_901), .Y(n_888) );
AOI211xp5_ASAP7_75t_L g1098 ( .A1(n_419), .A2(n_909), .B(n_1096), .C(n_1099), .Y(n_1098) );
BUFx2_ASAP7_75t_L g607 ( .A(n_420), .Y(n_607) );
BUFx3_ASAP7_75t_L g748 ( .A(n_420), .Y(n_748) );
BUFx2_ASAP7_75t_L g757 ( .A(n_420), .Y(n_757) );
INVx2_ASAP7_75t_L g803 ( .A(n_420), .Y(n_803) );
BUFx2_ASAP7_75t_L g886 ( .A(n_420), .Y(n_886) );
BUFx2_ASAP7_75t_L g921 ( .A(n_420), .Y(n_921) );
INVx1_ASAP7_75t_L g532 ( .A(n_421), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .B1(n_428), .B2(n_430), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_423), .A2(n_428), .B1(n_897), .B2(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g1100 ( .A(n_423), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_423), .A2(n_428), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
AND2x4_ASAP7_75t_L g428 ( .A(n_424), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g675 ( .A(n_424), .B(n_426), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g889 ( .A1(n_424), .A2(n_890), .B(n_893), .C(n_896), .Y(n_889) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_427), .A2(n_464), .B1(n_467), .B2(n_471), .Y(n_463) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_428), .Y(n_676) );
INVx1_ASAP7_75t_L g1101 ( .A(n_428), .Y(n_1101) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g670 ( .A(n_433), .Y(n_670) );
INVxp67_ASAP7_75t_L g976 ( .A(n_433), .Y(n_976) );
INVx2_ASAP7_75t_L g1220 ( .A(n_433), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_434), .Y(n_769) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_434), .Y(n_796) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g978 ( .A(n_436), .Y(n_978) );
INVx1_ASAP7_75t_L g1227 ( .A(n_436), .Y(n_1227) );
OAI31xp33_ASAP7_75t_L g666 ( .A1(n_437), .A2(n_667), .A3(n_671), .B(n_678), .Y(n_666) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_438), .B(n_440), .Y(n_437) );
AND2x2_ASAP7_75t_L g901 ( .A(n_438), .B(n_440), .Y(n_901) );
AND2x4_ASAP7_75t_L g983 ( .A(n_438), .B(n_440), .Y(n_983) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_438), .B(n_440), .Y(n_1228) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_450), .A3(n_459), .B(n_477), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_SL g619 ( .A(n_445), .Y(n_619) );
INVx4_ASAP7_75t_L g1231 ( .A(n_445), .Y(n_1231) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_448), .Y(n_511) );
BUFx3_ASAP7_75t_L g556 ( .A(n_448), .Y(n_556) );
INVx2_ASAP7_75t_L g704 ( .A(n_448), .Y(n_704) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_453), .Y(n_621) );
BUFx6f_ASAP7_75t_L g1240 ( .A(n_453), .Y(n_1240) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g623 ( .A(n_457), .Y(n_623) );
INVx1_ASAP7_75t_L g960 ( .A(n_457), .Y(n_960) );
AND2x4_ASAP7_75t_L g465 ( .A(n_458), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g956 ( .A(n_458), .B(n_543), .Y(n_956) );
AND2x2_ASAP7_75t_L g969 ( .A(n_458), .B(n_466), .Y(n_969) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g698 ( .A(n_462), .B(n_697), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_462), .B(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_462), .B(n_941), .Y(n_940) );
INVx2_ASAP7_75t_SL g1196 ( .A(n_462), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_464), .A2(n_467), .B1(n_615), .B2(n_616), .Y(n_614) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g1093 ( .A1(n_465), .A2(n_835), .B1(n_964), .B2(n_1094), .C1(n_1095), .C2(n_1096), .Y(n_1093) );
BUFx2_ASAP7_75t_L g547 ( .A(n_466), .Y(n_547) );
INVx1_ASAP7_75t_L g732 ( .A(n_466), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_466), .A2(n_549), .B1(n_785), .B2(n_812), .Y(n_833) );
INVx1_ASAP7_75t_L g872 ( .A(n_466), .Y(n_872) );
BUFx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g965 ( .A(n_468), .Y(n_965) );
INVx2_ASAP7_75t_L g1237 ( .A(n_468), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_469), .B(n_552), .Y(n_734) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g970 ( .A(n_473), .Y(n_970) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_474), .B(n_993), .Y(n_1234) );
AND2x4_ASAP7_75t_SL g579 ( .A(n_475), .B(n_493), .Y(n_579) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_475), .Y(n_706) );
BUFx3_ASAP7_75t_L g835 ( .A(n_475), .Y(n_835) );
BUFx3_ASAP7_75t_L g967 ( .A(n_475), .Y(n_967) );
AND2x6_ASAP7_75t_L g1035 ( .A(n_475), .B(n_552), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_475), .Y(n_1052) );
INVx1_ASAP7_75t_L g1263 ( .A(n_475), .Y(n_1263) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g994 ( .A(n_476), .Y(n_994) );
BUFx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OAI31xp33_ASAP7_75t_L g612 ( .A1(n_478), .A2(n_613), .A3(n_617), .B(n_620), .Y(n_612) );
BUFx2_ASAP7_75t_L g973 ( .A(n_478), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_478), .A2(n_983), .B1(n_1086), .B2(n_1097), .Y(n_1085) );
BUFx3_ASAP7_75t_L g1242 ( .A(n_478), .Y(n_1242) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g491 ( .A(n_480), .Y(n_491) );
INVxp67_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
OR2x2_ASAP7_75t_L g733 ( .A(n_480), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AO22x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_608), .B1(n_609), .B2(n_681), .Y(n_482) );
INVx1_ASAP7_75t_SL g681 ( .A(n_483), .Y(n_681) );
XNOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_486), .B(n_519), .Y(n_485) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_490), .A2(n_509), .B1(n_736), .B2(n_737), .Y(n_735) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g509 ( .A(n_491), .B(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g1038 ( .A(n_492), .Y(n_1038) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g510 ( .A(n_493), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g573 ( .A(n_493), .B(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g826 ( .A(n_493), .Y(n_826) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_493), .B(n_860), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1040 ( .A(n_493), .B(n_511), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_494), .Y(n_543) );
INVx3_ASAP7_75t_L g561 ( .A(n_494), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_494), .B(n_552), .Y(n_693) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx2_ASAP7_75t_SL g629 ( .A(n_497), .Y(n_629) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_497), .B(n_499), .Y(n_1284) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g593 ( .A(n_498), .Y(n_593) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g506 ( .A(n_500), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g535 ( .A(n_501), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g788 ( .A(n_501), .Y(n_788) );
INVx1_ASAP7_75t_L g760 ( .A(n_502), .Y(n_760) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g883 ( .A(n_507), .Y(n_883) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_511), .Y(n_568) );
INVx2_ASAP7_75t_L g829 ( .A(n_511), .Y(n_829) );
INVx1_ASAP7_75t_L g1134 ( .A(n_511), .Y(n_1134) );
INVx5_ASAP7_75t_L g844 ( .A(n_512), .Y(n_844) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .Y(n_512) );
OR2x2_ASAP7_75t_L g1527 ( .A(n_513), .B(n_518), .Y(n_1527) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
INVx8_ASAP7_75t_L g747 ( .A(n_514), .Y(n_747) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_514), .Y(n_753) );
BUFx3_ASAP7_75t_L g908 ( .A(n_514), .Y(n_908) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_514), .Y(n_1068) );
AND2x4_ASAP7_75t_L g525 ( .A(n_516), .B(n_526), .Y(n_525) );
AND2x6_ASAP7_75t_L g741 ( .A(n_516), .B(n_523), .Y(n_741) );
AND2x2_ASAP7_75t_L g743 ( .A(n_516), .B(n_531), .Y(n_743) );
INVx1_ASAP7_75t_L g750 ( .A(n_516), .Y(n_750) );
NAND3xp33_ASAP7_75t_SL g519 ( .A(n_520), .B(n_538), .C(n_584), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_527), .B1(n_528), .B2(n_533), .C(n_534), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
AND2x4_ASAP7_75t_SL g811 ( .A(n_523), .B(n_525), .Y(n_811) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_523), .B(n_525), .Y(n_1281) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g528 ( .A(n_525), .B(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g606 ( .A(n_525), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_SL g813 ( .A(n_525), .B(n_529), .Y(n_813) );
OR2x2_ASAP7_75t_L g692 ( .A(n_526), .B(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_527), .A2(n_547), .B1(n_548), .B2(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g1062 ( .A(n_528), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_528), .A2(n_606), .B1(n_811), .B2(n_1138), .C(n_1170), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_528), .A2(n_1280), .B1(n_1281), .B2(n_1282), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_528), .A2(n_1281), .B1(n_1522), .B2(n_1523), .Y(n_1521) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g790 ( .A(n_535), .Y(n_790) );
AND2x4_ASAP7_75t_L g1078 ( .A(n_535), .B(n_692), .Y(n_1078) );
INVx2_ASAP7_75t_L g784 ( .A(n_537), .Y(n_784) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_537), .B(n_733), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_537), .B(n_733), .Y(n_1128) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_571), .B(n_580), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_553), .C(n_564), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_544), .C(n_551), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_SL g867 ( .A1(n_542), .A2(n_551), .B(n_868), .C(n_869), .Y(n_867) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g818 ( .A(n_543), .Y(n_818) );
A2O1A1Ixp33_ASAP7_75t_L g831 ( .A1(n_543), .A2(n_551), .B(n_791), .C(n_832), .Y(n_831) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_543), .A2(n_915), .B(n_940), .C(n_942), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_547), .A2(n_549), .B1(n_913), .B2(n_924), .Y(n_941) );
INVx1_ASAP7_75t_L g873 ( .A(n_549), .Y(n_873) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g943 ( .A(n_552), .Y(n_943) );
BUFx2_ASAP7_75t_L g987 ( .A(n_556), .Y(n_987) );
HB1xp67_ASAP7_75t_L g1536 ( .A(n_556), .Y(n_1536) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_558), .A2(n_566), .B1(n_821), .B2(n_822), .C(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g864 ( .A(n_558), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_558), .A2(n_566), .B1(n_658), .B2(n_933), .C(n_934), .Y(n_932) );
INVx3_ASAP7_75t_L g1264 ( .A(n_558), .Y(n_1264) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g723 ( .A(n_561), .Y(n_723) );
INVx1_ASAP7_75t_L g990 ( .A(n_561), .Y(n_990) );
INVx2_ASAP7_75t_L g1136 ( .A(n_561), .Y(n_1136) );
BUFx3_ASAP7_75t_L g988 ( .A(n_562), .Y(n_988) );
INVx1_ASAP7_75t_SL g1117 ( .A(n_562), .Y(n_1117) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g575 ( .A(n_563), .Y(n_575) );
BUFx3_ASAP7_75t_L g819 ( .A(n_563), .Y(n_819) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_563), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B(n_567), .C(n_570), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_565), .A2(n_591), .B1(n_592), .B2(n_594), .Y(n_590) );
BUFx3_ASAP7_75t_L g1119 ( .A(n_568), .Y(n_1119) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g695 ( .A(n_574), .B(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g866 ( .A(n_575), .Y(n_866) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g1042 ( .A(n_577), .Y(n_1042) );
INVx2_ASAP7_75t_L g1540 ( .A(n_577), .Y(n_1540) );
INVx4_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g1137 ( .A(n_579), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g1266 ( .A(n_581), .Y(n_1266) );
BUFx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI31xp33_ASAP7_75t_L g815 ( .A1(n_582), .A2(n_816), .A3(n_824), .B(n_834), .Y(n_815) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_582), .Y(n_851) );
OAI31xp33_ASAP7_75t_L g928 ( .A1(n_582), .A2(n_929), .A3(n_935), .B(n_944), .Y(n_928) );
BUFx2_ASAP7_75t_L g1147 ( .A(n_582), .Y(n_1147) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g633 ( .A(n_586), .Y(n_633) );
INVx8_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx3_ASAP7_75t_L g1151 ( .A(n_587), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_588), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
BUFx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx3_ASAP7_75t_L g800 ( .A(n_589), .Y(n_800) );
BUFx12f_ASAP7_75t_L g891 ( .A(n_589), .Y(n_891) );
INVx5_ASAP7_75t_L g919 ( .A(n_589), .Y(n_919) );
BUFx4f_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g763 ( .A(n_595), .Y(n_763) );
INVx1_ASAP7_75t_L g1217 ( .A(n_595), .Y(n_1217) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx3_ASAP7_75t_L g637 ( .A(n_599), .Y(n_637) );
AND2x4_ASAP7_75t_L g808 ( .A(n_599), .B(n_788), .Y(n_808) );
OAI211xp5_ASAP7_75t_L g773 ( .A1(n_603), .A2(n_717), .B(n_774), .C(n_776), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g1006 ( .A(n_604), .B(n_1007), .C(n_1011), .Y(n_1006) );
AOI33xp33_ASAP7_75t_L g1105 ( .A1(n_604), .A2(n_1106), .A3(n_1107), .B1(n_1108), .B2(n_1109), .B3(n_1110), .Y(n_1105) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI33xp33_ASAP7_75t_L g792 ( .A1(n_605), .A2(n_793), .A3(n_795), .B1(n_797), .B2(n_801), .B3(n_804), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g905 ( .A(n_605), .B(n_906), .C(n_907), .Y(n_905) );
AOI33xp33_ASAP7_75t_L g1272 ( .A1(n_605), .A2(n_804), .A3(n_1273), .B1(n_1276), .B2(n_1277), .B3(n_1278), .Y(n_1272) );
AOI33xp33_ASAP7_75t_L g1513 ( .A1(n_605), .A2(n_804), .A3(n_1514), .B1(n_1517), .B2(n_1519), .B3(n_1520), .Y(n_1513) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_606), .A2(n_811), .B1(n_812), .B2(n_813), .C(n_814), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_606), .A2(n_811), .B1(n_813), .B2(n_924), .C(n_925), .Y(n_923) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_606), .Y(n_1079) );
INVx3_ASAP7_75t_L g1286 ( .A(n_606), .Y(n_1286) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_624), .C(n_666), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_615), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g1241 ( .A(n_623), .Y(n_1241) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_648), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_627), .A2(n_644), .B1(n_651), .B2(n_654), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_628), .A2(n_644), .B1(n_645), .B2(n_647), .Y(n_643) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_630), .A2(n_647), .B1(n_658), .B2(n_660), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_632), .A2(n_638), .B1(n_658), .B2(n_660), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_634), .A2(n_639), .B1(n_651), .B2(n_654), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_635), .A2(n_1071), .B1(n_1072), .B2(n_1073), .C(n_1074), .Y(n_1070) );
INVx1_ASAP7_75t_L g1015 ( .A(n_637), .Y(n_1015) );
OAI22xp5_ASAP7_75t_SL g1063 ( .A1(n_640), .A2(n_1064), .B1(n_1065), .B2(n_1070), .Y(n_1063) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_642), .Y(n_1109) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI33xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .A3(n_657), .B1(n_661), .B2(n_662), .B3(n_665), .Y(n_648) );
INVx1_ASAP7_75t_L g714 ( .A(n_649), .Y(n_714) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g1046 ( .A1(n_654), .A2(n_1047), .B1(n_1049), .B2(n_1050), .C(n_1051), .Y(n_1046) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_656), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_838) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g823 ( .A(n_659), .Y(n_823) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_674), .A2(n_676), .B1(n_966), .B2(n_968), .Y(n_980) );
BUFx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
XNOR2x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_950), .Y(n_682) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_846), .B2(n_949), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XOR2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_780), .Y(n_685) );
XNOR2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND4xp75_ASAP7_75t_L g688 ( .A(n_689), .B(n_699), .C(n_735), .D(n_738), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI211x1_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_714), .B(n_715), .C(n_729), .Y(n_699) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g1250 ( .A(n_702), .Y(n_1250) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_703), .Y(n_999) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g1031 ( .A(n_704), .Y(n_1031) );
BUFx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_706), .A2(n_807), .B1(n_814), .B2(n_828), .C(n_830), .Y(n_827) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_706), .A2(n_828), .B1(n_911), .B2(n_925), .C(n_937), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_711), .B2(n_713), .Y(n_707) );
BUFx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_710), .Y(n_1048) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_713), .A2(n_721), .B1(n_763), .B2(n_764), .C(n_765), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_724), .B(n_725), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_718), .A2(n_1194), .B1(n_1195), .B2(n_1197), .Y(n_1193) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g856 ( .A1(n_720), .A2(n_857), .B(n_858), .C(n_859), .Y(n_856) );
OAI211xp5_ASAP7_75t_SL g861 ( .A1(n_720), .A2(n_862), .B(n_863), .C(n_865), .Y(n_861) );
OAI33xp33_ASAP7_75t_L g1182 ( .A1(n_724), .A2(n_1113), .A3(n_1183), .B1(n_1188), .B2(n_1193), .B3(n_1198), .Y(n_1182) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2x2_ASAP7_75t_L g730 ( .A(n_727), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI31xp67_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_751), .A3(n_761), .B(n_778), .Y(n_738) );
INVx4_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_748), .C(n_749), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g777 ( .A(n_747), .Y(n_777) );
INVx2_ASAP7_75t_L g787 ( .A(n_747), .Y(n_787) );
INVx8_ASAP7_75t_L g794 ( .A(n_747), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_748), .A2(n_868), .B1(n_891), .B2(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B(n_758), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI21xp5_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_767), .B(n_773), .Y(n_761) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_770), .B1(n_771), .B2(n_772), .Y(n_767) );
OAI221xp5_ASAP7_75t_L g1159 ( .A1(n_768), .A2(n_1160), .B1(n_1161), .B2(n_1162), .C(n_1163), .Y(n_1159) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_SL g877 ( .A(n_769), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_771), .A2(n_877), .B1(n_878), .B2(n_879), .C(n_880), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g882 ( .A1(n_771), .A2(n_862), .B1(n_883), .B2(n_884), .C(n_885), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_771), .A2(n_1150), .B1(n_1151), .B2(n_1152), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_771), .A2(n_883), .B1(n_1189), .B2(n_1199), .Y(n_1211) );
INVx1_ASAP7_75t_L g1053 ( .A(n_778), .Y(n_1053) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g780 ( .A(n_781), .B(n_845), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_809), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_792), .C(n_806), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_786), .B2(n_789), .C1(n_790), .C2(n_791), .Y(n_783) );
AOI222xp33_ASAP7_75t_L g912 ( .A1(n_784), .A2(n_786), .B1(n_790), .B2(n_913), .C1(n_914), .C2(n_915), .Y(n_912) );
AND2x4_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
AND2x4_ASAP7_75t_L g1173 ( .A(n_787), .B(n_788), .Y(n_1173) );
INVx1_ASAP7_75t_L g1213 ( .A(n_796), .Y(n_1213) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g881 ( .A(n_803), .Y(n_881) );
INVx1_ASAP7_75t_L g909 ( .A(n_803), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_804), .B(n_917), .C(n_920), .Y(n_916) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_808), .B(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g1059 ( .A(n_808), .Y(n_1059) );
NAND3xp33_ASAP7_75t_SL g809 ( .A(n_810), .B(n_815), .C(n_842), .Y(n_809) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_818), .Y(n_1034) );
OAI21xp33_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_827), .B(n_831), .Y(n_824) );
OAI21xp5_ASAP7_75t_SL g935 ( .A1(n_825), .A2(n_936), .B(n_939), .Y(n_935) );
INVxp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g853 ( .A1(n_826), .A2(n_854), .B(n_855), .Y(n_853) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_844), .B(n_927), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_844), .B(n_1146), .Y(n_1171) );
XNOR2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_902), .Y(n_846) );
XOR2xp5_ASAP7_75t_L g949 ( .A(n_847), .B(n_902), .Y(n_949) );
XNOR2x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
AND2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_888), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B(n_875), .Y(n_850) );
NAND4xp25_ASAP7_75t_L g852 ( .A(n_853), .B(n_856), .C(n_861), .D(n_867), .Y(n_852) );
INVx1_ASAP7_75t_L g931 ( .A(n_860), .Y(n_931) );
BUFx2_ASAP7_75t_L g1005 ( .A(n_860), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1538 ( .A(n_860), .Y(n_1538) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NOR2x1_ASAP7_75t_L g1045 ( .A(n_872), .B(n_943), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_886), .Y(n_1010) );
XNOR2x1_ASAP7_75t_L g902 ( .A(n_903), .B(n_948), .Y(n_902) );
OR2x2_ASAP7_75t_L g903 ( .A(n_904), .B(n_922), .Y(n_903) );
NAND4xp25_ASAP7_75t_SL g904 ( .A(n_905), .B(n_910), .C(n_912), .D(n_916), .Y(n_904) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_908), .Y(n_1012) );
INVx2_ASAP7_75t_SL g1275 ( .A(n_908), .Y(n_1275) );
INVx1_ASAP7_75t_L g1516 ( .A(n_908), .Y(n_1516) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g1016 ( .A(n_919), .Y(n_1016) );
INVx2_ASAP7_75t_R g1518 ( .A(n_919), .Y(n_1518) );
NAND3xp33_ASAP7_75t_SL g922 ( .A(n_923), .B(n_926), .C(n_928), .Y(n_922) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g1018 ( .A(n_952), .Y(n_1018) );
NAND3xp33_ASAP7_75t_L g952 ( .A(n_953), .B(n_974), .C(n_984), .Y(n_952) );
OAI21xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_971), .B(n_973), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_962), .C(n_970), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_957), .B1(n_958), .B2(n_961), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_956), .A2(n_960), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
AOI222xp33_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_964), .B1(n_966), .B2(n_967), .C1(n_968), .C2(n_969), .Y(n_962) );
INVx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_969), .A2(n_1223), .B1(n_1236), .B2(n_1238), .Y(n_1235) );
NAND4xp25_ASAP7_75t_L g1086 ( .A(n_970), .B(n_1087), .C(n_1090), .D(n_1093), .Y(n_1086) );
OAI31xp33_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_979), .A3(n_981), .B(n_983), .Y(n_974) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_978), .A2(n_1088), .B1(n_1089), .B2(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_982), .Y(n_1103) );
AND4x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_997), .C(n_1006), .D(n_1013), .Y(n_984) );
NAND3xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .C(n_995), .Y(n_985) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_994), .Y(n_1003) );
INVx2_ASAP7_75t_SL g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx2_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_SL g1020 ( .A(n_1021), .Y(n_1020) );
XNOR2xp5_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1177), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1080), .B1(n_1175), .B2(n_1176), .Y(n_1022) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1023), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
O2A1O1Ixp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1041), .B(n_1053), .C(n_1054), .Y(n_1025) );
INVx3_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_1028), .A2(n_1040), .B1(n_1145), .B2(n_1146), .Y(n_1144) );
INVx2_ASAP7_75t_SL g1247 ( .A(n_1028), .Y(n_1247) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1033), .B(n_1035), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_1035), .A2(n_1132), .B1(n_1135), .B2(n_1137), .C(n_1138), .Y(n_1131) );
AOI21xp5_ASAP7_75t_SL g1248 ( .A1(n_1035), .A2(n_1249), .B(n_1251), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g1534 ( .A1(n_1035), .A2(n_1535), .B(n_1537), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1038), .B1(n_1039), .B2(n_1040), .Y(n_1036) );
AOI221xp5_ASAP7_75t_SL g1139 ( .A1(n_1038), .A2(n_1140), .B1(n_1141), .B2(n_1142), .C(n_1143), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_1038), .A2(n_1253), .B1(n_1254), .B2(n_1255), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_1038), .A2(n_1531), .B1(n_1532), .B2(n_1533), .Y(n_1530) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1040), .Y(n_1255) );
BUFx6f_ASAP7_75t_L g1533 ( .A(n_1040), .Y(n_1533) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx2_ASAP7_75t_L g1541 ( .A(n_1045), .Y(n_1541) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_1047), .A2(n_1199), .B1(n_1200), .B2(n_1201), .Y(n_1198) );
OAI221xp5_ASAP7_75t_L g1257 ( .A1(n_1047), .A2(n_1258), .B1(n_1259), .B2(n_1260), .C(n_1261), .Y(n_1257) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
OAI21xp5_ASAP7_75t_L g1065 ( .A1(n_1049), .A2(n_1066), .B(n_1069), .Y(n_1065) );
NAND3xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1060), .C(n_1075), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1058), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1063), .Y(n_1060) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1068), .Y(n_1165) );
AOI21xp5_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1077), .B(n_1079), .Y(n_1075) );
AOI21xp5_ASAP7_75t_L g1166 ( .A1(n_1077), .A2(n_1167), .B(n_1168), .Y(n_1166) );
AOI21xp33_ASAP7_75t_SL g1267 ( .A1(n_1077), .A2(n_1268), .B(n_1269), .Y(n_1267) );
AOI21xp33_ASAP7_75t_L g1524 ( .A1(n_1077), .A2(n_1525), .B(n_1526), .Y(n_1524) );
INVx8_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1080), .Y(n_1176) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B1(n_1122), .B2(n_1123), .Y(n_1080) );
INVx1_ASAP7_75t_SL g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NAND3x1_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1105), .C(n_1111), .Y(n_1084) );
NAND3xp33_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1102), .C(n_1104), .Y(n_1097) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_SL g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
XNOR2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1174), .Y(n_1124) );
NAND2xp5_ASAP7_75t_SL g1125 ( .A(n_1126), .B(n_1166), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_1127), .A2(n_1129), .B1(n_1130), .B2(n_1147), .C(n_1148), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND3xp33_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1139), .C(n_1144), .Y(n_1130) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_1134), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1142), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVxp67_ASAP7_75t_SL g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1157), .Y(n_1207) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
NAND3xp33_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1171), .C(n_1172), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1177 ( .A1(n_1178), .A2(n_1179), .B1(n_1243), .B2(n_1287), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NAND3xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1218), .C(n_1229), .Y(n_1180) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1203), .Y(n_1181) );
OAI22xp33_ASAP7_75t_L g1205 ( .A1(n_1184), .A2(n_1194), .B1(n_1206), .B2(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OAI22xp33_ASAP7_75t_L g1216 ( .A1(n_1187), .A2(n_1197), .B1(n_1206), .B2(n_1217), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1190), .B1(n_1191), .B2(n_1192), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_1191), .A2(n_1200), .B1(n_1213), .B2(n_1214), .Y(n_1212) );
INVx5_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVx5_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx3_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
OAI31xp33_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1221), .A3(n_1225), .B(n_1228), .Y(n_1218) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
OAI31xp33_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1232), .A3(n_1239), .B(n_1242), .Y(n_1229) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1243), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1267), .C(n_1270), .Y(n_1244) );
OAI21xp33_ASAP7_75t_L g1245 ( .A1(n_1246), .A2(n_1256), .B(n_1265), .Y(n_1245) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OAI21xp5_ASAP7_75t_SL g1528 ( .A1(n_1265), .A2(n_1529), .B(n_1539), .Y(n_1528) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
NOR3xp33_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1283), .C(n_1285), .Y(n_1270) );
NAND2xp5_ASAP7_75t_SL g1271 ( .A(n_1272), .B(n_1279), .Y(n_1271) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
NOR3xp33_ASAP7_75t_L g1510 ( .A(n_1285), .B(n_1511), .C(n_1512), .Y(n_1510) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_1286), .Y(n_1285) );
OAI221xp5_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1503), .B1(n_1507), .B2(n_1547), .C(n_1550), .Y(n_1289) );
AND3x1_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1440), .C(n_1477), .Y(n_1290) );
AOI211xp5_ASAP7_75t_SL g1291 ( .A1(n_1292), .A2(n_1313), .B(n_1367), .C(n_1416), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1308), .Y(n_1293) );
INVx3_ASAP7_75t_L g1388 ( .A(n_1294), .Y(n_1388) );
A2O1A1Ixp33_ASAP7_75t_L g1406 ( .A1(n_1294), .A2(n_1407), .B(n_1408), .C(n_1409), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1294), .B(n_1366), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1302), .Y(n_1294) );
AND2x6_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1297), .B(n_1301), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1297), .B(n_1304), .Y(n_1303) );
AND2x6_ASAP7_75t_L g1306 ( .A(n_1297), .B(n_1307), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1297), .B(n_1301), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1297), .B(n_1301), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1299), .B(n_1305), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g1506 ( .A(n_1300), .Y(n_1506) );
OAI21xp5_ASAP7_75t_L g1561 ( .A1(n_1301), .A2(n_1562), .B(n_1563), .Y(n_1561) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1308), .Y(n_1379) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1308), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1308), .B(n_1348), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1308), .B(n_1415), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1308), .B(n_1330), .Y(n_1448) );
NAND3xp33_ASAP7_75t_L g1454 ( .A(n_1308), .B(n_1424), .C(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1309), .B(n_1366), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1309), .B(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1309), .Y(n_1385) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1309), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1309), .B(n_1330), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1312), .Y(n_1309) );
OAI211xp5_ASAP7_75t_SL g1313 ( .A1(n_1314), .A2(n_1324), .B(n_1338), .C(n_1355), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1320), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1449 ( .A(n_1316), .B(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1317), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1317), .B(n_1343), .Y(n_1352) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1317), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1382 ( .A(n_1317), .B(n_1342), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1317), .B(n_1321), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1317), .B(n_1320), .Y(n_1393) );
NAND2x1_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1320), .B(n_1351), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1320), .B(n_1360), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1320), .B(n_1363), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1320), .B(n_1352), .Y(n_1412) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1320), .B(n_1382), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1320), .B(n_1400), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1320), .B(n_1341), .Y(n_1461) );
INVx2_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1321), .B(n_1335), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1321), .B(n_1354), .Y(n_1353) );
AOI22xp5_ASAP7_75t_L g1355 ( .A1(n_1321), .A2(n_1356), .B1(n_1358), .B2(n_1362), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1321), .B(n_1346), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1321), .B(n_1423), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1321), .B(n_1342), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1321), .B(n_1382), .Y(n_1468) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1321), .B(n_1343), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1493 ( .A(n_1321), .B(n_1343), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1324 ( .A(n_1325), .B(n_1334), .Y(n_1324) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1325), .Y(n_1415) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1325), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1330), .Y(n_1325) );
INVx2_ASAP7_75t_L g1348 ( .A(n_1326), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1326), .B(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1327), .B(n_1330), .Y(n_1357) );
INVx2_ASAP7_75t_SL g1365 ( .A(n_1327), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1327), .B(n_1363), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1327), .B(n_1366), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1327), .B(n_1369), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1329), .Y(n_1327) );
CKINVDCx5p33_ASAP7_75t_R g1366 ( .A(n_1330), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1368 ( .A1(n_1330), .A2(n_1341), .B1(n_1369), .B2(n_1372), .C(n_1376), .Y(n_1368) );
AOI221xp5_ASAP7_75t_L g1389 ( .A1(n_1330), .A2(n_1343), .B1(n_1390), .B2(n_1394), .C(n_1397), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1330), .B(n_1335), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1330), .B(n_1497), .Y(n_1496) );
AND2x4_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1333), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1334), .B(n_1341), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1334), .B(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1334), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1334), .B(n_1434), .Y(n_1433) );
OAI211xp5_ASAP7_75t_L g1442 ( .A1(n_1334), .A2(n_1443), .B(n_1445), .C(n_1447), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_1334), .B(n_1476), .Y(n_1475) );
OR2x2_ASAP7_75t_L g1495 ( .A(n_1334), .B(n_1393), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_1335), .Y(n_1334) );
INVx3_ASAP7_75t_L g1363 ( .A(n_1335), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1335), .B(n_1379), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1335), .B(n_1374), .Y(n_1499) );
AND2x4_ASAP7_75t_SL g1335 ( .A(n_1336), .B(n_1337), .Y(n_1335) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_1339), .A2(n_1348), .B1(n_1349), .B2(n_1353), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1348), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1347), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1341), .B(n_1411), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1346), .Y(n_1341) );
OAI322xp33_ASAP7_75t_L g1376 ( .A1(n_1342), .A2(n_1348), .A3(n_1377), .B1(n_1380), .B2(n_1382), .C1(n_1383), .C2(n_1386), .Y(n_1376) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1360 ( .A(n_1343), .B(n_1361), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1345), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1347), .B(n_1400), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1347), .B(n_1352), .Y(n_1463) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1348), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1348), .B(n_1446), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1348), .B(n_1463), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1485 ( .A(n_1348), .B(n_1358), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1348), .B(n_1379), .Y(n_1502) );
O2A1O1Ixp33_ASAP7_75t_L g1486 ( .A1(n_1349), .A2(n_1487), .B(n_1489), .C(n_1490), .Y(n_1486) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1351), .B(n_1371), .Y(n_1370) );
OAI22xp5_ASAP7_75t_SL g1478 ( .A1(n_1351), .A2(n_1383), .B1(n_1479), .B2(n_1480), .Y(n_1478) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1356), .B(n_1384), .Y(n_1383) );
AOI322xp5_ASAP7_75t_L g1404 ( .A1(n_1356), .A2(n_1378), .A3(n_1405), .B1(n_1406), .B2(n_1410), .C1(n_1412), .C2(n_1413), .Y(n_1404) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1358), .B(n_1363), .Y(n_1501) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1360), .Y(n_1400) );
NOR2xp33_ASAP7_75t_L g1444 ( .A(n_1360), .B(n_1429), .Y(n_1444) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1364), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1395 ( .A(n_1363), .B(n_1396), .Y(n_1395) );
CKINVDCx14_ASAP7_75t_R g1427 ( .A(n_1363), .Y(n_1427) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1363), .B(n_1374), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1363), .B(n_1365), .Y(n_1455) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1364), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1366), .Y(n_1364) );
INVx2_ASAP7_75t_L g1374 ( .A(n_1365), .Y(n_1374) );
A2O1A1Ixp33_ASAP7_75t_L g1459 ( .A1(n_1365), .A2(n_1460), .B(n_1462), .C(n_1464), .Y(n_1459) );
A2O1A1Ixp33_ASAP7_75t_L g1491 ( .A1(n_1365), .A2(n_1432), .B(n_1492), .C(n_1494), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1366), .B(n_1388), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1366), .B(n_1426), .Y(n_1425) );
OAI221xp5_ASAP7_75t_SL g1367 ( .A1(n_1368), .A2(n_1387), .B1(n_1389), .B2(n_1401), .C(n_1404), .Y(n_1367) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1371), .Y(n_1411) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1375), .Y(n_1373) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_1374), .B(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1375), .Y(n_1409) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1381), .Y(n_1437) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1382), .Y(n_1424) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
CKINVDCx14_ASAP7_75t_R g1441 ( .A(n_1387), .Y(n_1441) );
OAI221xp5_ASAP7_75t_L g1465 ( .A1(n_1387), .A2(n_1466), .B1(n_1469), .B2(n_1470), .C(n_1471), .Y(n_1465) );
OAI31xp33_ASAP7_75t_SL g1477 ( .A1(n_1387), .A2(n_1478), .A3(n_1481), .B(n_1484), .Y(n_1477) );
CKINVDCx14_ASAP7_75t_R g1387 ( .A(n_1388), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1388), .B(n_1403), .Y(n_1402) );
AOI322xp5_ASAP7_75t_L g1421 ( .A1(n_1390), .A2(n_1422), .A3(n_1425), .B1(n_1427), .B2(n_1428), .C1(n_1431), .C2(n_1433), .Y(n_1421) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1396), .B(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1396), .B(n_1467), .Y(n_1470) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
NOR2xp33_ASAP7_75t_L g1423 ( .A(n_1400), .B(n_1424), .Y(n_1423) );
CKINVDCx14_ASAP7_75t_R g1401 ( .A(n_1402), .Y(n_1401) );
OR2x2_ASAP7_75t_L g1429 ( .A(n_1403), .B(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1405), .Y(n_1498) );
OAI211xp5_ASAP7_75t_SL g1484 ( .A1(n_1409), .A2(n_1485), .B(n_1486), .C(n_1500), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1411), .B(n_1424), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_1412), .B(n_1452), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1412), .B(n_1419), .Y(n_1483) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
OAI211xp5_ASAP7_75t_SL g1416 ( .A1(n_1417), .A2(n_1418), .B(n_1421), .C(n_1435), .Y(n_1416) );
INVxp67_ASAP7_75t_SL g1464 ( .A(n_1417), .Y(n_1464) );
INVxp67_ASAP7_75t_L g1446 ( .A(n_1418), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1420), .Y(n_1418) );
INVx2_ASAP7_75t_L g1452 ( .A(n_1420), .Y(n_1452) );
AOI221xp5_ASAP7_75t_SL g1447 ( .A1(n_1425), .A2(n_1448), .B1(n_1449), .B2(n_1452), .C(n_1453), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1426), .B(n_1436), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1427), .B(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1430), .Y(n_1476) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1432), .Y(n_1458) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1438), .Y(n_1436) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
AOI211xp5_ASAP7_75t_L g1440 ( .A1(n_1441), .A2(n_1442), .B(n_1456), .C(n_1465), .Y(n_1440) );
INVxp67_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
OAI21xp5_ASAP7_75t_L g1471 ( .A1(n_1452), .A2(n_1472), .B(n_1474), .Y(n_1471) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
OAI21xp5_ASAP7_75t_L g1456 ( .A1(n_1457), .A2(n_1458), .B(n_1459), .Y(n_1456) );
OAI21xp33_ASAP7_75t_L g1500 ( .A1(n_1460), .A2(n_1501), .B(n_1502), .Y(n_1500) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
NAND2xp5_ASAP7_75t_SL g1490 ( .A(n_1491), .B(n_1496), .Y(n_1490) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
NOR2xp33_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1499), .Y(n_1497) );
CKINVDCx20_ASAP7_75t_R g1503 ( .A(n_1504), .Y(n_1503) );
CKINVDCx20_ASAP7_75t_R g1504 ( .A(n_1505), .Y(n_1504) );
INVx4_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
HB1xp67_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
HB1xp67_ASAP7_75t_L g1558 ( .A(n_1509), .Y(n_1558) );
AND3x1_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1524), .C(n_1528), .Y(n_1509) );
NAND2xp5_ASAP7_75t_SL g1512 ( .A(n_1513), .B(n_1521), .Y(n_1512) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
OAI211xp5_ASAP7_75t_SL g1542 ( .A1(n_1543), .A2(n_1544), .B(n_1545), .C(n_1546), .Y(n_1542) );
CKINVDCx5p33_ASAP7_75t_R g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
HB1xp67_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
BUFx3_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVxp33_ASAP7_75t_SL g1556 ( .A(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
endmodule