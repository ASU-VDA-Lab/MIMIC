module fake_jpeg_12691_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_44),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_51),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_11),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_59),
.B1(n_48),
.B2(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_59),
.B1(n_54),
.B2(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_50),
.B1(n_46),
.B2(n_58),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_50),
.B1(n_58),
.B2(n_20),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_98),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_2),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_95),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_4),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_93),
.B1(n_94),
.B2(n_85),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_22),
.C(n_10),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_9),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_106),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_110),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_110),
.B1(n_33),
.B2(n_39),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_23),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_26),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_28),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_29),
.C(n_31),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_102),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_122),
.B(n_109),
.Y(n_133)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_129),
.C(n_118),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_134),
.B(n_129),
.C(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_126),
.B1(n_104),
.B2(n_107),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_124),
.Y(n_138)
);


endmodule