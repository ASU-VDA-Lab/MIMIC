module fake_jpeg_28859_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_6),
.B(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_14),
.B(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_27),
.A2(n_8),
.B1(n_1),
.B2(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_5),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_27),
.B1(n_29),
.B2(n_17),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_8),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_23),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_83),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_22),
.B1(n_17),
.B2(n_32),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_25),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_69),
.B1(n_74),
.B2(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_32),
.B1(n_28),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_31),
.B1(n_23),
.B2(n_0),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_41),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_12),
.B1(n_13),
.B2(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_86),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_94),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_23),
.B1(n_11),
.B2(n_12),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_105),
.B1(n_107),
.B2(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_10),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_108),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_11),
.Y(n_101)
);

OR2x6_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_62),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_23),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_12),
.B1(n_78),
.B2(n_52),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_52),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_111),
.B1(n_93),
.B2(n_96),
.Y(n_141)
);

OAI22x1_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_84),
.B1(n_56),
.B2(n_79),
.Y(n_111)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_124),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_77),
.B1(n_68),
.B2(n_61),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_98),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_77),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_123),
.B(n_86),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_61),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_137),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_118),
.B1(n_130),
.B2(n_133),
.C(n_143),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_89),
.C(n_96),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_142),
.C(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_109),
.B1(n_118),
.B2(n_126),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_93),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_128),
.B(n_112),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_94),
.C(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_101),
.Y(n_145)
);

OAI221xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_118),
.B1(n_119),
.B2(n_111),
.C(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_156),
.C(n_133),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_113),
.C(n_122),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_150),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_159),
.B1(n_136),
.B2(n_131),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_134),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_118),
.B1(n_123),
.B2(n_105),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_158),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_123),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_107),
.B1(n_102),
.B2(n_129),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_162),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_136),
.C(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_146),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_156),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_152),
.B(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_147),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_139),
.B(n_138),
.C(n_148),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_163),
.B(n_149),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_158),
.B(n_140),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_177),
.B(n_161),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_179),
.B(n_181),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_162),
.C(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_138),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_168),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_112),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_171),
.B1(n_165),
.B2(n_146),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_185),
.C(n_114),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_86),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_187),
.B1(n_68),
.B2(n_70),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_70),
.C(n_71),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_87),
.Y(n_190)
);


endmodule