module fake_jpeg_11943_n_469 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_15),
.B1(n_7),
.B2(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_17),
.B1(n_27),
.B2(n_43),
.Y(n_101)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_48),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_77),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_7),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_79),
.B(n_11),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_93),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_42),
.B(n_8),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_24),
.B1(n_33),
.B2(n_40),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_98),
.A2(n_111),
.B1(n_44),
.B2(n_36),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_101),
.A2(n_44),
.B1(n_36),
.B2(n_16),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_31),
.B1(n_40),
.B2(n_33),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_106),
.A2(n_120),
.B(n_126),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_33),
.B1(n_40),
.B2(n_37),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_113),
.B(n_128),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_31),
.B1(n_40),
.B2(n_33),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_31),
.B1(n_46),
.B2(n_30),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_17),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_28),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_81),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_17),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_50),
.B(n_28),
.Y(n_148)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_51),
.C(n_89),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_106),
.C(n_134),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_31),
.B1(n_46),
.B2(n_19),
.Y(n_158)
);

OAI22x1_ASAP7_75t_L g226 ( 
.A1(n_158),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_166),
.B1(n_168),
.B2(n_172),
.Y(n_210)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

BUFx24_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_111),
.A2(n_59),
.B1(n_87),
.B2(n_84),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_57),
.B1(n_82),
.B2(n_76),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_63),
.B1(n_74),
.B2(n_69),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_176),
.Y(n_215)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_178),
.Y(n_222)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_192),
.B1(n_199),
.B2(n_200),
.Y(n_205)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_182),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_117),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_105),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_195),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_19),
.B1(n_27),
.B2(n_43),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_149),
.A2(n_27),
.B1(n_43),
.B2(n_29),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_107),
.A2(n_29),
.B1(n_34),
.B2(n_16),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_64),
.B1(n_62),
.B2(n_61),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_194),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_108),
.A2(n_29),
.B1(n_44),
.B2(n_36),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_103),
.B(n_25),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_104),
.B1(n_123),
.B2(n_124),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_136),
.B(n_30),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_140),
.A2(n_16),
.B1(n_37),
.B2(n_18),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_139),
.B1(n_135),
.B2(n_121),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_126),
.B(n_120),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_6),
.C(n_14),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_142),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_212),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_221),
.B1(n_159),
.B2(n_181),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_146),
.B(n_96),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_132),
.B1(n_123),
.B2(n_104),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_220),
.B1(n_225),
.B2(n_179),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_171),
.B1(n_157),
.B2(n_132),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_169),
.A2(n_151),
.B1(n_129),
.B2(n_134),
.Y(n_221)
);

MAJx3_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_30),
.C(n_1),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_0),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_30),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_224),
.B(n_1),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_124),
.B1(n_151),
.B2(n_138),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_173),
.B1(n_180),
.B2(n_161),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_155),
.A2(n_12),
.B(n_15),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_234),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_159),
.A2(n_30),
.B(n_135),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_121),
.B(n_37),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_165),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_259),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_174),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_178),
.B1(n_175),
.B2(n_170),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_153),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_267),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_255),
.B1(n_272),
.B2(n_224),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_203),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_269),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_254),
.A2(n_203),
.B1(n_236),
.B2(n_235),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_154),
.B1(n_201),
.B2(n_199),
.Y(n_255)
);

XOR2x2_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_241),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_177),
.B1(n_176),
.B2(n_198),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_257),
.A2(n_246),
.B(n_263),
.Y(n_308)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_167),
.B1(n_37),
.B2(n_18),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_264),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_164),
.B1(n_156),
.B2(n_165),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_204),
.Y(n_265)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_30),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_212),
.B(n_6),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_271),
.C(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_1),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_2),
.C(n_3),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_210),
.A2(n_205),
.B1(n_207),
.B2(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_9),
.B1(n_14),
.B2(n_5),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_14),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_2),
.C(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_215),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_234),
.B(n_226),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_278),
.A2(n_283),
.B(n_299),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_256),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_226),
.B1(n_221),
.B2(n_213),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_289),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_248),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_294),
.A2(n_296),
.B1(n_298),
.B2(n_307),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_262),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_300),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_297),
.B(n_4),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_210),
.B1(n_218),
.B2(n_237),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_244),
.A2(n_203),
.B(n_239),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_229),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_309),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_203),
.B(n_231),
.Y(n_305)
);

OAI31xp33_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_261),
.A3(n_245),
.B(n_265),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_255),
.A2(n_229),
.B1(n_236),
.B2(n_208),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_287),
.B1(n_301),
.B2(n_278),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_260),
.B(n_206),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_312),
.A2(n_304),
.B1(n_280),
.B2(n_290),
.Y(n_362)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_296),
.A2(n_264),
.B1(n_270),
.B2(n_275),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_332),
.B1(n_338),
.B2(n_301),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_335),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_277),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_323),
.C(n_327),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_298),
.A2(n_260),
.B1(n_266),
.B2(n_247),
.Y(n_320)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_320),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_322),
.A2(n_279),
.B(n_301),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_288),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_306),
.A2(n_245),
.B1(n_261),
.B2(n_271),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_324),
.A2(n_299),
.B(n_305),
.Y(n_346)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_333),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_268),
.C(n_250),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_257),
.B1(n_274),
.B2(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_258),
.Y(n_331)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_283),
.A2(n_278),
.B1(n_287),
.B2(n_289),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_309),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_341),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_339),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_257),
.B1(n_249),
.B2(n_236),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_337),
.A2(n_307),
.B1(n_308),
.B2(n_294),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_306),
.A2(n_257),
.B1(n_233),
.B2(n_231),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_295),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_208),
.C(n_206),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_314),
.Y(n_370)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_349),
.A2(n_352),
.B1(n_353),
.B2(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_351),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_321),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_312),
.A2(n_308),
.B1(n_279),
.B2(n_285),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_315),
.A2(n_337),
.B1(n_331),
.B2(n_324),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_291),
.Y(n_354)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_315),
.A2(n_292),
.B1(n_301),
.B2(n_311),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_340),
.B1(n_336),
.B2(n_328),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_332),
.A2(n_292),
.B1(n_311),
.B2(n_297),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_362),
.B1(n_293),
.B2(n_238),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_329),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_364),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

AO22x1_ASAP7_75t_L g365 ( 
.A1(n_314),
.A2(n_322),
.B1(n_338),
.B2(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_313),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_368),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_327),
.C(n_335),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_376),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_357),
.B(n_333),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_361),
.C(n_354),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_319),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_385),
.C(n_390),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_304),
.B1(n_284),
.B2(n_339),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_375),
.A2(n_382),
.B1(n_360),
.B2(n_358),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_323),
.C(n_341),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_367),
.C(n_346),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_380),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_280),
.C(n_317),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_280),
.C(n_316),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_383),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_325),
.C(n_284),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_290),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_293),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_349),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_293),
.C(n_233),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_393),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_377),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_397),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_390),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_365),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_399),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_400),
.B(n_407),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_344),
.B1(n_348),
.B2(n_343),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_384),
.A2(n_351),
.B1(n_366),
.B2(n_364),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_404),
.A2(n_374),
.B1(n_379),
.B2(n_347),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_383),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_406),
.B(n_409),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_359),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_369),
.C(n_381),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_412),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_378),
.C(n_380),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_393),
.A2(n_391),
.B(n_365),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_415),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_385),
.C(n_387),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_405),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_417),
.A2(n_420),
.B1(n_422),
.B2(n_344),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_396),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_399),
.A2(n_363),
.B(n_370),
.C(n_361),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_379),
.C(n_368),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_403),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_397),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_233),
.Y(n_436)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_427),
.B(n_428),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_407),
.C(n_396),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_421),
.A2(n_400),
.B1(n_403),
.B2(n_355),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_415),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_355),
.C(n_348),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_433),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_416),
.Y(n_433)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_414),
.B(n_343),
.CI(n_235),
.CON(n_434),
.SN(n_434)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_422),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_238),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_418),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_436),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_227),
.C(n_4),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_418),
.C(n_6),
.Y(n_446)
);

NAND2x1p5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_437),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_425),
.B(n_428),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_442),
.B(n_429),
.Y(n_452)
);

A2O1A1O1Ixp25_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_413),
.B(n_420),
.C(n_424),
.D(n_417),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_426),
.B(n_431),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_446),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_447),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_432),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_452),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_454),
.A2(n_456),
.B(n_439),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_455),
.A2(n_439),
.B(n_448),
.Y(n_457)
);

AOI21x1_ASAP7_75t_L g456 ( 
.A1(n_445),
.A2(n_434),
.B(n_227),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g462 ( 
.A1(n_457),
.A2(n_458),
.B(n_453),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_440),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_459),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_462),
.B(n_443),
.C(n_9),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_451),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_463),
.A2(n_443),
.B(n_12),
.Y(n_465)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_465),
.B(n_461),
.C(n_13),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_5),
.B(n_13),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_13),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_15),
.Y(n_469)
);


endmodule