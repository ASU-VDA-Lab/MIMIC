module fake_jpeg_4211_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_31),
.B(n_34),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_60),
.Y(n_67)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_30),
.Y(n_60)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_80),
.B1(n_54),
.B2(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_74),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_24),
.B1(n_17),
.B2(n_38),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_46),
.B1(n_55),
.B2(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_75),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_28),
.B(n_23),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_56),
.C(n_22),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_24),
.B1(n_28),
.B2(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_28),
.B1(n_31),
.B2(n_20),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_70),
.B1(n_65),
.B2(n_66),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_71),
.B(n_74),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_106),
.B(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_99),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_51),
.B1(n_82),
.B2(n_75),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_63),
.B1(n_58),
.B2(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_25),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_47),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_55),
.B1(n_51),
.B2(n_50),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_31),
.B1(n_36),
.B2(n_33),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_18),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_18),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_69),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_72),
.B1(n_67),
.B2(n_36),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_106),
.B(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_124),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_70),
.B1(n_73),
.B2(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_51),
.B1(n_73),
.B2(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_12),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_126),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_97),
.C(n_90),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_102),
.C(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_35),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_35),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_35),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_101),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_107),
.B(n_94),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_145),
.Y(n_177)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_155),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_159),
.B(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_86),
.C(n_92),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_86),
.C(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_129),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_89),
.C(n_53),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_125),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_112),
.A2(n_85),
.B(n_91),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_133),
.B(n_110),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_168),
.B1(n_153),
.B2(n_148),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_180),
.B(n_186),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_131),
.B(n_132),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_145),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_175),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_176),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_113),
.B1(n_117),
.B2(n_114),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_181),
.B1(n_182),
.B2(n_157),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_123),
.B1(n_114),
.B2(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_171),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_122),
.B(n_116),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_135),
.A2(n_123),
.B1(n_128),
.B2(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_184),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_157),
.C(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_136),
.A2(n_126),
.B1(n_119),
.B2(n_84),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_149),
.B1(n_144),
.B2(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_109),
.B1(n_100),
.B2(n_52),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_139),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_109),
.B(n_82),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_137),
.B1(n_148),
.B2(n_140),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_201),
.B1(n_209),
.B2(n_186),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_179),
.CI(n_163),
.CON(n_224),
.SN(n_224)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_140),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_203),
.C(n_211),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_158),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_205),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_142),
.C(n_137),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_142),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_208),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_212),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_158),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_158),
.B1(n_143),
.B2(n_84),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_18),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_45),
.C(n_52),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_177),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_224),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_27),
.B1(n_22),
.B2(n_15),
.Y(n_252)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_199),
.B(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_189),
.B(n_26),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_183),
.C(n_45),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_234),
.C(n_212),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_26),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_204),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_231),
.B(n_197),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_188),
.A2(n_16),
.B(n_27),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_82),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_75),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_45),
.C(n_52),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_215),
.B(n_210),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_240),
.C(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_253),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_242),
.B(n_219),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_209),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_217),
.C(n_215),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_198),
.C(n_188),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_187),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_191),
.C(n_206),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_240),
.C(n_235),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_202),
.B1(n_100),
.B2(n_16),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_222),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_19),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_19),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_218),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_260),
.B(n_262),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_236),
.B(n_232),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_257),
.B(n_265),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_243),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_263),
.B(n_1),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_227),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_18),
.C(n_3),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_224),
.A3(n_27),
.B1(n_22),
.B2(n_36),
.C1(n_15),
.C2(n_19),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_25),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_224),
.B(n_2),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_271),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.C(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_25),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_18),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_282),
.C(n_286),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_19),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_18),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_271),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_19),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_289),
.B(n_25),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_279),
.A2(n_257),
.B1(n_9),
.B2(n_11),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_2),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_8),
.C(n_12),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_8),
.C(n_11),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_9),
.C(n_3),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_9),
.Y(n_303)
);

A2O1A1O1Ixp25_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_277),
.B(n_282),
.C(n_286),
.D(n_281),
.Y(n_301)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_304),
.B(n_306),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_19),
.Y(n_304)
);

OAI21x1_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_287),
.B(n_288),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_293),
.C(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_2),
.C(n_3),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_300),
.B(n_19),
.C(n_6),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_315),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_311),
.C2(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.C(n_5),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_5),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_5),
.Y(n_319)
);


endmodule