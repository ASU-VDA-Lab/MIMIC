module fake_jpeg_3002_n_95 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_48),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_34),
.C(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_1),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_39),
.B1(n_41),
.B2(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_29),
.B1(n_38),
.B2(n_42),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_2),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_38),
.Y(n_59)
);

BUFx24_ASAP7_75t_SL g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_42),
.C(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_59),
.B1(n_29),
.B2(n_5),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_78),
.B1(n_26),
.B2(n_9),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_15),
.Y(n_75)
);

AO21x2_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_13),
.B(n_24),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_16),
.B(n_18),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_12),
.B1(n_22),
.B2(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_76),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_17),
.B(n_19),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_81),
.A3(n_76),
.B1(n_85),
.B2(n_82),
.C(n_77),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_88),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_75),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_87),
.B(n_78),
.C(n_10),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_8),
.Y(n_95)
);


endmodule