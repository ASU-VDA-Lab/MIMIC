module fake_netlist_6_17_n_2110 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2110);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2110;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_92),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_147),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_47),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_121),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_109),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_37),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_15),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_141),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_71),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_53),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_44),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_107),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_60),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_131),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_21),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_106),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_4),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_203),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_89),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_62),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_207),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_98),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_187),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_174),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_122),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_100),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_25),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_145),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_9),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_87),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_47),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_69),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_66),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_137),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_86),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_96),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_59),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_148),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_84),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_25),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_170),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_196),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_50),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_179),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_167),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_119),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_85),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_11),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_81),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_88),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_162),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_159),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_197),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_143),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_82),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_20),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_195),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_31),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_172),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_152),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_0),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_52),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_16),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_200),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_36),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_161),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_129),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_12),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_102),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_166),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_16),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_33),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_184),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_110),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_177),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_130),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_17),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_83),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_115),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_144),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_180),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_59),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_81),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_90),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_123),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_210),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_118),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_14),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_76),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_27),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_139),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_60),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_84),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_114),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_95),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_45),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_94),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_82),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_175),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_55),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_51),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_61),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_0),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_205),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_39),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_45),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_5),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_185),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_26),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_19),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_58),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_1),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_23),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_53),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_158),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_35),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_120),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_48),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_80),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_103),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_99),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_111),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_155),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_68),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_46),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_153),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_117),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_69),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_71),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_126),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_10),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_199),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_52),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_73),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_1),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_61),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_22),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_198),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_26),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_67),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_112),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_75),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_50),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_31),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_41),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_136),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_64),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_178),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_41),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_9),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_108),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_181),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_156),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_164),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_67),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_70),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_128),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_42),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_46),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_43),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_57),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_10),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_192),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_151),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_186),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_54),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_124),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_75),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_43),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_29),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_3),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_163),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_18),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_48),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_105),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_322),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_211),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_254),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_336),
.B(n_2),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_216),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_250),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_324),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_R g425 ( 
.A(n_218),
.B(n_2),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_5),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_316),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_6),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_221),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_222),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_353),
.B(n_6),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_347),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_316),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_226),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_R g437 ( 
.A(n_227),
.B(n_7),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_217),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_316),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_316),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_316),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_316),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_338),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_316),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_233),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_343),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_373),
.B(n_7),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_361),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_8),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_389),
.B(n_8),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_394),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_344),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_389),
.B(n_11),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_242),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_244),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_217),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_214),
.B(n_12),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_344),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_245),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_224),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_353),
.B(n_13),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_247),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_248),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_214),
.B(n_13),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_307),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_344),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_300),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_213),
.B(n_14),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_249),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_252),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_396),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_235),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_235),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_304),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_256),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_258),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_261),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_268),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_220),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_215),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_220),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_272),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_273),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_238),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_R g493 ( 
.A(n_275),
.B(n_140),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_238),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_307),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_276),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_257),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_257),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_259),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_280),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_231),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_281),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_232),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_259),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_286),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_289),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_293),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_260),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_260),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_297),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_301),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_303),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_312),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_313),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_262),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_262),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_314),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_318),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_319),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_325),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_334),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_282),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_469),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_421),
.B(n_291),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_445),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_427),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_429),
.A2(n_263),
.B(n_239),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_506),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_449),
.B(n_228),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_423),
.B(n_212),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_429),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_506),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_468),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_468),
.B(n_239),
.Y(n_544)
);

OA21x2_ASAP7_75t_L g545 ( 
.A1(n_472),
.A2(n_290),
.B(n_282),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_417),
.B(n_304),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_472),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_432),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_473),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_473),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_426),
.B(n_291),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_475),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_435),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_419),
.A2(n_234),
.B1(n_328),
.B2(n_269),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_475),
.B(n_263),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_495),
.B(n_213),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_476),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_477),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_477),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_435),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_506),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_489),
.Y(n_568)
);

BUFx8_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_506),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_489),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_418),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_439),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_428),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_439),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_440),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_467),
.B(n_219),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_440),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_451),
.B(n_308),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_492),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_506),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_492),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_511),
.B(n_441),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_441),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_494),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

AND3x2_ASAP7_75t_L g588 ( 
.A(n_452),
.B(n_287),
.C(n_265),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_497),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_497),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_433),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_498),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_453),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_498),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_422),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_442),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_442),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_444),
.B(n_265),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_499),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_444),
.B(n_287),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_478),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_459),
.A2(n_323),
.B(n_295),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_504),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_504),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_511),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_478),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_455),
.B(n_360),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_509),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_585),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_579),
.A2(n_527),
.B1(n_537),
.B2(n_609),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_572),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_536),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_531),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_537),
.B(n_430),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_531),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_597),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_531),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_585),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_531),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_574),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_538),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_536),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_609),
.B(n_431),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_579),
.A2(n_470),
.B1(n_466),
.B2(n_290),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_536),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_597),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_534),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_527),
.B(n_436),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_607),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_546),
.B(n_595),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_585),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_534),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_534),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_534),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_607),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_479),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_574),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_559),
.A2(n_292),
.B1(n_306),
.B2(n_294),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_559),
.B(n_583),
.C(n_545),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_539),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_597),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_525),
.B(n_462),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_607),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_536),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_559),
.A2(n_292),
.B1(n_306),
.B2(n_294),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_539),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_539),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_583),
.A2(n_309),
.B1(n_337),
.B2(n_329),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_598),
.B(n_295),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_547),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_607),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_539),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_545),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_577),
.B(n_219),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_549),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_526),
.B(n_446),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_536),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_526),
.B(n_503),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_591),
.B(n_456),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_597),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_549),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_591),
.B(n_457),
.Y(n_666)
);

AO22x2_ASAP7_75t_L g667 ( 
.A1(n_552),
.A2(n_329),
.B1(n_337),
.B2(n_309),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_549),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_553),
.Y(n_669)
);

AND2x6_ASAP7_75t_L g670 ( 
.A(n_598),
.B(n_323),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_553),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_553),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_SL g673 ( 
.A1(n_552),
.A2(n_225),
.B1(n_229),
.B2(n_223),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_577),
.B(n_479),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_604),
.B(n_461),
.Y(n_675)
);

CKINVDCx11_ASAP7_75t_R g676 ( 
.A(n_525),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_553),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_604),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_555),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_555),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_555),
.Y(n_681)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_538),
.B(n_424),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_555),
.Y(n_683)
);

CKINVDCx6p67_ASAP7_75t_R g684 ( 
.A(n_547),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_588),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_536),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_588),
.B(n_465),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_577),
.B(n_471),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_565),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_565),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_557),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_565),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_573),
.Y(n_695)
);

BUFx4f_ASAP7_75t_L g696 ( 
.A(n_545),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_603),
.B(n_223),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_536),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_573),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_541),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_573),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

NOR2x1_ASAP7_75t_L g703 ( 
.A(n_545),
.B(n_284),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_557),
.B(n_474),
.Y(n_705)
);

INVx6_ASAP7_75t_L g706 ( 
.A(n_569),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_541),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_481),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_569),
.B(n_483),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_541),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_575),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_575),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_569),
.B(n_490),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_547),
.B(n_496),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_545),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_576),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_598),
.A2(n_340),
.B1(n_355),
.B2(n_345),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_545),
.B(n_438),
.C(n_229),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_569),
.B(n_502),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_587),
.B(n_507),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_576),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_576),
.Y(n_722)
);

AND2x6_ASAP7_75t_L g723 ( 
.A(n_598),
.B(n_362),
.Y(n_723)
);

NOR2x1p5_ASAP7_75t_L g724 ( 
.A(n_564),
.B(n_340),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_538),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_576),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_569),
.B(n_508),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_525),
.A2(n_484),
.B1(n_485),
.B2(n_464),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_597),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_578),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_564),
.B(n_482),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_578),
.B(n_512),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_546),
.B(n_515),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_587),
.B(n_516),
.Y(n_734)
);

INVx5_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_587),
.B(n_519),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_556),
.B(n_521),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_578),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_578),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_556),
.B(n_522),
.Y(n_740)
);

INVx5_ASAP7_75t_L g741 ( 
.A(n_597),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_596),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_566),
.B(n_482),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_566),
.B(n_568),
.Y(n_744)
);

INVx5_ASAP7_75t_L g745 ( 
.A(n_597),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_598),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_568),
.B(n_523),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_596),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_596),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_600),
.B(n_480),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_600),
.B(n_480),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_593),
.B(n_376),
.C(n_230),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_571),
.B(n_458),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_596),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_567),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_541),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_528),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_600),
.B(n_366),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_528),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_600),
.B(n_362),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_674),
.B(n_571),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_684),
.B(n_236),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_640),
.B(n_580),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_759),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_612),
.B(n_600),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_616),
.B(n_661),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_708),
.B(n_544),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_732),
.B(n_544),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_747),
.B(n_544),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_666),
.B(n_640),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_582),
.B(n_584),
.C(n_580),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_630),
.A2(n_500),
.B1(n_505),
.B2(n_491),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_759),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_705),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_639),
.B(n_544),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_639),
.B(n_744),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_744),
.B(n_558),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_696),
.B(n_642),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_656),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_746),
.B(n_558),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_678),
.B(n_513),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_746),
.B(n_558),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_631),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_731),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_611),
.B(n_558),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_678),
.B(n_514),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_731),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_693),
.B(n_593),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_642),
.A2(n_603),
.B1(n_558),
.B2(n_237),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_631),
.B(n_582),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_656),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_757),
.Y(n_792)
);

BUFx8_ASAP7_75t_L g793 ( 
.A(n_645),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_715),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_611),
.B(n_529),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_757),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_620),
.B(n_529),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_743),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_620),
.B(n_530),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_743),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_689),
.B(n_520),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_696),
.B(n_715),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_696),
.B(n_395),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_626),
.A2(n_603),
.B1(n_237),
.B2(n_241),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_659),
.B(n_443),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_646),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_703),
.B(n_395),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_703),
.B(n_395),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_718),
.A2(n_241),
.B1(n_253),
.B2(n_225),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_652),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_615),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_614),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_674),
.B(n_584),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_633),
.B(n_532),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_638),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_638),
.B(n_533),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_637),
.B(n_533),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_693),
.B(n_593),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_615),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_617),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_675),
.B(n_447),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_617),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_737),
.B(n_450),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_622),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_657),
.B(n_540),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_753),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_654),
.B(n_586),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_625),
.A2(n_437),
.B1(n_425),
.B2(n_387),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_753),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_619),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_645),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_755),
.B(n_542),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_654),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_667),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_652),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_758),
.B(n_542),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_740),
.B(n_385),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_632),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_619),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_621),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_724),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_650),
.B(n_543),
.Y(n_843)
);

INVx8_ASAP7_75t_L g844 ( 
.A(n_652),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_650),
.B(n_543),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_685),
.B(n_240),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_665),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_685),
.B(n_243),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_750),
.B(n_246),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_751),
.B(n_251),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_718),
.A2(n_379),
.B1(n_253),
.B2(n_267),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_613),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_669),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_669),
.B(n_548),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_671),
.B(n_672),
.Y(n_856)
);

INVxp33_ASAP7_75t_L g857 ( 
.A(n_720),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_621),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_614),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_671),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_673),
.A2(n_610),
.B(n_606),
.C(n_605),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_688),
.B(n_395),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_623),
.B(n_725),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_672),
.B(n_550),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_629),
.B(n_370),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_736),
.B(n_255),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_677),
.B(n_550),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_663),
.A2(n_713),
.B1(n_719),
.B2(n_709),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_677),
.B(n_551),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_728),
.B(n_733),
.C(n_752),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_706),
.A2(n_393),
.B1(n_267),
.B2(n_277),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_679),
.B(n_551),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_652),
.A2(n_264),
.B1(n_382),
.B2(n_277),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_634),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_667),
.B(n_586),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_679),
.B(n_554),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_734),
.B(n_266),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_635),
.B(n_398),
.Y(n_878)
);

AOI22x1_ASAP7_75t_L g879 ( 
.A1(n_667),
.A2(n_363),
.B1(n_367),
.B2(n_296),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_641),
.A2(n_590),
.B(n_592),
.C(n_589),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_667),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_614),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_635),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_680),
.B(n_554),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_653),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_613),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_636),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_680),
.B(n_560),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_636),
.B(n_404),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_683),
.B(n_560),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_697),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_643),
.Y(n_892)
);

BUFx8_ASAP7_75t_L g893 ( 
.A(n_684),
.Y(n_893)
);

OAI22xp33_ASAP7_75t_L g894 ( 
.A1(n_706),
.A2(n_330),
.B1(n_326),
.B2(n_317),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_643),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_683),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_727),
.B(n_589),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_649),
.B(n_406),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_653),
.B(n_509),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_687),
.B(n_561),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_613),
.B(n_270),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_687),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_649),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_655),
.B(n_408),
.Y(n_904)
);

BUFx6f_ASAP7_75t_SL g905 ( 
.A(n_613),
.Y(n_905)
);

AND2x4_ASAP7_75t_SL g906 ( 
.A(n_648),
.B(n_291),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_690),
.B(n_561),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_682),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_655),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_697),
.B(n_590),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_697),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_SL g912 ( 
.A(n_706),
.B(n_541),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_676),
.B(n_274),
.C(n_271),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_658),
.B(n_413),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_692),
.B(n_562),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_682),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_806),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_766),
.A2(n_765),
.B(n_881),
.C(n_776),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_767),
.A2(n_768),
.B(n_803),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_779),
.B(n_644),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_853),
.B(n_886),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_774),
.B(n_341),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_770),
.B(n_694),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_769),
.B(n_694),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_857),
.B(n_356),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_764),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_838),
.A2(n_717),
.B(n_651),
.C(n_535),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_803),
.A2(n_628),
.B(n_644),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_778),
.A2(n_706),
.B1(n_697),
.B2(n_279),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_802),
.A2(n_697),
.B(n_695),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_777),
.A2(n_729),
.B(n_664),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_857),
.B(n_664),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_788),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_863),
.B(n_592),
.Y(n_934)
);

BUFx12f_ASAP7_75t_L g935 ( 
.A(n_893),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_792),
.B(n_695),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_792),
.B(n_796),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_779),
.B(n_791),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_779),
.B(n_664),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_796),
.B(n_701),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_866),
.B(n_701),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_802),
.A2(n_729),
.B(n_624),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_852),
.B(n_729),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_827),
.B(n_594),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_791),
.B(n_614),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_775),
.A2(n_624),
.B(n_614),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_816),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_761),
.B(n_702),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_807),
.A2(n_704),
.B(n_702),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_893),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_839),
.B(n_704),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_806),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_881),
.A2(n_862),
.B(n_875),
.C(n_771),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_836),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_L g955 ( 
.A(n_781),
.B(n_786),
.C(n_801),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_780),
.A2(n_686),
.B(n_624),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_849),
.A2(n_850),
.B(n_906),
.C(n_877),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_761),
.B(n_712),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_782),
.A2(n_686),
.B(n_624),
.Y(n_959)
);

O2A1O1Ixp5_ASAP7_75t_L g960 ( 
.A1(n_862),
.A2(n_662),
.B(n_668),
.C(n_658),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_814),
.B(n_712),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_794),
.B(n_624),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_807),
.A2(n_721),
.B(n_716),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_844),
.A2(n_691),
.B(n_686),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_788),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_L g966 ( 
.A1(n_824),
.A2(n_279),
.B(n_264),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_814),
.B(n_716),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_794),
.B(n_810),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_790),
.B(n_721),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_830),
.B(n_730),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_790),
.B(n_730),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_819),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_853),
.B(n_652),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_810),
.B(n_686),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_819),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_790),
.B(n_739),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_828),
.B(n_739),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_828),
.B(n_742),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_875),
.A2(n_742),
.B(n_748),
.C(n_754),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_764),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_828),
.B(n_748),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_844),
.A2(n_691),
.B(n_686),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_891),
.A2(n_371),
.B1(n_393),
.B2(n_392),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_910),
.A2(n_760),
.B1(n_670),
.B2(n_723),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_784),
.B(n_754),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_844),
.A2(n_710),
.B(n_691),
.Y(n_986)
);

OAI21xp33_ASAP7_75t_L g987 ( 
.A1(n_846),
.A2(n_298),
.B(n_278),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_910),
.A2(n_760),
.B1(n_670),
.B2(n_652),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_808),
.A2(n_789),
.B(n_804),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_836),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_787),
.B(n_681),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_899),
.B(n_594),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_910),
.A2(n_288),
.B(n_285),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_810),
.A2(n_710),
.B(n_691),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_798),
.B(n_699),
.Y(n_995)
);

OAI21xp33_ASAP7_75t_L g996 ( 
.A1(n_848),
.A2(n_302),
.B(n_299),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_891),
.A2(n_367),
.B1(n_392),
.B2(n_382),
.Y(n_997)
);

OAI321xp33_ASAP7_75t_L g998 ( 
.A1(n_868),
.A2(n_374),
.A3(n_345),
.B1(n_377),
.B2(n_368),
.C(n_365),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_785),
.A2(n_711),
.B(n_699),
.Y(n_999)
);

AO22x1_ASAP7_75t_L g1000 ( 
.A1(n_870),
.A2(n_346),
.B1(n_310),
.B2(n_414),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_906),
.A2(n_357),
.B(n_371),
.C(n_285),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_911),
.A2(n_357),
.B1(n_379),
.B2(n_288),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_899),
.B(n_711),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_783),
.B(n_599),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_831),
.A2(n_710),
.B(n_618),
.Y(n_1005)
);

AOI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_901),
.A2(n_305),
.B(n_296),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_800),
.B(n_722),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_806),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_863),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_836),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_879),
.A2(n_760),
.B1(n_652),
.B2(n_670),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_837),
.A2(n_710),
.B(n_618),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_763),
.B(n_722),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_818),
.B(n_726),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_773),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_L g1016 ( 
.A(n_836),
.B(n_670),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_911),
.B(n_627),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_861),
.A2(n_738),
.B(n_749),
.C(n_333),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_783),
.B(n_305),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_825),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_836),
.B(n_627),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_832),
.B(n_738),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_806),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_834),
.B(n_749),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_773),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_809),
.B(n_647),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_851),
.A2(n_333),
.B1(n_405),
.B2(n_330),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_886),
.B(n_599),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_826),
.B(n_647),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_835),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_806),
.B(n_647),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_833),
.A2(n_735),
.B(n_618),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_885),
.B(n_602),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_856),
.A2(n_741),
.B(n_735),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_847),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_835),
.B(n_660),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_854),
.A2(n_698),
.B(n_660),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_842),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_860),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_805),
.B(n_698),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_812),
.B(n_698),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_813),
.A2(n_741),
.B(n_735),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_812),
.B(n_700),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_813),
.A2(n_745),
.B(n_741),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_865),
.A2(n_700),
.B(n_756),
.C(n_707),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_896),
.B(n_700),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_813),
.A2(n_882),
.B(n_859),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_902),
.B(n_707),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_811),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_820),
.B(n_707),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_880),
.A2(n_405),
.B(n_311),
.C(n_317),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_897),
.A2(n_760),
.B1(n_723),
.B2(n_670),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_829),
.B(n_756),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_820),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_821),
.B(n_756),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_859),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_859),
.A2(n_882),
.B(n_797),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_772),
.Y(n_1058)
);

AO21x1_ASAP7_75t_L g1059 ( 
.A1(n_894),
.A2(n_326),
.B(n_311),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_762),
.B(n_602),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_882),
.A2(n_745),
.B(n_741),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_821),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_793),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_823),
.B(n_741),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_793),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_905),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_823),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_840),
.B(n_670),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_793),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_893),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_795),
.A2(n_745),
.B(n_741),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_799),
.A2(n_745),
.B(n_581),
.Y(n_1072)
);

AOI33xp33_ASAP7_75t_L g1073 ( 
.A1(n_873),
.A2(n_411),
.A3(n_384),
.B1(n_374),
.B2(n_368),
.B3(n_365),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_840),
.B(n_670),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_841),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_815),
.A2(n_581),
.B(n_541),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_817),
.A2(n_581),
.B(n_567),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_822),
.A2(n_384),
.B(n_415),
.C(n_355),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_865),
.A2(n_889),
.B(n_878),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_841),
.A2(n_399),
.B(n_377),
.C(n_409),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_858),
.B(n_723),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_858),
.A2(n_760),
.B(n_723),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_889),
.A2(n_363),
.B(n_354),
.C(n_610),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_898),
.A2(n_354),
.B(n_606),
.C(n_605),
.Y(n_1084)
);

AO21x1_ASAP7_75t_L g1085 ( 
.A1(n_871),
.A2(n_403),
.B(n_409),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_913),
.B(n_510),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_898),
.A2(n_562),
.B(n_563),
.C(n_352),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_908),
.B(n_304),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_919),
.A2(n_912),
.B(n_845),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1009),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1003),
.B(n_874),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1035),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_934),
.B(n_916),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_954),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_957),
.A2(n_904),
.B(n_914),
.C(n_887),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_SL g1096 ( 
.A(n_973),
.B(n_905),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1058),
.A2(n_879),
.B1(n_914),
.B2(n_905),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_989),
.A2(n_883),
.B1(n_909),
.B2(n_887),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_922),
.B(n_883),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_935),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_925),
.B(n_320),
.C(n_315),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_966),
.A2(n_892),
.B(n_909),
.C(n_895),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1039),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_937),
.B(n_892),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_965),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_922),
.B(n_895),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_954),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1003),
.B(n_903),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1062),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_939),
.A2(n_915),
.B(n_907),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_925),
.B(n_972),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1016),
.A2(n_869),
.B(n_900),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_968),
.A2(n_867),
.B(n_890),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1062),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_968),
.A2(n_855),
.B(n_888),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1006),
.A2(n_903),
.B(n_884),
.C(n_876),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1063),
.A2(n_383),
.B1(n_321),
.B2(n_327),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1020),
.B(n_872),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1069),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_927),
.A2(n_864),
.B1(n_843),
.B2(n_359),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_955),
.A2(n_283),
.B(n_349),
.C(n_359),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_927),
.A2(n_399),
.B1(n_403),
.B2(n_411),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1067),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1004),
.B(n_1038),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_947),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_954),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_924),
.A2(n_974),
.B(n_920),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1040),
.A2(n_932),
.B1(n_992),
.B2(n_933),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_965),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_933),
.B(n_493),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_975),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1028),
.B(n_291),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_923),
.B(n_723),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1056),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1030),
.A2(n_760),
.B1(n_723),
.B2(n_304),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_950),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1056),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_948),
.A2(n_390),
.B1(n_332),
.B2(n_335),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_1065),
.B(n_517),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1004),
.B(n_331),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_975),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1030),
.A2(n_723),
.B1(n_760),
.B2(n_563),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1049),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_942),
.A2(n_570),
.B(n_601),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1022),
.B(n_339),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1040),
.A2(n_601),
.B1(n_388),
.B2(n_386),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_921),
.A2(n_342),
.B1(n_350),
.B2(n_351),
.Y(n_1147)
);

BUFx8_ASAP7_75t_SL g1148 ( 
.A(n_1070),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1033),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1054),
.Y(n_1150)
);

INVx6_ASAP7_75t_L g1151 ( 
.A(n_1066),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_926),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1022),
.B(n_358),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1078),
.A2(n_524),
.B(n_518),
.C(n_517),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_980),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1015),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_932),
.A2(n_951),
.B1(n_1086),
.B2(n_1038),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_944),
.Y(n_1158)
);

BUFx2_ASAP7_75t_SL g1159 ( 
.A(n_1066),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_954),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_951),
.B(n_601),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_1088),
.B(n_364),
.Y(n_1162)
);

AND2x6_ASAP7_75t_L g1163 ( 
.A(n_990),
.B(n_1010),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1056),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_920),
.A2(n_608),
.B(n_518),
.Y(n_1165)
);

BUFx5_ASAP7_75t_L g1166 ( 
.A(n_1060),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_958),
.B(n_608),
.Y(n_1167)
);

BUFx4f_ASAP7_75t_L g1168 ( 
.A(n_1060),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1000),
.B(n_486),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_970),
.B(n_608),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_994),
.A2(n_608),
.B(n_486),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_917),
.B(n_952),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_973),
.B(n_369),
.Y(n_1173)
);

OA22x2_ASAP7_75t_L g1174 ( 
.A1(n_1086),
.A2(n_412),
.B1(n_410),
.B2(n_407),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_SL g1175 ( 
.A1(n_1053),
.A2(n_193),
.B(n_188),
.C(n_183),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1025),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_990),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1056),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1036),
.A2(n_608),
.B1(n_401),
.B2(n_400),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1075),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_928),
.A2(n_608),
.B(n_154),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1075),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_990),
.B(n_608),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_961),
.B(n_372),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1075),
.Y(n_1185)
);

BUFx8_ASAP7_75t_SL g1186 ( 
.A(n_990),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_987),
.B(n_375),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1036),
.A2(n_391),
.B1(n_381),
.B2(n_380),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_938),
.A2(n_138),
.B(n_97),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_996),
.B(n_397),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_SL g1191 ( 
.A(n_1019),
.B(n_378),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_943),
.B(n_15),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_943),
.B(n_176),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1001),
.A2(n_18),
.B(n_21),
.C(n_23),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_L g1195 ( 
.A(n_998),
.B(n_1027),
.C(n_918),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1010),
.Y(n_1196)
);

INVx3_ASAP7_75t_SL g1197 ( 
.A(n_917),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_991),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_941),
.B(n_24),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_970),
.A2(n_169),
.B(n_165),
.C(n_157),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_967),
.B(n_150),
.Y(n_1201)
);

AO22x1_ASAP7_75t_L g1202 ( 
.A1(n_1023),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_985),
.B(n_146),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1011),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1011),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_936),
.B(n_135),
.Y(n_1206)
);

NOR3xp33_ASAP7_75t_SL g1207 ( 
.A(n_1080),
.B(n_36),
.C(n_38),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1014),
.B(n_39),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_995),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1010),
.B(n_134),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_984),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1075),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_952),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_969),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1010),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_938),
.A2(n_132),
.B(n_127),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1079),
.B(n_116),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1007),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_940),
.B(n_113),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1008),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1008),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_931),
.A2(n_104),
.B(n_101),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1024),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_953),
.A2(n_40),
.B(n_49),
.C(n_51),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_971),
.B(n_49),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_976),
.B(n_93),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_988),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_977),
.B(n_56),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_SL g1229 ( 
.A(n_993),
.B(n_83),
.C(n_58),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_978),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_983),
.A2(n_57),
.B(n_62),
.C(n_63),
.Y(n_1231)
);

AOI221xp5_ASAP7_75t_L g1232 ( 
.A1(n_997),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.C(n_66),
.Y(n_1232)
);

O2A1O1Ixp5_ASAP7_75t_L g1233 ( 
.A1(n_929),
.A2(n_65),
.B(n_68),
.C(n_72),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_981),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_946),
.A2(n_80),
.B(n_77),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_SL g1236 ( 
.A(n_930),
.B(n_76),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1002),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.C(n_1051),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1017),
.A2(n_78),
.B1(n_79),
.B2(n_1021),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_R g1239 ( 
.A(n_949),
.B(n_1041),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_964),
.A2(n_982),
.B(n_986),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1029),
.B(n_979),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1018),
.A2(n_1084),
.B(n_1045),
.C(n_1083),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1050),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1013),
.B(n_1052),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1145),
.B(n_1073),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1153),
.B(n_1087),
.C(n_1080),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1122),
.A2(n_1120),
.A3(n_1095),
.B(n_1242),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1199),
.A2(n_1121),
.B1(n_1122),
.B2(n_1111),
.C(n_1138),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1148),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_1059),
.A3(n_1085),
.B(n_1057),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1092),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1196),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1198),
.B(n_1043),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1149),
.B(n_1017),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1098),
.A2(n_956),
.A3(n_959),
.B(n_1012),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1186),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1103),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_1151),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1100),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1158),
.B(n_1031),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1112),
.A2(n_1082),
.B(n_1037),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1215),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1209),
.B(n_1055),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1144),
.A2(n_960),
.B(n_1047),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1127),
.A2(n_999),
.B(n_963),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1218),
.B(n_1046),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1093),
.B(n_1021),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1134),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1098),
.A2(n_1076),
.A3(n_1026),
.B(n_1077),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1125),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1224),
.A2(n_1211),
.B(n_1227),
.C(n_1187),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1230),
.B(n_1214),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1102),
.A2(n_1116),
.A3(n_1110),
.B(n_1241),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1192),
.A2(n_1081),
.B(n_1074),
.C(n_1068),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1244),
.A2(n_1005),
.B(n_962),
.Y(n_1275)
);

AOI31xp67_ASAP7_75t_L g1276 ( 
.A1(n_1217),
.A2(n_945),
.A3(n_962),
.B(n_1064),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1157),
.B(n_1048),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1118),
.B(n_1031),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1124),
.B(n_945),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1241),
.A2(n_1072),
.A3(n_1032),
.B(n_1034),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1131),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1136),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1151),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_1163),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1113),
.A2(n_1071),
.B(n_1064),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1123),
.Y(n_1286)
);

AO32x2_ASAP7_75t_L g1287 ( 
.A1(n_1211),
.A2(n_1042),
.A3(n_1044),
.B1(n_1061),
.B2(n_1227),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1141),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_SL g1289 ( 
.A1(n_1204),
.A2(n_1205),
.B(n_1235),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1143),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1115),
.A2(n_1133),
.B(n_1219),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1150),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1152),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1196),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1133),
.A2(n_1195),
.B(n_1128),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1181),
.A2(n_1167),
.B(n_1171),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1160),
.B(n_1099),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1155),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1167),
.A2(n_1165),
.B(n_1222),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1239),
.A2(n_1170),
.B(n_1161),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1206),
.A2(n_1219),
.B(n_1091),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_SL g1302 ( 
.A(n_1101),
.B(n_1124),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1206),
.A2(n_1108),
.B(n_1203),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_SL g1304 ( 
.A1(n_1204),
.A2(n_1205),
.B(n_1194),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1226),
.A2(n_1201),
.B(n_1104),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1184),
.B(n_1105),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1231),
.A2(n_1132),
.B(n_1236),
.C(n_1229),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1156),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1200),
.A2(n_1210),
.B(n_1193),
.C(n_1097),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1106),
.A2(n_1208),
.B(n_1226),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1104),
.A2(n_1160),
.B(n_1223),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1243),
.A2(n_1189),
.B(n_1216),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1169),
.A2(n_1162),
.B(n_1184),
.C(n_1233),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1160),
.A2(n_1142),
.B(n_1183),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1176),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1238),
.A2(n_1228),
.B(n_1225),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1180),
.A2(n_1185),
.B(n_1182),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1109),
.B(n_1114),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1160),
.A2(n_1183),
.B(n_1096),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1151),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1212),
.A2(n_1094),
.B(n_1107),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1090),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1183),
.A2(n_1175),
.B(n_1135),
.Y(n_1323)
);

INVx3_ASAP7_75t_SL g1324 ( 
.A(n_1139),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1168),
.B(n_1188),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1159),
.B(n_1119),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1129),
.B(n_1140),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1138),
.B(n_1190),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1139),
.Y(n_1329)
);

CKINVDCx6p67_ASAP7_75t_R g1330 ( 
.A(n_1139),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1163),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1173),
.A2(n_1130),
.B(n_1107),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1174),
.A2(n_1237),
.B1(n_1168),
.B2(n_1147),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_SL g1334 ( 
.A(n_1163),
.B(n_1166),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1166),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1213),
.B(n_1221),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1134),
.B(n_1137),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1094),
.A2(n_1126),
.B(n_1177),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1166),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1220),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1154),
.A2(n_1174),
.B(n_1146),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1163),
.A2(n_1134),
.B(n_1137),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_1164),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1166),
.B(n_1164),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1164),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1178),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1166),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1178),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1166),
.B(n_1179),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1178),
.Y(n_1350)
);

AO21x1_ASAP7_75t_L g1351 ( 
.A1(n_1234),
.A2(n_1191),
.B(n_1202),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1232),
.A2(n_1172),
.B(n_1197),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1117),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1207),
.A2(n_1240),
.B(n_1144),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1122),
.A2(n_1120),
.A3(n_1095),
.B(n_1242),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1148),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1240),
.A2(n_1144),
.B(n_1089),
.Y(n_1357)
);

CKINVDCx8_ASAP7_75t_R g1358 ( 
.A(n_1159),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1093),
.B(n_863),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1240),
.A2(n_1144),
.B(n_1089),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1186),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1092),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1145),
.B(n_766),
.C(n_955),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1198),
.B(n_1209),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1121),
.A2(n_612),
.B(n_766),
.C(n_957),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1148),
.Y(n_1367)
);

NAND2x1p5_ASAP7_75t_L g1368 ( 
.A(n_1160),
.B(n_1168),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1127),
.A2(n_919),
.B(n_957),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1100),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1095),
.A2(n_919),
.B(n_1242),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1121),
.A2(n_612),
.B(n_766),
.C(n_957),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1131),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1196),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_SL g1375 ( 
.A(n_1159),
.B(n_935),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1121),
.A2(n_612),
.B(n_766),
.C(n_957),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1093),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1122),
.A2(n_1120),
.A3(n_1095),
.B(n_1242),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1090),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_SL g1381 ( 
.A1(n_1224),
.A2(n_957),
.B(n_966),
.C(n_1006),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1240),
.A2(n_1144),
.B(n_1089),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1122),
.A2(n_1120),
.A3(n_1095),
.B(n_1242),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1131),
.Y(n_1385)
);

AO32x2_ASAP7_75t_L g1386 ( 
.A1(n_1122),
.A2(n_1120),
.A3(n_1227),
.B1(n_1211),
.B2(n_1204),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1198),
.B(n_1209),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1149),
.B(n_1158),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1186),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1100),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1198),
.B(n_1209),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1186),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1198),
.B(n_1209),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1145),
.B(n_766),
.C(n_955),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1122),
.A2(n_1120),
.A3(n_1095),
.B(n_1242),
.Y(n_1397)
);

BUFx8_ASAP7_75t_L g1398 ( 
.A(n_1131),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1240),
.A2(n_1144),
.B(n_1089),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1093),
.B(n_863),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1198),
.B(n_1209),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1240),
.A2(n_1144),
.B(n_1089),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1199),
.A2(n_766),
.B(n_957),
.C(n_955),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1236),
.A2(n_766),
.B1(n_612),
.B2(n_955),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1089),
.A2(n_919),
.B(n_957),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1273),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1388),
.B(n_1254),
.Y(n_1411)
);

INVx3_ASAP7_75t_SL g1412 ( 
.A(n_1367),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1408),
.A2(n_1364),
.B1(n_1396),
.B2(n_1407),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1362),
.A2(n_1383),
.B(n_1380),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1284),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1258),
.Y(n_1416)
);

CKINVDCx11_ASAP7_75t_R g1417 ( 
.A(n_1249),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1356),
.Y(n_1418)
);

INVx2_ASAP7_75t_R g1419 ( 
.A(n_1284),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1251),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1284),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1398),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1365),
.B(n_1387),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1257),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1398),
.Y(n_1425)
);

BUFx8_ASAP7_75t_SL g1426 ( 
.A(n_1370),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1283),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1304),
.B2(n_1353),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1408),
.A2(n_1248),
.B1(n_1339),
.B2(n_1328),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1351),
.A2(n_1316),
.B1(n_1289),
.B2(n_1333),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1273),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1320),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1281),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1288),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1373),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1256),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1365),
.A2(n_1392),
.B1(n_1387),
.B2(n_1395),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1392),
.A2(n_1395),
.B1(n_1403),
.B2(n_1377),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1282),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1359),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1316),
.A2(n_1245),
.B1(n_1246),
.B2(n_1310),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1403),
.A2(n_1306),
.B1(n_1353),
.B2(n_1272),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1325),
.A2(n_1246),
.B1(n_1278),
.B2(n_1327),
.Y(n_1443)
);

INVx6_ASAP7_75t_L g1444 ( 
.A(n_1258),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1270),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1363),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1259),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1345),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1260),
.B(n_1267),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1290),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1292),
.Y(n_1451)
);

INVx4_ASAP7_75t_L g1452 ( 
.A(n_1331),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_SL g1453 ( 
.A(n_1358),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1310),
.A2(n_1295),
.B1(n_1277),
.B2(n_1302),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1272),
.B(n_1253),
.Y(n_1455)
);

INVx4_ASAP7_75t_L g1456 ( 
.A(n_1331),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1253),
.B(n_1402),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1295),
.A2(n_1341),
.B1(n_1298),
.B2(n_1293),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1271),
.A2(n_1329),
.B1(n_1366),
.B2(n_1372),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1308),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1315),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1317),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1266),
.A2(n_1369),
.B1(n_1371),
.B2(n_1279),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1268),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1376),
.A2(n_1307),
.B(n_1313),
.Y(n_1465)
);

BUFx2_ASAP7_75t_SL g1466 ( 
.A(n_1256),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1352),
.A2(n_1322),
.B1(n_1379),
.B2(n_1330),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1369),
.A2(n_1371),
.B1(n_1279),
.B2(n_1303),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1361),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1385),
.A2(n_1324),
.B1(n_1297),
.B2(n_1326),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1394),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1297),
.A2(n_1326),
.B1(n_1314),
.B2(n_1263),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1391),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_1256),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1390),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1390),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1368),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1301),
.A2(n_1263),
.B1(n_1286),
.B2(n_1349),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1318),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1336),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1334),
.A2(n_1390),
.B1(n_1386),
.B2(n_1323),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1336),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1326),
.Y(n_1483)
);

INVx5_ASAP7_75t_L g1484 ( 
.A(n_1268),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1340),
.B(n_1348),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1321),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1350),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1337),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1262),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1262),
.Y(n_1490)
);

BUFx2_ASAP7_75t_SL g1491 ( 
.A(n_1262),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1344),
.A2(n_1346),
.B1(n_1347),
.B2(n_1335),
.Y(n_1492)
);

CKINVDCx6p67_ASAP7_75t_R g1493 ( 
.A(n_1268),
.Y(n_1493)
);

OAI21xp33_ASAP7_75t_L g1494 ( 
.A1(n_1332),
.A2(n_1311),
.B(n_1375),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1338),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1344),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1265),
.A2(n_1386),
.B1(n_1406),
.B2(n_1405),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1346),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1337),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1265),
.A2(n_1386),
.B1(n_1409),
.B2(n_1401),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1389),
.A2(n_1393),
.B1(n_1399),
.B2(n_1300),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1300),
.A2(n_1305),
.B1(n_1261),
.B2(n_1381),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1252),
.B(n_1294),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1274),
.A2(n_1291),
.B(n_1275),
.Y(n_1504)
);

CKINVDCx9p33_ASAP7_75t_R g1505 ( 
.A(n_1334),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1294),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1285),
.A2(n_1354),
.B1(n_1312),
.B2(n_1374),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1319),
.A2(n_1397),
.B1(n_1247),
.B2(n_1378),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1342),
.Y(n_1509)
);

CKINVDCx6p67_ASAP7_75t_R g1510 ( 
.A(n_1343),
.Y(n_1510)
);

BUFx10_ASAP7_75t_L g1511 ( 
.A(n_1309),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1247),
.A2(n_1378),
.B1(n_1355),
.B2(n_1397),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1287),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1285),
.A2(n_1247),
.B1(n_1384),
.B2(n_1378),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1355),
.A2(n_1384),
.B1(n_1299),
.B2(n_1296),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1357),
.A2(n_1404),
.B1(n_1400),
.B2(n_1382),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1360),
.A2(n_1264),
.B1(n_1250),
.B2(n_1287),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_SL g1518 ( 
.A1(n_1250),
.A2(n_1287),
.B(n_1276),
.Y(n_1518)
);

BUFx2_ASAP7_75t_SL g1519 ( 
.A(n_1280),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1250),
.B(n_1269),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1280),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1280),
.A2(n_955),
.B1(n_766),
.B2(n_1364),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1255),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1269),
.A2(n_1364),
.B1(n_1396),
.B2(n_1408),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1255),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1255),
.A2(n_1408),
.B1(n_1236),
.B2(n_1396),
.Y(n_1526)
);

BUFx2_ASAP7_75t_SL g1527 ( 
.A(n_1282),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1364),
.A2(n_955),
.B1(n_766),
.B2(n_1396),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1365),
.B(n_766),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1532)
);

CKINVDCx11_ASAP7_75t_R g1533 ( 
.A(n_1249),
.Y(n_1533)
);

INVx8_ASAP7_75t_L g1534 ( 
.A(n_1283),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1362),
.A2(n_1383),
.B(n_1380),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1365),
.B(n_766),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1256),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1258),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1541)
);

BUFx10_ASAP7_75t_L g1542 ( 
.A(n_1256),
.Y(n_1542)
);

BUFx8_ASAP7_75t_SL g1543 ( 
.A(n_1249),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1283),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1364),
.A2(n_632),
.B1(n_1396),
.B2(n_766),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1284),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1284),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1364),
.A2(n_632),
.B1(n_1396),
.B2(n_766),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1365),
.B(n_766),
.Y(n_1549)
);

BUFx8_ASAP7_75t_SL g1550 ( 
.A(n_1249),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1364),
.A2(n_632),
.B1(n_1396),
.B2(n_766),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1408),
.A2(n_1364),
.B1(n_1396),
.B2(n_766),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1408),
.A2(n_1364),
.B1(n_1396),
.B2(n_766),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1398),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1364),
.A2(n_1396),
.B1(n_1408),
.B2(n_1248),
.Y(n_1555)
);

BUFx10_ASAP7_75t_L g1556 ( 
.A(n_1256),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1284),
.Y(n_1557)
);

BUFx8_ASAP7_75t_L g1558 ( 
.A(n_1256),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1256),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1353),
.A2(n_766),
.B1(n_682),
.B2(n_824),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1306),
.B(n_1359),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1258),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1408),
.A2(n_1236),
.B1(n_1396),
.B2(n_1364),
.Y(n_1563)
);

BUFx8_ASAP7_75t_L g1564 ( 
.A(n_1256),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1283),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1449),
.B(n_1524),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1410),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1560),
.B(n_1440),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_SL g1569 ( 
.A(n_1511),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1410),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1524),
.B(n_1496),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1414),
.A2(n_1536),
.B(n_1516),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1434),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1431),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1431),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1437),
.B(n_1423),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1521),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1455),
.B(n_1438),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1504),
.A2(n_1516),
.B(n_1501),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1529),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1495),
.B(n_1486),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1435),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1528),
.B(n_1529),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1523),
.B(n_1462),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1525),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1507),
.A2(n_1501),
.B(n_1502),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1415),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1444),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1520),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1552),
.A2(n_1553),
.B(n_1530),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1532),
.B(n_1535),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1523),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1532),
.A2(n_1539),
.B(n_1535),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1513),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1512),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1461),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1519),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1539),
.A2(n_1555),
.B(n_1541),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1421),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1420),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1424),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1561),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1411),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1444),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1512),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1505),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1541),
.B(n_1555),
.Y(n_1607)
);

AO21x2_ASAP7_75t_L g1608 ( 
.A1(n_1526),
.A2(n_1508),
.B(n_1518),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1517),
.A2(n_1468),
.B(n_1497),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1508),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1468),
.A2(n_1497),
.B(n_1500),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1433),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1500),
.A2(n_1514),
.B(n_1463),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1445),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1465),
.A2(n_1514),
.B(n_1522),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1446),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1481),
.B(n_1413),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1450),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1451),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1441),
.A2(n_1430),
.B(n_1458),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1505),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1460),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1441),
.B(n_1463),
.Y(n_1623)
);

AOI21xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1563),
.A2(n_1551),
.B(n_1548),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1479),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1430),
.A2(n_1478),
.B(n_1454),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1459),
.A2(n_1478),
.B(n_1472),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1531),
.B(n_1537),
.Y(n_1629)
);

CKINVDCx6p67_ASAP7_75t_R g1630 ( 
.A(n_1436),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1454),
.B(n_1428),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1452),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1515),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1487),
.Y(n_1634)
);

AOI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1429),
.A2(n_1470),
.B(n_1467),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1545),
.A2(n_1563),
.B(n_1526),
.Y(n_1636)
);

AOI21xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1549),
.A2(n_1442),
.B(n_1412),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1492),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1511),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1439),
.B(n_1480),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1442),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1509),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1482),
.B(n_1457),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1494),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1456),
.Y(n_1645)
);

CKINVDCx16_ASAP7_75t_R g1646 ( 
.A(n_1453),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1510),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1527),
.B(n_1412),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1485),
.B(n_1499),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1419),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1419),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1483),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1503),
.A2(n_1506),
.B(n_1488),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1456),
.A2(n_1477),
.B(n_1416),
.Y(n_1654)
);

INVx3_ASAP7_75t_SL g1655 ( 
.A(n_1444),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1546),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1546),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1477),
.A2(n_1416),
.B(n_1562),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1547),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1484),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1557),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1557),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1464),
.B(n_1484),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1425),
.A2(n_1554),
.B1(n_1422),
.B2(n_1466),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1447),
.B(n_1498),
.Y(n_1665)
);

CKINVDCx16_ASAP7_75t_R g1666 ( 
.A(n_1436),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1464),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1540),
.Y(n_1668)
);

OA21x2_ASAP7_75t_L g1669 ( 
.A1(n_1489),
.A2(n_1476),
.B(n_1493),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1538),
.A2(n_1559),
.B1(n_1490),
.B2(n_1565),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1540),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1562),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1448),
.B(n_1491),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1448),
.B(n_1565),
.Y(n_1674)
);

OR2x2_ASAP7_75t_SL g1675 ( 
.A(n_1646),
.B(n_1550),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1593),
.A2(n_1475),
.B1(n_1469),
.B2(n_1471),
.Y(n_1676)
);

AO32x2_ASAP7_75t_L g1677 ( 
.A1(n_1667),
.A2(n_1594),
.A3(n_1604),
.B1(n_1588),
.B2(n_1653),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1580),
.A2(n_1544),
.B1(n_1427),
.B2(n_1432),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1566),
.B(n_1544),
.Y(n_1679)
);

A2O1A1Ixp33_ASAP7_75t_SL g1680 ( 
.A1(n_1590),
.A2(n_1556),
.B(n_1542),
.C(n_1534),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1593),
.A2(n_1534),
.B(n_1432),
.C(n_1427),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1566),
.B(n_1556),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1602),
.B(n_1534),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1577),
.B(n_1542),
.Y(n_1684)
);

AND2x4_ASAP7_75t_SL g1685 ( 
.A(n_1612),
.B(n_1564),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1624),
.A2(n_1564),
.B(n_1558),
.C(n_1474),
.Y(n_1686)
);

A2O1A1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1598),
.A2(n_1558),
.B(n_1474),
.C(n_1559),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1624),
.A2(n_1538),
.B1(n_1533),
.B2(n_1473),
.C(n_1418),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1674),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1586),
.A2(n_1533),
.B(n_1426),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1598),
.A2(n_1417),
.B1(n_1543),
.B2(n_1590),
.C(n_1636),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1577),
.B(n_1603),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1584),
.B(n_1650),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1606),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1634),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1578),
.B(n_1629),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_SL g1697 ( 
.A(n_1576),
.B(n_1578),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1606),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1621),
.B(n_1649),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1621),
.B(n_1649),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1643),
.B(n_1571),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1646),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1628),
.B(n_1613),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1571),
.B(n_1617),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1582),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1653),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_SL g1707 ( 
.A(n_1576),
.B(n_1642),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1653),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1669),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1655),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_SL g1711 ( 
.A1(n_1580),
.A2(n_1607),
.B(n_1636),
.C(n_1637),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1607),
.A2(n_1642),
.B1(n_1638),
.B2(n_1583),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1583),
.A2(n_1591),
.B1(n_1631),
.B2(n_1617),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1666),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1655),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1629),
.B(n_1591),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1637),
.A2(n_1631),
.B(n_1628),
.C(n_1626),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1647),
.A2(n_1626),
.B1(n_1638),
.B2(n_1568),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1647),
.A2(n_1642),
.B1(n_1569),
.B2(n_1615),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1671),
.B(n_1623),
.Y(n_1720)
);

AO21x1_ASAP7_75t_L g1721 ( 
.A1(n_1639),
.A2(n_1641),
.B(n_1635),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1623),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1600),
.B(n_1601),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1596),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1628),
.A2(n_1635),
.B(n_1644),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_SL g1726 ( 
.A1(n_1639),
.A2(n_1641),
.B(n_1660),
.C(n_1672),
.Y(n_1726)
);

O2A1O1Ixp33_ASAP7_75t_L g1727 ( 
.A1(n_1644),
.A2(n_1573),
.B(n_1639),
.C(n_1615),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1615),
.A2(n_1627),
.B(n_1633),
.C(n_1672),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1579),
.A2(n_1658),
.B(n_1611),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1615),
.A2(n_1627),
.B(n_1633),
.C(n_1668),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1599),
.Y(n_1731)
);

OAI31xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1611),
.A2(n_1613),
.A3(n_1609),
.B(n_1610),
.Y(n_1732)
);

OR2x6_ASAP7_75t_L g1733 ( 
.A(n_1613),
.B(n_1609),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1619),
.B(n_1622),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1664),
.A2(n_1670),
.B1(n_1569),
.B2(n_1630),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1567),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1614),
.B(n_1616),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1666),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1614),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1584),
.B(n_1650),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1584),
.B(n_1651),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1655),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1610),
.B(n_1595),
.Y(n_1743)
);

AO32x2_ASAP7_75t_L g1744 ( 
.A1(n_1667),
.A2(n_1605),
.A3(n_1595),
.B1(n_1608),
.B2(n_1589),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1584),
.B(n_1651),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1618),
.B(n_1605),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1630),
.Y(n_1747)
);

AO21x2_ASAP7_75t_L g1748 ( 
.A1(n_1572),
.A2(n_1597),
.B(n_1608),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1693),
.B(n_1581),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1739),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1706),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1724),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1736),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1720),
.B(n_1625),
.Y(n_1754)
);

INVx3_ASAP7_75t_SL g1755 ( 
.A(n_1747),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1691),
.A2(n_1654),
.B1(n_1648),
.B2(n_1674),
.C(n_1673),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1733),
.B(n_1608),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1736),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1733),
.B(n_1608),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1706),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1722),
.B(n_1625),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1733),
.B(n_1703),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1709),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1693),
.Y(n_1764)
);

AND2x4_ASAP7_75t_SL g1765 ( 
.A(n_1693),
.B(n_1592),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1697),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1710),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1677),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1696),
.B(n_1585),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1716),
.B(n_1640),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1703),
.B(n_1581),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1737),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1705),
.B(n_1567),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1727),
.B(n_1669),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1677),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1703),
.B(n_1581),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1677),
.B(n_1581),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1708),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1712),
.A2(n_1627),
.B1(n_1620),
.B2(n_1569),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1688),
.A2(n_1678),
.B1(n_1735),
.B2(n_1679),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1705),
.B(n_1570),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1723),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1695),
.B(n_1570),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1708),
.B(n_1575),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1690),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1677),
.B(n_1592),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1718),
.A2(n_1627),
.B1(n_1620),
.B2(n_1569),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1682),
.A2(n_1620),
.B1(n_1665),
.B2(n_1656),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1734),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1695),
.B(n_1574),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1727),
.B(n_1669),
.Y(n_1791)
);

A2O1A1Ixp33_ASAP7_75t_SL g1792 ( 
.A1(n_1686),
.A2(n_1599),
.B(n_1632),
.C(n_1645),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1774),
.B(n_1731),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1717),
.C(n_1711),
.Y(n_1795)
);

INVx4_ASAP7_75t_L g1796 ( 
.A(n_1755),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1769),
.B(n_1701),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1769),
.B(n_1704),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1764),
.B(n_1740),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1792),
.A2(n_1711),
.B(n_1717),
.Y(n_1800)
);

CKINVDCx14_ASAP7_75t_R g1801 ( 
.A(n_1770),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1702),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1772),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1771),
.B(n_1740),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

OAI222xp33_ASAP7_75t_L g1806 ( 
.A1(n_1756),
.A2(n_1713),
.B1(n_1719),
.B2(n_1743),
.C1(n_1676),
.C2(n_1686),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1771),
.B(n_1740),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1764),
.B(n_1741),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1752),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1764),
.B(n_1741),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1784),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1749),
.B(n_1745),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1763),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1784),
.Y(n_1814)
);

AOI322xp5_ASAP7_75t_L g1815 ( 
.A1(n_1780),
.A2(n_1687),
.A3(n_1681),
.B1(n_1738),
.B2(n_1692),
.C1(n_1699),
.C2(n_1700),
.Y(n_1815)
);

AND2x4_ASAP7_75t_SL g1816 ( 
.A(n_1793),
.B(n_1738),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1768),
.A2(n_1725),
.B1(n_1730),
.B2(n_1728),
.C(n_1729),
.Y(n_1817)
);

AOI322xp5_ASAP7_75t_L g1818 ( 
.A1(n_1779),
.A2(n_1687),
.A3(n_1681),
.B1(n_1702),
.B2(n_1694),
.C1(n_1698),
.C2(n_1684),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1749),
.B(n_1690),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1752),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1754),
.B(n_1743),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1753),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1765),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1749),
.B(n_1690),
.Y(n_1824)
);

INVx5_ASAP7_75t_SL g1825 ( 
.A(n_1785),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1752),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1768),
.A2(n_1728),
.B1(n_1730),
.B2(n_1721),
.C(n_1726),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1755),
.A2(n_1714),
.B1(n_1675),
.B2(n_1747),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1753),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1777),
.B(n_1744),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1774),
.B(n_1731),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1758),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1758),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1754),
.B(n_1746),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1766),
.B(n_1714),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1777),
.B(n_1744),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1750),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1777),
.B(n_1744),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_L g1839 ( 
.A(n_1787),
.B(n_1732),
.C(n_1680),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1761),
.B(n_1789),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1771),
.B(n_1744),
.Y(n_1841)
);

NOR2x1p5_ASAP7_75t_L g1842 ( 
.A(n_1767),
.B(n_1710),
.Y(n_1842)
);

AND3x1_ASAP7_75t_L g1843 ( 
.A(n_1787),
.B(n_1673),
.C(n_1689),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1789),
.B(n_1748),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1788),
.A2(n_1620),
.B1(n_1685),
.B2(n_1654),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1765),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1789),
.B(n_1748),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1830),
.B(n_1775),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1837),
.Y(n_1849)
);

AND2x4_ASAP7_75t_SL g1850 ( 
.A(n_1796),
.B(n_1793),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1842),
.B(n_1762),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1809),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1837),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1842),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1799),
.B(n_1762),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1822),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1799),
.B(n_1762),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1811),
.B(n_1775),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1816),
.Y(n_1859)
);

OAI33xp33_ASAP7_75t_L g1860 ( 
.A1(n_1795),
.A2(n_1783),
.A3(n_1790),
.B1(n_1781),
.B2(n_1773),
.B3(n_1766),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1800),
.B(n_1791),
.C(n_1785),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1808),
.B(n_1757),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1822),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1808),
.B(n_1757),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1811),
.B(n_1778),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1801),
.B(n_1683),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_R g1867 ( 
.A(n_1796),
.B(n_1715),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1809),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1820),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1814),
.B(n_1772),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1830),
.B(n_1757),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1836),
.B(n_1759),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1814),
.B(n_1778),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1820),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1836),
.B(n_1759),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1839),
.B(n_1791),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1803),
.B(n_1751),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1826),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1838),
.B(n_1759),
.Y(n_1879)
);

INVxp67_ASAP7_75t_L g1880 ( 
.A(n_1805),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1829),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1829),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1832),
.B(n_1751),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1832),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1819),
.B(n_1776),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1816),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1810),
.B(n_1776),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1833),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1819),
.B(n_1776),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1794),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1838),
.B(n_1786),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1840),
.B(n_1760),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1826),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1840),
.B(n_1760),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1833),
.B(n_1782),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1880),
.B(n_1798),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1881),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1851),
.B(n_1824),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1858),
.B(n_1844),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1881),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1856),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1880),
.B(n_1797),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1851),
.B(n_1854),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1856),
.Y(n_1904)
);

O2A1O1Ixp33_ASAP7_75t_SL g1905 ( 
.A1(n_1861),
.A2(n_1680),
.B(n_1806),
.C(n_1815),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1852),
.Y(n_1906)
);

AOI322xp5_ASAP7_75t_L g1907 ( 
.A1(n_1848),
.A2(n_1827),
.A3(n_1817),
.B1(n_1841),
.B2(n_1786),
.C1(n_1835),
.C2(n_1845),
.Y(n_1907)
);

INVxp33_ASAP7_75t_L g1908 ( 
.A(n_1867),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1851),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1863),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1859),
.B(n_1821),
.Y(n_1911)
);

NAND2xp67_ASAP7_75t_SL g1912 ( 
.A(n_1848),
.B(n_1824),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1859),
.B(n_1821),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1858),
.B(n_1844),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1863),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1852),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1851),
.B(n_1841),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1873),
.B(n_1847),
.Y(n_1918)
);

NOR2xp67_ASAP7_75t_L g1919 ( 
.A(n_1861),
.B(n_1796),
.Y(n_1919)
);

INVx4_ASAP7_75t_L g1920 ( 
.A(n_1876),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1854),
.B(n_1804),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1882),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1882),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1852),
.Y(n_1924)
);

AND2x4_ASAP7_75t_SL g1925 ( 
.A(n_1854),
.B(n_1813),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1873),
.B(n_1847),
.Y(n_1926)
);

NAND2x1p5_ASAP7_75t_L g1927 ( 
.A(n_1890),
.B(n_1843),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1884),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1850),
.B(n_1804),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1884),
.Y(n_1930)
);

NAND2x1p5_ASAP7_75t_L g1931 ( 
.A(n_1890),
.B(n_1785),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1888),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1888),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1855),
.B(n_1804),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1849),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1855),
.B(n_1807),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1886),
.B(n_1834),
.Y(n_1937)
);

NOR3xp33_ASAP7_75t_L g1938 ( 
.A(n_1860),
.B(n_1828),
.C(n_1802),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1857),
.B(n_1807),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1857),
.B(n_1807),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1886),
.B(n_1834),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1849),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1850),
.B(n_1812),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1876),
.B(n_1818),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1876),
.A2(n_1845),
.B1(n_1828),
.B2(n_1785),
.Y(n_1945)
);

NAND2x1_ASAP7_75t_L g1946 ( 
.A(n_1920),
.B(n_1876),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1901),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1904),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1938),
.B(n_1876),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1907),
.B(n_1876),
.C(n_1785),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1910),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1925),
.B(n_1850),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1917),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1929),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1915),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1911),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1937),
.B(n_1865),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1929),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1941),
.B(n_1865),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1944),
.B(n_1870),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1905),
.A2(n_1860),
.B(n_1785),
.C(n_1866),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1925),
.B(n_1848),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1903),
.B(n_1890),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1913),
.B(n_1870),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1902),
.B(n_1887),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1896),
.B(n_1887),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1918),
.B(n_1877),
.Y(n_1967)
);

INVx4_ASAP7_75t_L g1968 ( 
.A(n_1920),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1927),
.B(n_1871),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1927),
.B(n_1871),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1919),
.B(n_1877),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1918),
.B(n_1892),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1945),
.A2(n_1785),
.B1(n_1885),
.B2(n_1889),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1922),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1917),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1908),
.B(n_1871),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1903),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1908),
.B(n_1872),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1920),
.B(n_1872),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1912),
.B(n_1853),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1927),
.B(n_1872),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1921),
.B(n_1875),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_SL g1983 ( 
.A(n_1897),
.B(n_1883),
.C(n_1895),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1934),
.B(n_1936),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1905),
.B(n_1685),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1929),
.B(n_1812),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1951),
.Y(n_1987)
);

AOI22xp33_ASAP7_75t_SL g1988 ( 
.A1(n_1950),
.A2(n_1909),
.B1(n_1921),
.B2(n_1707),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1951),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1949),
.B(n_1934),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1974),
.Y(n_1991)
);

AOI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1961),
.A2(n_1909),
.B1(n_1900),
.B2(n_1942),
.C(n_1923),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1974),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1947),
.Y(n_1994)
);

OAI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1946),
.A2(n_1909),
.B1(n_1831),
.B2(n_1794),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1962),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1985),
.A2(n_1943),
.B1(n_1898),
.B2(n_1889),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1948),
.Y(n_1998)
);

INVxp67_ASAP7_75t_SL g1999 ( 
.A(n_1954),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1962),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1977),
.B(n_1936),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1955),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1956),
.B(n_1939),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1960),
.A2(n_1831),
.B(n_1794),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1984),
.B(n_1943),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1976),
.B(n_1943),
.Y(n_2006)
);

INVxp33_ASAP7_75t_SL g2007 ( 
.A(n_1978),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_1952),
.Y(n_2008)
);

INVxp67_ASAP7_75t_L g2009 ( 
.A(n_1971),
.Y(n_2009)
);

NAND3xp33_ASAP7_75t_L g2010 ( 
.A(n_1983),
.B(n_1930),
.C(n_1928),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1954),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1957),
.B(n_1932),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1984),
.B(n_1939),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1952),
.B(n_1940),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1952),
.A2(n_1898),
.B1(n_1940),
.B2(n_1831),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1973),
.A2(n_1825),
.B1(n_1885),
.B2(n_1889),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1999),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1992),
.A2(n_1946),
.B(n_1980),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2007),
.B(n_2008),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_SL g2020 ( 
.A1(n_2007),
.A2(n_1968),
.B1(n_1954),
.B2(n_1958),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1996),
.B(n_1953),
.Y(n_2021)
);

XNOR2x2_ASAP7_75t_L g2022 ( 
.A(n_2010),
.B(n_1969),
.Y(n_2022)
);

O2A1O1Ixp5_ASAP7_75t_L g2023 ( 
.A1(n_2011),
.A2(n_1968),
.B(n_1958),
.C(n_1979),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1990),
.B(n_1965),
.Y(n_2024)
);

NAND3x2_ASAP7_75t_L g2025 ( 
.A(n_2014),
.B(n_1970),
.C(n_1969),
.Y(n_2025)
);

NAND3xp33_ASAP7_75t_L g2026 ( 
.A(n_2009),
.B(n_1968),
.C(n_1959),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_2005),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1987),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1996),
.B(n_1953),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1987),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1988),
.A2(n_1964),
.B(n_1970),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2000),
.B(n_1975),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_1998),
.A2(n_1981),
.B1(n_1957),
.B2(n_1959),
.C(n_1967),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2000),
.B(n_1975),
.Y(n_2034)
);

AOI222xp33_ASAP7_75t_L g2035 ( 
.A1(n_2003),
.A2(n_1981),
.B1(n_1982),
.B2(n_1966),
.C1(n_1958),
.C2(n_1963),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1993),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2011),
.B(n_1963),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_2006),
.A2(n_1986),
.B1(n_1963),
.B2(n_1967),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1993),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_2014),
.B(n_1972),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_2019),
.B(n_2001),
.Y(n_2041)
);

AOI21xp33_ASAP7_75t_SL g2042 ( 
.A1(n_2020),
.A2(n_1995),
.B(n_2016),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2040),
.B(n_2013),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_2022),
.A2(n_1994),
.B1(n_2002),
.B2(n_1991),
.Y(n_2044)
);

AOI222xp33_ASAP7_75t_L g2045 ( 
.A1(n_2033),
.A2(n_2002),
.B1(n_1994),
.B2(n_1989),
.C1(n_1997),
.C2(n_2005),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2033),
.A2(n_2004),
.B1(n_2012),
.B2(n_2015),
.C(n_2013),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_2017),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2025),
.A2(n_2012),
.B1(n_1972),
.B2(n_1825),
.Y(n_2048)
);

O2A1O1Ixp33_ASAP7_75t_SL g2049 ( 
.A1(n_2018),
.A2(n_1935),
.B(n_1933),
.C(n_1883),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2027),
.B(n_1875),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2021),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2029),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2023),
.Y(n_2053)
);

AOI322xp5_ASAP7_75t_L g2054 ( 
.A1(n_2038),
.A2(n_1891),
.A3(n_1875),
.B1(n_1879),
.B2(n_1786),
.C1(n_1912),
.C2(n_1885),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2035),
.B(n_1879),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2032),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_2047),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2044),
.A2(n_2026),
.B1(n_2031),
.B2(n_2024),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_2047),
.Y(n_2059)
);

NOR2xp67_ASAP7_75t_L g2060 ( 
.A(n_2053),
.B(n_2037),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_2041),
.B(n_2034),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_2043),
.Y(n_2062)
);

NAND4xp25_ASAP7_75t_L g2063 ( 
.A(n_2044),
.B(n_2023),
.C(n_2031),
.D(n_2036),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2045),
.B(n_2028),
.Y(n_2064)
);

NOR2xp67_ASAP7_75t_L g2065 ( 
.A(n_2042),
.B(n_2030),
.Y(n_2065)
);

NAND4xp25_ASAP7_75t_L g2066 ( 
.A(n_2046),
.B(n_2039),
.C(n_1742),
.D(n_1715),
.Y(n_2066)
);

NOR3x1_ASAP7_75t_L g2067 ( 
.A(n_2048),
.B(n_1926),
.C(n_1914),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_SL g2068 ( 
.A(n_2055),
.B(n_1931),
.C(n_1926),
.Y(n_2068)
);

AND4x1_ASAP7_75t_L g2069 ( 
.A(n_2051),
.B(n_1879),
.C(n_1891),
.D(n_1864),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2050),
.Y(n_2070)
);

NAND5xp2_ASAP7_75t_L g2071 ( 
.A(n_2058),
.B(n_2049),
.C(n_2052),
.D(n_2056),
.E(n_2054),
.Y(n_2071)
);

NOR3xp33_ASAP7_75t_L g2072 ( 
.A(n_2064),
.B(n_1916),
.C(n_1906),
.Y(n_2072)
);

O2A1O1Ixp33_ASAP7_75t_L g2073 ( 
.A1(n_2063),
.A2(n_1931),
.B(n_1924),
.C(n_1916),
.Y(n_2073)
);

AOI221xp5_ASAP7_75t_SL g2074 ( 
.A1(n_2066),
.A2(n_1924),
.B1(n_1906),
.B2(n_1914),
.C(n_1899),
.Y(n_2074)
);

NAND4xp25_ASAP7_75t_SL g2075 ( 
.A(n_2070),
.B(n_1899),
.C(n_1891),
.D(n_1862),
.Y(n_2075)
);

OAI211xp5_ASAP7_75t_L g2076 ( 
.A1(n_2065),
.A2(n_1767),
.B(n_1742),
.C(n_1894),
.Y(n_2076)
);

AOI32xp33_ASAP7_75t_L g2077 ( 
.A1(n_2061),
.A2(n_1885),
.A3(n_1889),
.B1(n_1864),
.B2(n_1862),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2060),
.B(n_1853),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_R g2079 ( 
.A(n_2059),
.B(n_1599),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2078),
.Y(n_2080)
);

OAI221xp5_ASAP7_75t_L g2081 ( 
.A1(n_2074),
.A2(n_2062),
.B1(n_2057),
.B2(n_2068),
.C(n_2069),
.Y(n_2081)
);

NAND4xp75_ASAP7_75t_L g2082 ( 
.A(n_2071),
.B(n_2067),
.C(n_2057),
.D(n_1846),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2073),
.A2(n_1931),
.B(n_1895),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_L g2084 ( 
.A(n_2076),
.B(n_1767),
.C(n_1658),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2072),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2075),
.A2(n_1825),
.B1(n_1846),
.B2(n_1823),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2079),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_2087),
.Y(n_2088)
);

OAI322xp33_ASAP7_75t_L g2089 ( 
.A1(n_2081),
.A2(n_2077),
.A3(n_1894),
.B1(n_1892),
.B2(n_1878),
.C1(n_1893),
.C2(n_1874),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2085),
.Y(n_2090)
);

XOR2xp5_ASAP7_75t_L g2091 ( 
.A(n_2082),
.B(n_1656),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2080),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2084),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2090),
.B(n_2086),
.Y(n_2094)
);

NOR3xp33_ASAP7_75t_SL g2095 ( 
.A(n_2089),
.B(n_2083),
.C(n_1790),
.Y(n_2095)
);

AOI21xp33_ASAP7_75t_SL g2096 ( 
.A1(n_2088),
.A2(n_1823),
.B(n_1878),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_2088),
.B(n_1825),
.Y(n_2097)
);

AOI221xp5_ASAP7_75t_SL g2098 ( 
.A1(n_2096),
.A2(n_2093),
.B1(n_2091),
.B2(n_2092),
.C(n_1878),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2094),
.B(n_1868),
.Y(n_2099)
);

AO22x2_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_2097),
.B1(n_2095),
.B2(n_1893),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_2100),
.B(n_2098),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2100),
.Y(n_2102)
);

INVx1_ASAP7_75t_SL g2103 ( 
.A(n_2101),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_2102),
.A2(n_1893),
.B1(n_1874),
.B2(n_1869),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2103),
.A2(n_1874),
.B(n_1869),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2105),
.A2(n_2104),
.B1(n_1869),
.B2(n_1868),
.Y(n_2106)
);

AOI31xp33_ASAP7_75t_L g2107 ( 
.A1(n_2106),
.A2(n_1663),
.A3(n_1659),
.B(n_1657),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2107),
.Y(n_2108)
);

AOI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_2108),
.A2(n_1868),
.B1(n_1726),
.B2(n_1783),
.C(n_1781),
.Y(n_2109)
);

AOI211xp5_ASAP7_75t_L g2110 ( 
.A1(n_2109),
.A2(n_1661),
.B(n_1662),
.C(n_1587),
.Y(n_2110)
);


endmodule