module real_jpeg_17429_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_662, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_662;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_634;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_431;
wire n_357;
wire n_420;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_1),
.A2(n_141),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_1),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_1),
.A2(n_194),
.B1(n_341),
.B2(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_1),
.A2(n_341),
.B1(n_418),
.B2(n_479),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_1),
.A2(n_275),
.B1(n_341),
.B2(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_2),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_2),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_3),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_63),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_3),
.A2(n_63),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_3),
.A2(n_63),
.B1(n_580),
.B2(n_583),
.Y(n_579)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_5),
.A2(n_107),
.B1(n_212),
.B2(n_223),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_5),
.A2(n_107),
.B1(n_601),
.B2(n_604),
.Y(n_600)
);

AO22x1_ASAP7_75t_L g643 ( 
.A1(n_5),
.A2(n_107),
.B1(n_644),
.B2(n_647),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_6),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_8),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_8),
.A2(n_140),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_8),
.A2(n_140),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_8),
.A2(n_140),
.B1(n_485),
.B2(n_488),
.Y(n_484)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g395 ( 
.A(n_9),
.Y(n_395)
);

AOI22x1_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_152),
.B1(n_158),
.B2(n_160),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_10),
.A2(n_148),
.B1(n_160),
.B2(n_239),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_10),
.A2(n_160),
.B1(n_266),
.B2(n_270),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_10),
.A2(n_160),
.B1(n_389),
.B2(n_393),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_11),
.A2(n_147),
.B1(n_190),
.B2(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_11),
.A2(n_147),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_11),
.A2(n_147),
.B1(n_393),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_12),
.B(n_261),
.Y(n_401)
);

OAI32xp33_ASAP7_75t_L g422 ( 
.A1(n_12),
.A2(n_169),
.A3(n_423),
.B1(n_426),
.B2(n_431),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_12),
.B(n_199),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_12),
.A2(n_82),
.B1(n_443),
.B2(n_528),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_12),
.A2(n_314),
.B1(n_547),
.B2(n_550),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_13),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_13),
.A2(n_96),
.B1(n_212),
.B2(n_217),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_13),
.A2(n_96),
.B1(n_152),
.B2(n_588),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_13),
.A2(n_96),
.B1(n_258),
.B2(n_634),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_14),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_15),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_15),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_15),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_15),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_16),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_16),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_16),
.A2(n_257),
.B1(n_355),
.B2(n_358),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_16),
.A2(n_257),
.B1(n_498),
.B2(n_500),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_16),
.A2(n_257),
.B1(n_489),
.B2(n_510),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_17),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_17),
.A2(n_74),
.B1(n_158),
.B2(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_17),
.A2(n_74),
.B1(n_275),
.B2(n_280),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_17),
.A2(n_74),
.B1(n_364),
.B2(n_595),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_18),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_18),
.Y(n_177)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_19),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_19),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g149 ( 
.A(n_19),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g597 ( 
.A(n_19),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_656),
.B(n_658),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_570),
.B(n_649),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_405),
.B(n_565),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_294),
.C(n_344),
.Y(n_27)
);

A2O1A1O1Ixp25_ASAP7_75t_L g565 ( 
.A1(n_28),
.A2(n_294),
.B(n_566),
.C(n_568),
.D(n_569),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_244),
.Y(n_28)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_29),
.B(n_244),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_200),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_30),
.B(n_621),
.C(n_622),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_108),
.C(n_150),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_31),
.B(n_247),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_64),
.B(n_80),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_32),
.B(n_64),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_57),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_33),
.A2(n_65),
.B1(n_210),
.B2(n_222),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_33),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_33),
.A2(n_65),
.B1(n_368),
.B2(n_373),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_33),
.A2(n_65),
.B1(n_474),
.B2(n_478),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_33),
.A2(n_65),
.B1(n_478),
.B2(n_497),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_33),
.A2(n_65),
.B1(n_415),
.B2(n_497),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g576 ( 
.A1(n_33),
.A2(n_65),
.B(n_222),
.Y(n_576)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_46),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_40),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_41),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_43),
.Y(n_487)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_43),
.Y(n_512)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_46)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_47),
.Y(n_416)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_47),
.Y(n_477)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_48),
.Y(n_372)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_48),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_53),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_56),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_58),
.A2(n_66),
.B1(n_242),
.B2(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_60),
.Y(n_499)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_66),
.A2(n_68),
.B1(n_211),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_66),
.A2(n_242),
.B1(n_414),
.B2(n_419),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_66),
.B(n_314),
.Y(n_536)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_73),
.Y(n_272)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_78),
.Y(n_226)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_79),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_80),
.B(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_91),
.B1(n_101),
.B2(n_103),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_81),
.A2(n_331),
.B1(n_388),
.B2(n_396),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_81),
.A2(n_388),
.B1(n_438),
.B2(n_442),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_81),
.A2(n_508),
.B1(n_513),
.B2(n_514),
.Y(n_507)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_82),
.A2(n_104),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_82),
.A2(n_92),
.B1(n_274),
.B2(n_283),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_82),
.A2(n_274),
.B1(n_330),
.B2(n_337),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_82),
.A2(n_484),
.B1(n_491),
.B2(n_492),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_82),
.A2(n_509),
.B1(n_528),
.B2(n_535),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_83),
.Y(n_491)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_87),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_89),
.Y(n_441)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_90),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_90),
.Y(n_336)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_90),
.Y(n_456)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_100),
.Y(n_279)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_100),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_102),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_109),
.B(n_150),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_123),
.B1(n_136),
.B2(n_144),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_110),
.A2(n_123),
.B1(n_144),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_110),
.A2(n_136),
.B1(n_253),
.B2(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_110),
.A2(n_238),
.B1(n_260),
.B2(n_579),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_110),
.A2(n_260),
.B1(n_632),
.B2(n_633),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_110),
.A2(n_260),
.B1(n_633),
.B2(n_642),
.Y(n_641)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_111),
.A2(n_261),
.B1(n_340),
.B2(n_343),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_111),
.A2(n_261),
.B1(n_340),
.B2(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_111),
.A2(n_261),
.B1(n_593),
.B2(n_594),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_111),
.A2(n_261),
.B(n_643),
.Y(n_657)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_119),
.B(n_123),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_116),
.Y(n_634)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_118),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_119),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_123),
.Y(n_261)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_128),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_129),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_129),
.Y(n_323)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_135),
.Y(n_319)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_139),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_139),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_141),
.B(n_314),
.Y(n_313)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_148),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

OAI22x1_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_161),
.B1(n_189),
.B2(n_198),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_151),
.A2(n_161),
.B1(n_198),
.B2(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_157),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_161),
.A2(n_198),
.B1(n_286),
.B2(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_161),
.A2(n_198),
.B1(n_382),
.B2(n_546),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_161),
.A2(n_198),
.B1(n_206),
.B2(n_587),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_161),
.A2(n_198),
.B1(n_587),
.B2(n_600),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_169),
.B(n_178),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_175),
.Y(n_603)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_176),
.Y(n_360)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_176),
.Y(n_430)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_176),
.Y(n_549)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_177),
.Y(n_310)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_177),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_181),
.B1(n_185),
.B2(n_187),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_180),
.Y(n_454)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_185),
.Y(n_464)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_196),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_197),
.Y(n_357)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_199),
.A2(n_203),
.B1(n_307),
.B2(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_199),
.A2(n_203),
.B1(n_354),
.B2(n_381),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_199),
.A2(n_203),
.B(n_630),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_228),
.Y(n_200)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_201),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_209),
.B(n_227),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_209),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_213),
.Y(n_370)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_227),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_227),
.A2(n_613),
.B1(n_615),
.B2(n_625),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_228),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_240),
.B2(n_243),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_231),
.A2(n_232),
.B1(n_241),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_231),
.A2(n_243),
.B1(n_617),
.B2(n_662),
.Y(n_616)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_234),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_236),
.Y(n_618)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_250),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.C(n_285),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_252),
.B(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_273),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_264),
.B(n_273),
.Y(n_351)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_265),
.Y(n_373)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_267),
.Y(n_418)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_295),
.B(n_298),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_303),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_301),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_311),
.C(n_339),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_339),
.Y(n_350)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_329),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_329),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_315),
.B1(n_324),
.B2(n_328),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_SL g362 ( 
.A1(n_313),
.A2(n_314),
.B(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_314),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_314),
.B(n_463),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_SL g474 ( 
.A1(n_314),
.A2(n_462),
.B(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_314),
.B(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_337),
.Y(n_513)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_347),
.B(n_374),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_345),
.B(n_347),
.C(n_567),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.C(n_352),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_348),
.A2(n_349),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_352),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_361),
.C(n_367),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_367),
.Y(n_377)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx2_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g584 ( 
.A(n_365),
.Y(n_584)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_366),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_368),
.Y(n_419)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_402),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_375),
.B(n_402),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.C(n_379),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_379),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_387),
.C(n_401),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_383),
.Y(n_551)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_401),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_399),
.Y(n_444)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_403),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_445),
.B(n_564),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_407),
.B(n_409),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_413),
.C(n_420),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_410),
.A2(n_411),
.B1(n_559),
.B2(n_560),
.Y(n_558)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_413),
.A2(n_420),
.B1(n_421),
.B2(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_413),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_436),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_422),
.A2(n_436),
.B1(n_437),
.B2(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_422),
.Y(n_555)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_557),
.B(n_563),
.Y(n_445)
);

AOI21x1_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_540),
.B(n_556),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_505),
.B(n_539),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_482),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_449),
.B(n_482),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_472),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_450),
.A2(n_472),
.B1(n_473),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

OAI32xp33_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_455),
.A3(n_457),
.B1(n_462),
.B2(n_465),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx8_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_493),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_483),
.B(n_495),
.C(n_504),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_484),
.Y(n_514)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_504),
.Y(n_493)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_517),
.B(n_538),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_515),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_515),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_512),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_533),
.B(n_537),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_527),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_525),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_536),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_536),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_542),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_542),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_554),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_544),
.A2(n_545),
.B1(n_552),
.B2(n_553),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_553),
.C(n_554),
.Y(n_562)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_562),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_558),
.B(n_562),
.Y(n_563)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NOR3xp33_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_626),
.C(n_639),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_619),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_573),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_573),
.A2(n_652),
.B(n_653),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_SL g573 ( 
.A(n_574),
.B(n_612),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_574),
.B(n_612),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_590),
.Y(n_574)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_575),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_577),
.C(n_585),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_576),
.A2(n_599),
.B1(n_608),
.B2(n_609),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_576),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_576),
.B(n_586),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_576),
.B(n_592),
.C(n_609),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_577),
.A2(n_591),
.B1(n_610),
.B2(n_611),
.Y(n_590)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_577),
.Y(n_610)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

XNOR2x1_ASAP7_75t_L g613 ( 
.A(n_578),
.B(n_614),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_579),
.Y(n_593)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_591),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_591),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_598),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_594),
.Y(n_632)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_599),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_600),
.Y(n_630)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_610),
.B(n_637),
.C(n_638),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_615),
.C(n_616),
.Y(n_612)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_613),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_616),
.B(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_620),
.B(n_623),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_620),
.B(n_623),
.Y(n_652)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

A2O1A1O1Ixp25_ASAP7_75t_L g650 ( 
.A1(n_627),
.A2(n_640),
.B(n_651),
.C(n_654),
.D(n_655),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_628),
.B(n_636),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_628),
.B(n_636),
.Y(n_654)
);

BUFx24_ASAP7_75t_SL g661 ( 
.A(n_628),
.Y(n_661)
);

FAx1_ASAP7_75t_SL g628 ( 
.A(n_629),
.B(n_631),
.CI(n_635),
.CON(n_628),
.SN(n_628)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_631),
.C(n_635),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_634),
.Y(n_647)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_648),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_648),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_641),
.B(n_657),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_641),
.B(n_657),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g642 ( 
.A(n_643),
.Y(n_642)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g658 ( 
.A(n_659),
.Y(n_658)
);


endmodule