module fake_jpeg_21396_n_54 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_54);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_54;

wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_8),
.B1(n_20),
.B2(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_26),
.B1(n_11),
.B2(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_7),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_25),
.B(n_27),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_24),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_24),
.C(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

XNOR2x1_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_47),
.B1(n_42),
.B2(n_39),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_40),
.C(n_5),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_9),
.C1(n_13),
.C2(n_15),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_21),
.B(n_4),
.C(n_6),
.Y(n_54)
);


endmodule