module fake_jpeg_8806_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_4),
.B(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_17),
.C(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_50),
.C(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_55),
.B1(n_19),
.B2(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_17),
.C(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_22),
.B1(n_23),
.B2(n_17),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.C(n_37),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_19),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_0),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_27),
.B1(n_24),
.B2(n_39),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_40),
.B(n_37),
.C(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_81),
.B1(n_82),
.B2(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_38),
.B1(n_23),
.B2(n_25),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_83),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_25),
.B1(n_64),
.B2(n_60),
.Y(n_76)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_94),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_2),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_40),
.Y(n_107)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_31),
.B1(n_30),
.B2(n_20),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_11),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_58),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_73),
.C(n_74),
.Y(n_141)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_111),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_1),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_80),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_77),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_78),
.B1(n_84),
.B2(n_90),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_117),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_1),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_121),
.Y(n_144)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_21),
.B(n_26),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_83),
.B1(n_89),
.B2(n_91),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_137),
.B1(n_152),
.B2(n_112),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_151),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_81),
.B1(n_92),
.B2(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_136),
.B1(n_138),
.B2(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_130),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_134),
.B(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_73),
.B(n_72),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_148),
.B(n_111),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_102),
.B1(n_117),
.B2(n_105),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_75),
.B1(n_72),
.B2(n_69),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_72),
.B1(n_85),
.B2(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_100),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_109),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_153),
.Y(n_166)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_72),
.B(n_26),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_2),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_123),
.B(n_97),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_112),
.B(n_110),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_2),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_90),
.B1(n_26),
.B2(n_6),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_3),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_155),
.B(n_164),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_159),
.B(n_168),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_171),
.C(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_141),
.B1(n_125),
.B2(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_173),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_115),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_178),
.B(n_127),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_101),
.C(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_150),
.B1(n_131),
.B2(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_SL g178 ( 
.A(n_128),
.B(n_121),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_101),
.C(n_110),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_182),
.C(n_149),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_129),
.B(n_3),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_104),
.B(n_6),
.C(n_7),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_96),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_208),
.B1(n_211),
.B2(n_182),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_154),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_164),
.B1(n_174),
.B2(n_158),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_8),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_163),
.B1(n_155),
.B2(n_167),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_233)
);

OAI221xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_143),
.B1(n_150),
.B2(n_149),
.C(n_110),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_142),
.B1(n_143),
.B2(n_96),
.Y(n_208)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_227),
.B1(n_205),
.B2(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_228),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_187),
.B(n_172),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_187),
.B(n_195),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_171),
.B1(n_161),
.B2(n_165),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_165),
.C(n_7),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_234),
.C(n_204),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_235),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_195),
.B1(n_211),
.B2(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_193),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_245),
.C(n_252),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_207),
.B1(n_197),
.B2(n_188),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_250),
.B1(n_251),
.B2(n_215),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_210),
.C(n_196),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_247),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_199),
.B(n_189),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_224),
.B(n_221),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_189),
.B1(n_209),
.B2(n_203),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_211),
.B1(n_200),
.B2(n_10),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_211),
.C(n_9),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_233),
.B1(n_226),
.B2(n_223),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_264),
.B1(n_253),
.B2(n_243),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_262),
.B(n_267),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_230),
.C(n_216),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_229),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_224),
.C(n_222),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_240),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_211),
.C(n_9),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_10),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_8),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_10),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_239),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_271),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_239),
.Y(n_271)
);

AOI321xp33_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_249),
.A3(n_256),
.B1(n_259),
.B2(n_236),
.C(n_242),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_266),
.B(n_13),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_11),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_285),
.B(n_12),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_12),
.Y(n_285)
);

CKINVDCx12_ASAP7_75t_R g286 ( 
.A(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_271),
.C(n_270),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_293),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_12),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_296),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_283),
.A3(n_290),
.B1(n_292),
.B2(n_280),
.C1(n_281),
.C2(n_16),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_301),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_302),
.B(n_297),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_13),
.B1(n_15),
.B2(n_298),
.Y(n_304)
);


endmodule