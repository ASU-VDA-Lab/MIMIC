module fake_jpeg_2819_n_436 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_436);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_436;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx11_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_50),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_19),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_66),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_64),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_76),
.Y(n_93)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_35),
.A2(n_12),
.B(n_1),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_69),
.Y(n_103)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_72),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_71),
.B(n_73),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_77),
.Y(n_110)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_24),
.B(n_32),
.CON(n_75),
.SN(n_75)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_78),
.B1(n_80),
.B2(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_79),
.B(n_83),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_82),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_34),
.B(n_12),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_12),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_46),
.B1(n_30),
.B2(n_41),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_24),
.B(n_0),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_37),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_0),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_67),
.B1(n_51),
.B2(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_95),
.A2(n_98),
.B1(n_106),
.B2(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_32),
.B1(n_21),
.B2(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_26),
.B1(n_25),
.B2(n_43),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_100),
.A2(n_118),
.B1(n_139),
.B2(n_7),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_38),
.B1(n_44),
.B2(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_39),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_115),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_54),
.A2(n_38),
.B1(n_40),
.B2(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_40),
.B1(n_25),
.B2(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_46),
.B1(n_30),
.B2(n_41),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_46),
.B1(n_22),
.B2(n_41),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_81),
.B1(n_47),
.B2(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_46),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_22),
.B1(n_46),
.B2(n_36),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_46),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_128),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_36),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_49),
.B(n_36),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_137),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_31),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_52),
.A2(n_22),
.B1(n_31),
.B2(n_29),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_57),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_6),
.Y(n_175)
);

NOR4xp25_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_72),
.C(n_71),
.D(n_66),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_145),
.B(n_148),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_146),
.A2(n_166),
.B1(n_170),
.B2(n_94),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_161),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_104),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_152),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_107),
.A2(n_27),
.B1(n_18),
.B2(n_45),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_164),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_96),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_154),
.B(n_158),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_64),
.C(n_50),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_188),
.C(n_191),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_63),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_113),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_63),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_142),
.Y(n_165)
);

BUFx8_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_103),
.A2(n_18),
.B1(n_45),
.B2(n_2),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_187),
.B1(n_144),
.B2(n_134),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_0),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_184),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_170)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_121),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_189),
.Y(n_196)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_95),
.B1(n_123),
.B2(n_143),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_7),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_192),
.Y(n_208)
);

AO22x2_ASAP7_75t_L g186 ( 
.A1(n_103),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_186)
);

FAx1_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_190),
.CI(n_135),
.CON(n_222),
.SN(n_222)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_103),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_124),
.B(n_11),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_107),
.A2(n_116),
.B(n_115),
.C(n_127),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_101),
.A2(n_132),
.B(n_133),
.C(n_105),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_94),
.B(n_143),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_123),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_101),
.B(n_105),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_109),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_229),
.B1(n_165),
.B2(n_153),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_186),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_223),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_163),
.B(n_192),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_125),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_216),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_129),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_129),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_219),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_151),
.A2(n_102),
.B1(n_114),
.B2(n_97),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_163),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_148),
.B(n_114),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_166),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_144),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_230),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_102),
.B1(n_97),
.B2(n_135),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_135),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_168),
.C(n_162),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_150),
.C(n_181),
.Y(n_257)
);

AOI32xp33_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_189),
.A3(n_160),
.B1(n_172),
.B2(n_193),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_164),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_236),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_164),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_237),
.B(n_265),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_242),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_156),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_264),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_214),
.B(n_188),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_199),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_246),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_188),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_251),
.B(n_257),
.C(n_258),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_220),
.Y(n_252)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_216),
.B(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_194),
.B1(n_203),
.B2(n_238),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_205),
.B(n_149),
.C(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_174),
.B(n_186),
.C(n_171),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_222),
.B(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_196),
.B(n_150),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_176),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_269),
.B(n_213),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_209),
.B(n_159),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_273),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_196),
.B(n_159),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_207),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_245),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_296),
.C(n_306),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_224),
.B1(n_222),
.B2(n_226),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_276),
.A2(n_308),
.B1(n_294),
.B2(n_287),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_250),
.A2(n_270),
.B1(n_273),
.B2(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_300),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_201),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_264),
.C(n_200),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_250),
.A2(n_259),
.B(n_267),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_307),
.B(n_308),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_254),
.A2(n_226),
.B1(n_202),
.B2(n_234),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_246),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_248),
.A2(n_203),
.B(n_236),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_261),
.A2(n_224),
.B(n_230),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_237),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_310),
.B(n_314),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_284),
.B(n_257),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_251),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_323),
.C(n_327),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_336),
.B1(n_286),
.B2(n_283),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_307),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_SL g358 ( 
.A(n_317),
.B(n_271),
.C(n_272),
.Y(n_358)
);

NAND5xp2_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_249),
.C(n_223),
.D(n_227),
.E(n_253),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_318),
.A2(n_299),
.B1(n_300),
.B2(n_298),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_288),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_322),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_249),
.Y(n_320)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_263),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_244),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_332),
.C(n_335),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_285),
.A2(n_247),
.B(n_256),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_330),
.A2(n_285),
.B(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_331),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_243),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_291),
.B(n_208),
.Y(n_333)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_242),
.C(n_240),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_206),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_315),
.B(n_279),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_349),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_348),
.B1(n_352),
.B2(n_354),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_298),
.C(n_203),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_359),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_341),
.A2(n_351),
.B(n_330),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_313),
.A2(n_194),
.B1(n_298),
.B2(n_203),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_332),
.B(n_289),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_295),
.C(n_289),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_355),
.C(n_325),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_305),
.B(n_295),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_260),
.B1(n_262),
.B2(n_286),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_278),
.C(n_281),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_309),
.A2(n_281),
.B1(n_278),
.B2(n_301),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_356),
.A2(n_342),
.B1(n_312),
.B2(n_331),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_301),
.Y(n_357)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_319),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_335),
.B(n_255),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_362),
.B(n_366),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_312),
.Y(n_363)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_375),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_346),
.C(n_355),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_229),
.C(n_207),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_344),
.Y(n_366)
);

AO21x1_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_380),
.B(n_199),
.Y(n_387)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_372),
.A2(n_378),
.B1(n_370),
.B2(n_363),
.Y(n_393)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_376),
.Y(n_389)
);

OAI322xp33_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_320),
.A3(n_318),
.B1(n_309),
.B2(n_326),
.C1(n_334),
.C2(n_328),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_374),
.B(n_379),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_326),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_356),
.A2(n_339),
.B1(n_351),
.B2(n_341),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_378),
.A2(n_311),
.B1(n_297),
.B2(n_324),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_199),
.C(n_297),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_369),
.A2(n_338),
.B1(n_345),
.B2(n_353),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_384),
.B1(n_385),
.B2(n_393),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_380),
.A2(n_359),
.B(n_349),
.Y(n_383)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_343),
.B1(n_340),
.B2(n_311),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_372),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_266),
.B(n_239),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_390),
.A2(n_371),
.B(n_252),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_364),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_399),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_398),
.Y(n_412)
);

NOR2x1_ASAP7_75t_R g399 ( 
.A(n_393),
.B(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_400),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_401),
.B(n_405),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_365),
.C(n_375),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_391),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_386),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_406),
.Y(n_414)
);

OAI221xp5_ASAP7_75t_L g405 ( 
.A1(n_381),
.A2(n_358),
.B1(n_377),
.B2(n_371),
.C(n_252),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_388),
.A2(n_377),
.B(n_302),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_395),
.B(n_290),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_407),
.B(n_394),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_382),
.B1(n_392),
.B2(n_391),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_408),
.B(n_390),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_413),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_384),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_387),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_416),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_411),
.A2(n_401),
.B(n_398),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_418),
.A2(n_411),
.B(n_412),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_399),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_421),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_397),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_232),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_420),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_426),
.B(n_428),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_417),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_429),
.C(n_228),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_232),
.Y(n_429)
);

AOI221xp5_ASAP7_75t_L g430 ( 
.A1(n_425),
.A2(n_228),
.B1(n_218),
.B2(n_210),
.C(n_179),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_430),
.A2(n_426),
.B(n_157),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_432),
.Y(n_434)
);

OAI31xp33_ASAP7_75t_L g435 ( 
.A1(n_433),
.A2(n_431),
.A3(n_155),
.B(n_182),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_434),
.Y(n_436)
);


endmodule