module real_aes_17799_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_733;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g112 ( .A(n_0), .B(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_1), .A2(n_4), .B1(n_281), .B2(n_282), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_2), .A2(n_44), .B1(n_182), .B2(n_230), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_3), .A2(n_25), .B1(n_230), .B2(n_264), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_5), .A2(n_17), .B1(n_531), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_6), .A2(n_62), .B1(n_167), .B2(n_168), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_7), .A2(n_18), .B1(n_182), .B2(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_9), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_10), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_11), .A2(n_19), .B1(n_532), .B2(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_12), .A2(n_66), .B1(n_140), .B2(n_141), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
BUFx2_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
OR2x2_ASAP7_75t_L g130 ( .A(n_13), .B(n_39), .Y(n_130) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_14), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_15), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_16), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_20), .A2(n_99), .B1(n_282), .B2(n_531), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_21), .A2(n_40), .B1(n_160), .B2(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_22), .B(n_158), .Y(n_592) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_23), .A2(n_60), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_24), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_26), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_27), .B(n_155), .Y(n_222) );
INVx4_ASAP7_75t_R g206 ( .A(n_28), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_29), .A2(n_48), .B1(n_186), .B2(n_279), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_30), .A2(n_55), .B1(n_186), .B2(n_531), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_31), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_32), .B(n_556), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_33), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_34), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g286 ( .A(n_35), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_SL g261 ( .A1(n_36), .A2(n_154), .B(n_182), .C(n_262), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_37), .A2(n_56), .B1(n_182), .B2(n_186), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_38), .Y(n_809) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_41), .A2(n_87), .B1(n_182), .B2(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g827 ( .A1(n_42), .A2(n_54), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g829 ( .A(n_42), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_43), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_45), .A2(n_47), .B1(n_182), .B2(n_183), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_46), .A2(n_61), .B1(n_531), .B2(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g226 ( .A(n_49), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_50), .B(n_182), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_51), .Y(n_240) );
INVx2_ASAP7_75t_L g135 ( .A(n_52), .Y(n_135) );
BUFx3_ASAP7_75t_L g116 ( .A(n_53), .Y(n_116) );
INVx1_ASAP7_75t_L g128 ( .A(n_53), .Y(n_128) );
INVx1_ASAP7_75t_L g828 ( .A(n_54), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_57), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_58), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_59), .A2(n_88), .B1(n_182), .B2(n_186), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_63), .A2(n_76), .B1(n_279), .B2(n_548), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_64), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_65), .A2(n_79), .B1(n_182), .B2(n_183), .Y(n_533) );
INVx1_ASAP7_75t_L g141 ( .A(n_66), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_67), .A2(n_98), .B1(n_531), .B2(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g173 ( .A(n_68), .Y(n_173) );
AND2x4_ASAP7_75t_L g176 ( .A(n_69), .B(n_177), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_70), .A2(n_90), .B1(n_186), .B2(n_279), .Y(n_278) );
AO22x1_ASAP7_75t_L g156 ( .A1(n_71), .A2(n_77), .B1(n_157), .B2(n_160), .Y(n_156) );
INVx1_ASAP7_75t_L g177 ( .A(n_72), .Y(n_177) );
AND2x2_ASAP7_75t_L g265 ( .A(n_73), .B(n_218), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_74), .B(n_167), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_75), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_78), .B(n_230), .Y(n_241) );
INVx2_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_81), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_82), .B(n_218), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_83), .A2(n_97), .B1(n_167), .B2(n_186), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_84), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_85), .B(n_171), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_86), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_89), .B(n_218), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_91), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_92), .B(n_218), .Y(n_237) );
INVx1_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_93), .B(n_127), .Y(n_126) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_94), .B(n_158), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_95), .A2(n_167), .B(n_188), .C(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g211 ( .A(n_96), .B(n_212), .Y(n_211) );
NAND2xp33_ASAP7_75t_L g245 ( .A(n_100), .B(n_207), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_117), .B(n_830), .Y(n_101) );
BUFx4f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx8_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx8_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_105), .B(n_831), .Y(n_830) );
AND2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_110), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
NOR3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_114), .C(n_116), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g503 ( .A(n_115), .Y(n_503) );
INVx1_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
NOR2x1_ASAP7_75t_L g815 ( .A(n_116), .B(n_130), .Y(n_815) );
NAND2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_816), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_131), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_120), .A2(n_822), .B(n_824), .Y(n_821) );
NOR2x1_ASAP7_75t_R g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx4_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx3_ASAP7_75t_L g823 ( .A(n_123), .Y(n_823) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
CKINVDCx8_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_SL g125 ( .A(n_126), .B(n_129), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_129), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_138), .B(n_808), .Y(n_131) );
BUFx12f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_SL g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_135), .B(n_813), .Y(n_812) );
INVx3_ASAP7_75t_L g820 ( .A(n_135), .Y(n_820) );
OAI22xp33_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_142), .B1(n_143), .B2(n_807), .Y(n_138) );
INVx1_ASAP7_75t_L g807 ( .A(n_139), .Y(n_807) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI22x1_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_501), .B1(n_504), .B2(n_806), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_411), .Y(n_145) );
NOR3xp33_ASAP7_75t_L g146 ( .A(n_147), .B(n_340), .C(n_382), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_314), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_213), .B1(n_289), .B2(n_300), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_194), .Y(n_150) );
AOI21xp33_ASAP7_75t_L g333 ( .A1(n_151), .A2(n_334), .B(n_336), .Y(n_333) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_151), .A2(n_407), .B(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_178), .Y(n_151) );
INVx2_ASAP7_75t_L g326 ( .A(n_152), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_152), .B(n_179), .Y(n_356) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_162), .C(n_174), .Y(n_153) );
INVx6_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_154), .A2(n_245), .B(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_154), .B(n_156), .Y(n_298) );
O2A1O1Ixp5_ASAP7_75t_L g590 ( .A1(n_154), .A2(n_183), .B(n_591), .C(n_592), .Y(n_590) );
BUFx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g165 ( .A(n_155), .Y(n_165) );
INVx1_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
INVx1_ASAP7_75t_L g225 ( .A(n_155), .Y(n_225) );
INVxp67_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g531 ( .A(n_158), .Y(n_531) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g161 ( .A(n_159), .Y(n_161) );
INVx1_ASAP7_75t_L g167 ( .A(n_159), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_159), .Y(n_169) );
INVx3_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_159), .Y(n_230) );
INVx1_ASAP7_75t_L g258 ( .A(n_159), .Y(n_258) );
INVx2_ASAP7_75t_L g264 ( .A(n_159), .Y(n_264) );
OAI21xp33_ASAP7_75t_SL g221 ( .A1(n_160), .A2(n_222), .B(n_223), .Y(n_221) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g297 ( .A(n_162), .Y(n_297) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_170), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_163), .A2(n_228), .B(n_229), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_163), .A2(n_184), .B1(n_269), .B2(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g514 ( .A(n_164), .Y(n_514) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g243 ( .A(n_165), .Y(n_243) );
INVx1_ASAP7_75t_L g576 ( .A(n_168), .Y(n_576) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_169), .B(n_203), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g174 ( .A1(n_170), .A2(n_171), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g189 ( .A(n_171), .Y(n_189) );
INVx2_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
INVx2_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
INVx1_ASAP7_75t_L g299 ( .A(n_174), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_175), .A2(n_254), .B(n_261), .Y(n_253) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx10_ASAP7_75t_L g190 ( .A(n_176), .Y(n_190) );
BUFx10_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
INVx1_ASAP7_75t_L g284 ( .A(n_176), .Y(n_284) );
AND2x2_ASAP7_75t_L g396 ( .A(n_178), .B(n_235), .Y(n_396) );
INVx1_ASAP7_75t_L g429 ( .A(n_178), .Y(n_429) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g291 ( .A(n_179), .B(n_236), .Y(n_291) );
AND2x2_ASAP7_75t_L g322 ( .A(n_179), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g331 ( .A(n_179), .Y(n_331) );
OR2x2_ASAP7_75t_L g350 ( .A(n_179), .B(n_196), .Y(n_350) );
AND2x2_ASAP7_75t_L g365 ( .A(n_179), .B(n_196), .Y(n_365) );
AO31x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_189), .A3(n_190), .B(n_191), .Y(n_179) );
OAI22x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B1(n_185), .B2(n_187), .Y(n_180) );
INVx4_ASAP7_75t_L g183 ( .A(n_182), .Y(n_183) );
INVx1_ASAP7_75t_L g532 ( .A(n_182), .Y(n_532) );
INVx1_ASAP7_75t_L g548 ( .A(n_182), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_183), .A2(n_240), .B(n_241), .C(n_242), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_184), .A2(n_187), .B1(n_278), .B2(n_280), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_184), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_184), .A2(n_187), .B1(n_522), .B2(n_524), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_184), .A2(n_530), .B1(n_533), .B2(n_534), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_184), .A2(n_514), .B1(n_546), .B2(n_547), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_184), .A2(n_514), .B1(n_555), .B2(n_557), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_184), .A2(n_514), .B1(n_565), .B2(n_566), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_184), .A2(n_534), .B1(n_575), .B2(n_577), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_184), .A2(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_186), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g281 ( .A(n_186), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_187), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_SL g534 ( .A(n_188), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_189), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_189), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g210 ( .A(n_190), .Y(n_210) );
AO31x2_ASAP7_75t_L g511 ( .A1(n_190), .A2(n_271), .A3(n_512), .B(n_516), .Y(n_511) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_190), .A2(n_520), .A3(n_554), .B(n_559), .Y(n_553) );
AO31x2_ASAP7_75t_L g573 ( .A1(n_190), .A2(n_252), .A3(n_574), .B(n_578), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx2_ASAP7_75t_L g212 ( .A(n_193), .Y(n_212) );
BUFx2_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_193), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_193), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_195), .B(n_364), .Y(n_407) );
OR2x2_ASAP7_75t_L g495 ( .A(n_195), .B(n_356), .Y(n_495) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g323 ( .A(n_196), .Y(n_323) );
AND2x2_ASAP7_75t_L g332 ( .A(n_196), .B(n_295), .Y(n_332) );
AND2x2_ASAP7_75t_L g335 ( .A(n_196), .B(n_236), .Y(n_335) );
AND2x2_ASAP7_75t_L g354 ( .A(n_196), .B(n_235), .Y(n_354) );
AND2x4_ASAP7_75t_L g373 ( .A(n_196), .B(n_296), .Y(n_373) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_200), .B(n_211), .Y(n_196) );
AO31x2_ASAP7_75t_L g544 ( .A1(n_197), .A2(n_535), .A3(n_545), .B(n_549), .Y(n_544) );
AO31x2_ASAP7_75t_L g563 ( .A1(n_197), .A2(n_283), .A3(n_564), .B(n_567), .Y(n_563) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_199), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_SL g578 ( .A(n_199), .B(n_579), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_204), .B(n_210), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_205) );
INVx2_ASAP7_75t_L g279 ( .A(n_207), .Y(n_279) );
INVx1_ASAP7_75t_L g556 ( .A(n_207), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_208), .Y(n_558) );
INVx1_ASAP7_75t_L g535 ( .A(n_210), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_233), .B(n_274), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_214), .B(n_368), .Y(n_471) );
CKINVDCx14_ASAP7_75t_R g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_216), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g304 ( .A(n_216), .Y(n_304) );
OR2x2_ASAP7_75t_L g312 ( .A(n_216), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_216), .B(n_305), .Y(n_337) );
AND2x2_ASAP7_75t_L g362 ( .A(n_216), .B(n_276), .Y(n_362) );
AND2x2_ASAP7_75t_L g380 ( .A(n_216), .B(n_310), .Y(n_380) );
INVx1_ASAP7_75t_L g419 ( .A(n_216), .Y(n_419) );
AND2x2_ASAP7_75t_L g421 ( .A(n_216), .B(n_422), .Y(n_421) );
NAND2x1p5_ASAP7_75t_SL g440 ( .A(n_216), .B(n_361), .Y(n_440) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_220), .Y(n_216) );
NOR2x1_ASAP7_75t_L g247 ( .A(n_218), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g271 ( .A(n_218), .Y(n_271) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g231 ( .A(n_219), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_219), .B(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g520 ( .A(n_219), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_219), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_219), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_SL g588 ( .A(n_219), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_227), .B(n_231), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
BUFx4f_ASAP7_75t_L g260 ( .A(n_225), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_230), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_232), .A2(n_268), .A3(n_271), .B(n_272), .Y(n_267) );
OAI32xp33_ASAP7_75t_L g324 ( .A1(n_233), .A2(n_316), .A3(n_325), .B1(n_327), .B2(n_329), .Y(n_324) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_249), .Y(n_233) );
INVx1_ASAP7_75t_L g364 ( .A(n_234), .Y(n_364) );
AND2x2_ASAP7_75t_L g372 ( .A(n_234), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g371 ( .A(n_235), .B(n_295), .Y(n_371) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx3_ASAP7_75t_L g321 ( .A(n_236), .Y(n_321) );
AND2x2_ASAP7_75t_L g330 ( .A(n_236), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g436 ( .A(n_236), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_244), .B(n_247), .Y(n_238) );
INVx2_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g306 ( .A(n_249), .Y(n_306) );
OR2x2_ASAP7_75t_L g316 ( .A(n_249), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g438 ( .A(n_249), .Y(n_438) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_266), .Y(n_249) );
AND2x2_ASAP7_75t_L g339 ( .A(n_250), .B(n_267), .Y(n_339) );
INVx2_ASAP7_75t_L g361 ( .A(n_250), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_250), .B(n_276), .Y(n_381) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g288 ( .A(n_251), .Y(n_288) );
AOI21x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_265), .Y(n_251) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_252), .A2(n_277), .A3(n_283), .B(n_285), .Y(n_276) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_252), .A2(n_529), .A3(n_535), .B(n_536), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_257), .B(n_260), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_SL g523 ( .A(n_264), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_266), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g370 ( .A(n_266), .Y(n_370) );
INVx2_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
BUFx2_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
OR2x2_ASAP7_75t_L g376 ( .A(n_267), .B(n_276), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_267), .B(n_276), .Y(n_409) );
INVx2_ASAP7_75t_L g357 ( .A(n_274), .Y(n_357) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_287), .Y(n_274) );
OR2x2_ASAP7_75t_L g344 ( .A(n_275), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g422 ( .A(n_275), .Y(n_422) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
INVx1_ASAP7_75t_L g313 ( .A(n_276), .Y(n_313) );
INVx1_ASAP7_75t_L g328 ( .A(n_276), .Y(n_328) );
AO31x2_ASAP7_75t_L g519 ( .A1(n_283), .A2(n_520), .A3(n_521), .B(n_525), .Y(n_519) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_SL g596 ( .A(n_284), .Y(n_596) );
OR2x2_ASAP7_75t_L g432 ( .A(n_287), .B(n_409), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_288), .B(n_304), .Y(n_345) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_288), .Y(n_347) );
OR2x2_ASAP7_75t_L g446 ( .A(n_288), .B(n_370), .Y(n_446) );
INVxp67_ASAP7_75t_L g470 ( .A(n_288), .Y(n_470) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2x1_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_291), .B(n_332), .Y(n_399) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g348 ( .A(n_293), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g461 ( .A(n_294), .Y(n_461) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g490 ( .A(n_295), .B(n_323), .Y(n_490) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g416 ( .A(n_296), .B(n_323), .Y(n_416) );
AOI21x1_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_307), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_303), .B(n_339), .Y(n_453) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx2_ASAP7_75t_L g317 ( .A(n_304), .Y(n_317) );
AND2x2_ASAP7_75t_L g367 ( .A(n_304), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_304), .B(n_361), .Y(n_410) );
OR2x2_ASAP7_75t_L g482 ( .A(n_304), .B(n_369), .Y(n_482) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g402 ( .A(n_308), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx2_ASAP7_75t_L g393 ( .A(n_309), .Y(n_393) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g383 ( .A(n_312), .B(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_312), .Y(n_394) );
OR2x2_ASAP7_75t_L g445 ( .A(n_312), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g500 ( .A(n_312), .Y(n_500) );
AOI211xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_324), .C(n_333), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g389 ( .A(n_317), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_317), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g462 ( .A(n_317), .B(n_339), .Y(n_462) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_320), .B(n_365), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_320), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g472 ( .A(n_320), .B(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g415 ( .A(n_321), .Y(n_415) );
AND2x2_ASAP7_75t_L g443 ( .A(n_322), .B(n_371), .Y(n_443) );
INVx2_ASAP7_75t_L g466 ( .A(n_322), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_322), .B(n_364), .Y(n_498) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_325), .B(n_330), .Y(n_452) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g405 ( .A(n_326), .B(n_331), .Y(n_405) );
OR2x2_ASAP7_75t_L g457 ( .A(n_326), .B(n_350), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_327), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_327), .B(n_339), .Y(n_493) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g441 ( .A(n_328), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_L g424 ( .A(n_330), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_330), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g474 ( .A(n_331), .Y(n_474) );
BUFx2_ASAP7_75t_L g342 ( .A(n_332), .Y(n_342) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g460 ( .A(n_335), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_339), .Y(n_401) );
NAND3xp33_ASAP7_75t_SL g340 ( .A(n_341), .B(n_351), .C(n_366), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_343), .B1(n_346), .B2(n_348), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_348), .A2(n_374), .B1(n_455), .B2(n_458), .C1(n_460), .C2(n_462), .Y(n_454) );
AND2x2_ASAP7_75t_L g486 ( .A(n_349), .B(n_435), .Y(n_486) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g434 ( .A(n_350), .B(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_357), .B1(n_358), .B2(n_363), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx2_ASAP7_75t_SL g430 ( .A(n_354), .Y(n_430) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
AND2x2_ASAP7_75t_L g417 ( .A(n_359), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g375 ( .A(n_360), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g369 ( .A(n_361), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g484 ( .A(n_362), .Y(n_484) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_365), .B(n_461), .Y(n_480) );
INVx1_ASAP7_75t_L g497 ( .A(n_365), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_372), .B2(n_374), .C1(n_377), .C2(n_378), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_373), .Y(n_377) );
AND2x2_ASAP7_75t_L g395 ( .A(n_373), .B(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g426 ( .A(n_373), .Y(n_426) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
OR2x2_ASAP7_75t_L g459 ( .A(n_376), .B(n_440), .Y(n_459) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B(n_388), .C(n_397), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_395), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_389), .A2(n_427), .B1(n_476), .B2(n_479), .C(n_481), .Y(n_475) );
AND2x4_ASAP7_75t_L g418 ( .A(n_390), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g449 ( .A(n_396), .Y(n_449) );
AOI211x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_402), .C(n_406), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g467 ( .A(n_405), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_408), .B(n_456), .C(n_457), .Y(n_455) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g491 ( .A(n_409), .Y(n_491) );
NOR2x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_463), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_413), .B(n_420), .C(n_442), .D(n_454), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AND2x2_ASAP7_75t_L g473 ( .A(n_416), .B(n_474), .Y(n_473) );
AOI221x1_ASAP7_75t_L g442 ( .A1(n_418), .A2(n_443), .B1(n_444), .B2(n_447), .C(n_450), .Y(n_442) );
AND2x2_ASAP7_75t_L g468 ( .A(n_418), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g478 ( .A(n_419), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_427), .B2(n_431), .C(n_433), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_425), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_430), .A2(n_434), .B1(n_437), .B2(n_439), .Y(n_433) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_434), .A2(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g456 ( .A(n_436), .Y(n_456) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_459), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .C(n_487), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B1(n_471), .B2(n_472), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g483 ( .A(n_470), .B(n_484), .Y(n_483) );
NAND2x1_ASAP7_75t_L g499 ( .A(n_470), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_485), .Y(n_481) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B1(n_492), .B2(n_494), .C(n_496), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
INVx4_ASAP7_75t_L g806 ( .A(n_501), .Y(n_806) );
BUFx12f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g814 ( .A(n_503), .B(n_815), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g826 ( .A(n_504), .B(n_827), .Y(n_826) );
NOR2x1p5_ASAP7_75t_L g504 ( .A(n_505), .B(n_716), .Y(n_504) );
NAND4xp75_ASAP7_75t_L g505 ( .A(n_506), .B(n_661), .C(n_681), .D(n_697), .Y(n_505) );
NOR2x1p5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_631), .Y(n_506) );
NAND4xp75_ASAP7_75t_L g507 ( .A(n_508), .B(n_569), .C(n_608), .D(n_617), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_538), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .Y(n_509) );
AND2x4_ASAP7_75t_L g741 ( .A(n_510), .B(n_668), .Y(n_741) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_511), .Y(n_584) );
INVx2_ASAP7_75t_L g602 ( .A(n_511), .Y(n_602) );
AND2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_587), .Y(n_625) );
OR2x2_ASAP7_75t_L g680 ( .A(n_511), .B(n_519), .Y(n_680) );
AND2x2_ASAP7_75t_L g598 ( .A(n_518), .B(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g748 ( .A(n_518), .B(n_625), .Y(n_748) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
OR2x2_ASAP7_75t_L g585 ( .A(n_519), .B(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g616 ( .A(n_519), .Y(n_616) );
AND2x2_ASAP7_75t_L g622 ( .A(n_519), .B(n_528), .Y(n_622) );
INVx1_ASAP7_75t_L g640 ( .A(n_519), .Y(n_640) );
INVx2_ASAP7_75t_L g669 ( .A(n_519), .Y(n_669) );
INVx3_ASAP7_75t_L g645 ( .A(n_527), .Y(n_645) );
INVx2_ASAP7_75t_L g650 ( .A(n_527), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_527), .B(n_601), .Y(n_655) );
AND2x2_ASAP7_75t_L g678 ( .A(n_527), .B(n_657), .Y(n_678) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_527), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_527), .B(n_733), .Y(n_732) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g667 ( .A(n_528), .Y(n_667) );
AND2x2_ASAP7_75t_L g715 ( .A(n_528), .B(n_669), .Y(n_715) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_551), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_540), .B(n_659), .Y(n_706) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2x1p5_ASAP7_75t_L g703 ( .A(n_541), .B(n_659), .Y(n_703) );
INVx1_ASAP7_75t_L g804 ( .A(n_541), .Y(n_804) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g754 ( .A(n_542), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
OR2x2_ASAP7_75t_L g688 ( .A(n_543), .B(n_562), .Y(n_688) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g630 ( .A(n_544), .Y(n_630) );
AND2x4_ASAP7_75t_L g636 ( .A(n_544), .B(n_637), .Y(n_636) );
AOI32xp33_ASAP7_75t_L g774 ( .A1(n_551), .A2(n_677), .A3(n_775), .B1(n_777), .B2(n_778), .Y(n_774) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g723 ( .A(n_552), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_553), .Y(n_571) );
OR2x2_ASAP7_75t_L g605 ( .A(n_553), .B(n_563), .Y(n_605) );
INVx1_ASAP7_75t_L g620 ( .A(n_553), .Y(n_620) );
AND2x2_ASAP7_75t_L g629 ( .A(n_553), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g635 ( .A(n_553), .Y(n_635) );
INVx2_ASAP7_75t_L g660 ( .A(n_553), .Y(n_660) );
AND2x2_ASAP7_75t_L g779 ( .A(n_553), .B(n_573), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_561), .B(n_612), .Y(n_699) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_563), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g628 ( .A(n_563), .Y(n_628) );
INVx2_ASAP7_75t_L g637 ( .A(n_563), .Y(n_637) );
AND2x4_ASAP7_75t_L g659 ( .A(n_563), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_563), .Y(n_751) );
AOI22x1_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_580), .B1(n_598), .B2(n_603), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_572), .B(n_729), .C(n_730), .D(n_731), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_572), .B(n_629), .Y(n_759) );
INVx4_ASAP7_75t_SL g612 ( .A(n_573), .Y(n_612) );
BUFx2_ASAP7_75t_L g675 ( .A(n_573), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_573), .B(n_620), .Y(n_738) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g700 ( .A(n_582), .B(n_649), .Y(n_700) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g623 ( .A(n_586), .B(n_601), .Y(n_623) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_587), .B(n_602), .Y(n_647) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_597), .Y(n_587) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_588), .A2(n_589), .B(n_597), .Y(n_642) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .B(n_596), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_599), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g665 ( .A(n_599), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g704 ( .A(n_600), .B(n_622), .Y(n_704) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g747 ( .A(n_602), .B(n_657), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_603), .A2(n_720), .B1(n_722), .B2(n_725), .C(n_727), .Y(n_719) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx2_ASAP7_75t_L g613 ( .A(n_605), .Y(n_613) );
OR2x2_ASAP7_75t_L g713 ( .A(n_605), .B(n_652), .Y(n_713) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_614), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_609), .A2(n_735), .B1(n_739), .B2(n_742), .Y(n_734) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
AND2x4_ASAP7_75t_L g658 ( .A(n_610), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g770 ( .A(n_610), .B(n_688), .Y(n_770) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g618 ( .A(n_612), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g634 ( .A(n_612), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g693 ( .A(n_612), .B(n_630), .Y(n_693) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_612), .Y(n_710) );
INVx1_ASAP7_75t_L g724 ( .A(n_612), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_612), .B(n_637), .Y(n_767) );
AND2x4_ASAP7_75t_L g674 ( .A(n_613), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g672 ( .A(n_615), .Y(n_672) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_616), .B(n_657), .Y(n_656) );
NAND2x1_ASAP7_75t_L g776 ( .A(n_616), .B(n_678), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B1(n_624), .B2(n_626), .Y(n_617) );
AND2x2_ASAP7_75t_L g643 ( .A(n_618), .B(n_636), .Y(n_643) );
INVx1_ASAP7_75t_L g684 ( .A(n_618), .Y(n_684) );
AND2x2_ASAP7_75t_L g791 ( .A(n_618), .B(n_652), .Y(n_791) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_SL g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g624 ( .A(n_622), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g764 ( .A(n_622), .Y(n_764) );
AND2x2_ASAP7_75t_L g781 ( .A(n_622), .B(n_641), .Y(n_781) );
AND2x2_ASAP7_75t_L g797 ( .A(n_622), .B(n_747), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_623), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g720 ( .A(n_623), .B(n_721), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_623), .A2(n_713), .B1(n_728), .B2(n_732), .Y(n_727) );
INVx1_ASAP7_75t_L g683 ( .A(n_625), .Y(n_683) );
AND2x2_ASAP7_75t_L g714 ( .A(n_625), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_625), .B(n_721), .Y(n_743) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g749 ( .A(n_629), .B(n_750), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_629), .A2(n_653), .B1(n_758), .B2(n_760), .Y(n_757) );
INVx3_ASAP7_75t_L g652 ( .A(n_630), .Y(n_652) );
AND2x2_ASAP7_75t_L g784 ( .A(n_630), .B(n_637), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_648), .Y(n_631) );
AOI32xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_638), .A3(n_641), .B1(n_643), .B2(n_644), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_635), .Y(n_730) );
INVx1_ASAP7_75t_L g755 ( .A(n_635), .Y(n_755) );
INVx3_ASAP7_75t_L g711 ( .A(n_636), .Y(n_711) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g786 ( .A1(n_639), .A2(n_787), .B1(n_788), .B2(n_789), .C(n_790), .Y(n_786) );
BUFx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g763 ( .A(n_641), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g799 ( .A(n_641), .B(n_760), .Y(n_799) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g657 ( .A(n_642), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_644), .B(n_672), .Y(n_671) );
AO22x1_ASAP7_75t_L g701 ( .A1(n_644), .A2(n_702), .B1(n_704), .B2(n_705), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g805 ( .A(n_644), .B(n_672), .Y(n_805) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx2_ASAP7_75t_L g721 ( .A(n_645), .Y(n_721) );
INVx1_ASAP7_75t_L g731 ( .A(n_645), .Y(n_731) );
AND2x2_ASAP7_75t_L g651 ( .A(n_646), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_SL g733 ( .A(n_647), .Y(n_733) );
INVx1_ASAP7_75t_L g773 ( .A(n_647), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B(n_653), .C(n_658), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2x1p5_ASAP7_75t_L g760 ( .A(n_650), .B(n_680), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_651), .B(n_710), .Y(n_787) );
AOI31xp33_ASAP7_75t_L g670 ( .A1(n_652), .A2(n_671), .A3(n_673), .B(n_676), .Y(n_670) );
INVx4_ASAP7_75t_L g729 ( .A(n_652), .Y(n_729) );
OR2x2_ASAP7_75t_L g766 ( .A(n_652), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AND2x4_ASAP7_75t_L g668 ( .A(n_657), .B(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_659), .Y(n_664) );
AND2x2_ASAP7_75t_L g695 ( .A(n_659), .B(n_693), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g661 ( .A(n_662), .B(n_670), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g788 ( .A(n_665), .Y(n_788) );
INVx1_ASAP7_75t_L g696 ( .A(n_666), .Y(n_696) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g726 ( .A(n_667), .Y(n_726) );
AND2x2_ASAP7_75t_L g725 ( .A(n_668), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .A3(n_685), .B1(n_689), .B2(n_692), .C1(n_694), .C2(n_696), .Y(n_682) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI211x1_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B(n_701), .C(n_707), .Y(n_697) );
INVx1_ASAP7_75t_L g802 ( .A(n_698), .Y(n_802) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g756 ( .A(n_700), .Y(n_756) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OA21x2_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_712), .B(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx2_ASAP7_75t_L g777 ( .A(n_711), .Y(n_777) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp33_ASAP7_75t_L g772 ( .A(n_715), .B(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_785), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_752), .C(n_768), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_734), .C(n_744), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_721), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI21xp33_ASAP7_75t_L g780 ( .A1(n_725), .A2(n_781), .B(n_782), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_729), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_729), .B(n_779), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_730), .B(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_731), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g790 ( .A1(n_741), .A2(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_749), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B(n_757), .C(n_761), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_SL g771 ( .A(n_763), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_767), .Y(n_789) );
OAI211xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B(n_774), .C(n_780), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_779), .B(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g800 ( .A(n_779), .Y(n_800) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g796 ( .A(n_784), .Y(n_796) );
NOR3xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_794), .C(n_801), .Y(n_785) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI21xp33_ASAP7_75t_SL g794 ( .A1(n_795), .A2(n_798), .B(n_800), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AOI21xp33_ASAP7_75t_R g801 ( .A1(n_802), .A2(n_803), .B(n_805), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx6_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
BUFx10_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OR2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_821), .Y(n_816) );
INVxp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
endmodule