module real_jpeg_27958_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_181;
wire n_85;
wire n_102;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_0),
.B(n_215),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_3),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_118),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_118),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_3),
.A2(n_51),
.B1(n_53),
.B2(n_118),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_5),
.A2(n_45),
.B1(n_49),
.B2(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_5),
.A2(n_51),
.B1(n_53),
.B2(n_69),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_29),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_45),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_6),
.B(n_20),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_45),
.B(n_64),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_6),
.A2(n_48),
.B(n_51),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_6),
.B(n_66),
.Y(n_210)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_10),
.A2(n_31),
.B1(n_45),
.B2(n_49),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_31),
.B1(n_51),
.B2(n_53),
.Y(n_103)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_11),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_126),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_124),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_94),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_15),
.B(n_94),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_15),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_73),
.CI(n_81),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_38),
.B2(n_39),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_19),
.B(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_20),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_22),
.B(n_29),
.C(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_21),
.A2(n_34),
.B(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_21),
.B(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_23),
.B(n_26),
.Y(n_157)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_24),
.A2(n_61),
.B(n_62),
.C(n_66),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_24),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_24),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_24),
.A2(n_57),
.B(n_61),
.C(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_28),
.B(n_34),
.Y(n_259)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_33),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_35),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_36),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_37),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_40),
.B(n_139),
.C(n_141),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_40),
.A2(n_41),
.B1(n_141),
.B2(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_54),
.B(n_55),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_42),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_43),
.B(n_56),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_43),
.B(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_49),
.B1(n_61),
.B2(n_64),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_45),
.A2(n_47),
.B(n_57),
.C(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_50),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_53),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_79),
.B(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_54),
.B(n_57),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_57),
.B(n_88),
.Y(n_230)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_67),
.B(n_70),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_60),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_60),
.B(n_144),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_60),
.Y(n_262)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_66),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_71),
.B(n_154),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_75),
.A2(n_152),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_78),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_79),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_93),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_83),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_85),
.B1(n_93),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_84),
.A2(n_85),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_85),
.B(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_86),
.B(n_89),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_86),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_103),
.Y(n_135)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_90),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_92),
.B(n_197),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_119),
.C(n_120),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_95),
.A2(n_96),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.C(n_110),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_97),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_105),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_98),
.B(n_105),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_99),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_100),
.A2(n_134),
.B(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_101),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_119),
.B(n_120),
.Y(n_283)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_279),
.B(n_284),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_266),
.B(n_278),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_174),
.B(n_248),
.C(n_265),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_162),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_130),
.B(n_162),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_145),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_132),
.B(n_138),
.C(n_145),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_133),
.B(n_136),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_137),
.B(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_140),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_147),
.B(n_150),
.C(n_155),
.Y(n_263)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_163),
.A2(n_164),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_173),
.B(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_247),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_240),
.B(n_246),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_199),
.B(n_239),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_189),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_178),
.B(n_189),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_185),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_179),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_237)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_196),
.C(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_234),
.B(n_238),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_216),
.B(n_233),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_232),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_227),
.B(n_231),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_225),
.B(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_250),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_263),
.B2(n_264),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.C(n_264),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_258),
.C(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_275),
.C(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);


endmodule