module real_jpeg_7066_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_12;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_42),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_2),
.A2(n_42),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_42),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_126),
.C(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_222),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_2),
.A2(n_229),
.B(n_231),
.C(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_2),
.B(n_243),
.C(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_133),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_2),
.B(n_75),
.Y(n_269)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_4),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_6),
.A2(n_69),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_6),
.A2(n_69),
.B1(n_160),
.B2(n_164),
.Y(n_159)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_9),
.A2(n_35),
.B1(n_67),
.B2(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_171),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_169),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_151),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_14),
.B(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_98),
.C(n_135),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_15),
.B(n_98),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_71),
.B2(n_72),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_16),
.A2(n_74),
.B(n_97),
.Y(n_168)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_36),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_18),
.A2(n_73),
.B1(n_74),
.B2(n_97),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_18),
.A2(n_36),
.B1(n_97),
.B2(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_27),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_20),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_22),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_23),
.A2(n_27),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_23),
.A2(n_139),
.B1(n_186),
.B2(n_192),
.Y(n_185)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_25),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_28),
.Y(n_141)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_30),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_30),
.Y(n_191)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_33),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_46),
.B1(n_54),
.B2(n_63),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_38),
.B(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_40),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_42),
.A2(n_70),
.B(n_114),
.Y(n_231)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_46),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_46),
.B(n_54),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_46),
.A2(n_54),
.B(n_131),
.Y(n_156)
);

NAND2x1_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_54),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_50),
.Y(n_244)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_55),
.B(n_253),
.Y(n_252)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_64),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_128)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_73),
.A2(n_74),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_73),
.A2(n_100),
.B(n_150),
.C(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_73),
.A2(n_74),
.B1(n_225),
.B2(n_236),
.Y(n_280)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_74),
.B(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_74),
.B(n_99),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_74),
.B(n_100),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_74),
.B(n_146),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_85),
.B(n_94),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_86),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_81),
.Y(n_234)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_127),
.B(n_134),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_99),
.A2(n_100),
.B1(n_146),
.B2(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_99),
.A2(n_100),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_99),
.A2(n_146),
.B(n_227),
.C(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_99),
.B(n_146),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_99),
.B(n_212),
.C(n_268),
.Y(n_283)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_128),
.Y(n_134)
);

AO21x2_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_113),
.B(n_123),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_102)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_123),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

OA22x2_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

FAx1_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_152),
.CI(n_168),
.CON(n_151),
.SN(n_151)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_135),
.A2(n_136),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_148),
.B(n_149),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_146),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_146),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_146),
.A2(n_201),
.B1(n_221),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_146),
.A2(n_201),
.B1(n_240),
.B2(n_241),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_146),
.A2(n_201),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_146),
.A2(n_185),
.B1(n_201),
.B2(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_149),
.B(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AND3x1_ASAP7_75t_L g298 ( 
.A(n_150),
.B(n_275),
.C(n_299),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_151),
.Y(n_311)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_167),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI211xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_215),
.B(n_305),
.C(n_310),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_197),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_175),
.A2(n_197),
.B(n_306),
.C(n_309),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_194),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_176),
.B(n_194),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_183),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_184),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_178),
.A2(n_179),
.B1(n_204),
.B2(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_185),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_213),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_198),
.B(n_213),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.C(n_203),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_199),
.B(n_200),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_221),
.C(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_265),
.C(n_272),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_203),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_223),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_212),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_223),
.B1(n_228),
.B2(n_235),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_212),
.A2(n_223),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_212),
.B(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_287),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_277),
.B(n_286),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_263),
.B(n_276),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_237),
.B(n_262),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_223),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_236),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_249),
.B(n_261),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_246),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_259),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_273),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_273),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_297),
.C(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_300),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_303),
.Y(n_308)
);


endmodule