module fake_jpeg_13521_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_1),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_18),
.B1(n_15),
.B2(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_19),
.B1(n_17),
.B2(n_10),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_18),
.B1(n_15),
.B2(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_26),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_12),
.B1(n_16),
.B2(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_17),
.B1(n_33),
.B2(n_23),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_32),
.B(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_16),
.C(n_4),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_47),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_19),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_34),
.B1(n_31),
.B2(n_28),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_47),
.Y(n_62)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_21),
.B1(n_25),
.B2(n_23),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_58),
.B(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_29),
.B1(n_21),
.B2(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_65),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_44),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.C(n_64),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_42),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_9),
.A3(n_7),
.B1(n_6),
.B2(n_53),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_56),
.B(n_57),
.C(n_48),
.D(n_52),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_41),
.C(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_73),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_60),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_35),
.C(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_56),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_75),
.B(n_63),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_7),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_6),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_81),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_71),
.C(n_35),
.Y(n_84)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_71),
.B1(n_72),
.B2(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_78),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_76),
.Y(n_88)
);

OAI31xp33_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_80),
.A3(n_2),
.B(n_4),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_4),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_89),
.Y(n_93)
);


endmodule