module real_jpeg_21593_n_17 (n_8, n_0, n_2, n_10, n_9, n_79, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_81, n_1, n_80, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_79;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_81;
input n_1;
input n_80;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_12),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_2),
.B(n_80),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_81),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_45),
.B1(n_48),
.B2(n_59),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_8),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_11),
.B(n_79),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_25),
.C(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_12),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_19),
.B1(n_20),
.B2(n_43),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_14),
.A2(n_43),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

AOI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_44),
.B1(n_60),
.B2(n_72),
.C(n_77),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_41),
.Y(n_20)
);

OAI211xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B(n_27),
.C(n_37),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_26),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_26),
.A2(n_37),
.B(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B(n_32),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_29),
.B(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_30),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_57),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.C(n_71),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);


endmodule