module real_jpeg_886_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_1),
.B(n_58),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_1),
.B(n_83),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_1),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_1),
.A2(n_58),
.B(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_1),
.B(n_27),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_1),
.A2(n_36),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_1),
.B(n_45),
.C(n_48),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_221),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_1),
.B(n_101),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_43),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_65),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_65),
.Y(n_188)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_34),
.B1(n_36),
.B2(n_70),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_5),
.A2(n_45),
.B1(n_49),
.B2(n_70),
.Y(n_212)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_9),
.A2(n_38),
.B1(n_58),
.B2(n_59),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_9),
.A2(n_38),
.B1(n_45),
.B2(n_49),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_34),
.B1(n_36),
.B2(n_67),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_67),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_45),
.B1(n_49),
.B2(n_67),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_11),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_111),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_111),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_11),
.A2(n_45),
.B1(n_49),
.B2(n_111),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_12),
.A2(n_34),
.B1(n_36),
.B2(n_150),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_150),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_12),
.A2(n_45),
.B1(n_49),
.B2(n_150),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_13),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_176),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_176),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_13),
.A2(n_45),
.B1(n_49),
.B2(n_176),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_15),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_15),
.A2(n_34),
.B1(n_36),
.B2(n_195),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_15),
.A2(n_45),
.B1(n_49),
.B2(n_195),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_16),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_16),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.C(n_71),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_22),
.A2(n_68),
.B1(n_119),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_22),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_53),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_25),
.B(n_42),
.C(n_54),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_25)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_26),
.A2(n_39),
.B1(n_116),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_26),
.A2(n_39),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_26),
.A2(n_39),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_26),
.A2(n_39),
.B1(n_191),
.B2(n_207),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_26),
.A2(n_39),
.B1(n_206),
.B2(n_253),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_27),
.A2(n_74),
.B(n_79),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_27),
.A2(n_73),
.B1(n_74),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_27),
.A2(n_74),
.B1(n_146),
.B2(n_173),
.Y(n_172)
);

AO22x2_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_28),
.B(n_32),
.Y(n_222)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_29),
.A2(n_31),
.A3(n_36),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_29),
.B(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_34),
.B(n_61),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_34),
.B(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_36),
.A2(n_59),
.A3(n_62),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_68),
.C(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_42),
.A2(n_53),
.B1(n_72),
.B2(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_50),
.B(n_52),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_43),
.A2(n_50),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_43),
.A2(n_50),
.B1(n_52),
.B2(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_43),
.A2(n_50),
.B1(n_106),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_43),
.A2(n_50),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_43),
.A2(n_50),
.B1(n_217),
.B2(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_43),
.A2(n_50),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_43),
.A2(n_50),
.B1(n_244),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_44),
.A2(n_143),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_44),
.A2(n_169),
.B1(n_216),
.B2(n_256),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_45),
.B(n_272),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_50),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_63),
.B1(n_69),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_63),
.B1(n_110),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_55),
.A2(n_63),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_55),
.A2(n_63),
.B1(n_194),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_56),
.A2(n_83),
.B1(n_149),
.B2(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_156),
.B(n_311),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_151),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_125),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_93),
.B(n_125),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_112),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_118),
.C(n_123),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_108),
.B(n_109),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_96),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_108),
.B1(n_109),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_98),
.A2(n_100),
.B1(n_139),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_98),
.A2(n_100),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_98),
.A2(n_100),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_101),
.B1(n_103),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_99),
.A2(n_101),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_99),
.A2(n_101),
.B1(n_188),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_99),
.A2(n_101),
.B1(n_225),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_99),
.A2(n_101),
.B1(n_221),
.B2(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_99),
.A2(n_101),
.B1(n_274),
.B2(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_118),
.B1(n_123),
.B2(n_124),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_114),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_133),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.C(n_147),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_135),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_147),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_151),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_152),
.B(n_155),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_177),
.B(n_310),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_158),
.B(n_160),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.C(n_174),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_167),
.B(n_170),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_174),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_200),
.B(n_309),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_198),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_179),
.B(n_198),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_197),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_180),
.B(n_197),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_182),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.C(n_193),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_183),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_187),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_190),
.B(n_193),
.Y(n_300)
);

AOI31xp33_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_294),
.A3(n_303),
.B(n_306),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_239),
.B(n_293),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_227),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_203),
.B(n_227),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.C(n_218),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_204),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_209),
.C(n_213),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_214),
.B(n_218),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_223),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_227),
.B(n_304),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.CI(n_230),
.CON(n_227),
.SN(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_231),
.B(n_234),
.C(n_238),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_288),
.B(n_292),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_257),
.B(n_287),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_246),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_252),
.C(n_255),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_268),
.B(n_286),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_280),
.B(n_285),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B(n_279),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_284),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);


endmodule