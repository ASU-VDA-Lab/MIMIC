module fake_jpeg_23447_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_1),
.CON(n_31),
.SN(n_31)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_14),
.Y(n_48)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_17),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_39),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_44),
.B1(n_15),
.B2(n_28),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_20),
.B1(n_18),
.B2(n_14),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_39),
.B1(n_30),
.B2(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_34),
.B(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_65),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_34),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_70),
.B1(n_76),
.B2(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_43),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

NOR2xp67_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_81),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_63),
.C(n_61),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.C(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_76),
.B1(n_67),
.B2(n_66),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_54),
.C(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_90),
.C(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_79),
.B1(n_80),
.B2(n_71),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_9),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_85),
.C(n_90),
.Y(n_95)
);

AO221x1_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_73),
.B1(n_51),
.B2(n_9),
.C(n_8),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_4),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.C(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_97),
.B(n_92),
.C(n_91),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_98),
.B(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_55),
.Y(n_102)
);


endmodule