module fake_jpeg_3808_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_22),
.B1(n_16),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_56),
.B1(n_37),
.B2(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_59),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_31),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_58),
.B1(n_38),
.B2(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_31),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_62),
.B1(n_53),
.B2(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_33),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_78),
.B1(n_63),
.B2(n_50),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_38),
.B1(n_26),
.B2(n_28),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_38),
.B1(n_17),
.B2(n_18),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_87),
.B1(n_43),
.B2(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_28),
.B1(n_26),
.B2(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_44),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_62),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_36),
.B1(n_39),
.B2(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_94),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_55),
.B1(n_43),
.B2(n_42),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_105),
.B1(n_108),
.B2(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_96),
.B1(n_74),
.B2(n_82),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_63),
.C(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_103),
.Y(n_113)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_63),
.B(n_62),
.C(n_60),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_76),
.B(n_79),
.Y(n_122)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_63),
.C(n_39),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_36),
.B1(n_50),
.B2(n_46),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_110),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_124),
.Y(n_157)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_115),
.Y(n_138)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_81),
.B1(n_86),
.B2(n_72),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_126),
.B1(n_65),
.B2(n_104),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_126),
.B1(n_97),
.B2(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_122),
.B1(n_135),
.B2(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_133),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_101),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_84),
.B1(n_86),
.B2(n_80),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_67),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_110),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_84),
.B1(n_78),
.B2(n_67),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_142),
.Y(n_165)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_144),
.B1(n_156),
.B2(n_77),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_125),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_145),
.B(n_32),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_101),
.B(n_94),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_127),
.B(n_120),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_152),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_94),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_63),
.C(n_32),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_155),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_153),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_103),
.B(n_65),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_117),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_122),
.B1(n_130),
.B2(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_159),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_114),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_91),
.B1(n_99),
.B2(n_105),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_83),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_167),
.B1(n_182),
.B2(n_161),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_151),
.C(n_147),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_87),
.B1(n_131),
.B2(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_46),
.B1(n_36),
.B2(n_49),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_87),
.C(n_39),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_183),
.C(n_188),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_175),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_82),
.B1(n_106),
.B2(n_46),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_39),
.C(n_106),
.Y(n_183)
);

AND2x4_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_32),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_145),
.B(n_162),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_187),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_39),
.Y(n_188)
);

INVx5_ASAP7_75t_SL g189 ( 
.A(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_190),
.B(n_200),
.C(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_199),
.B1(n_211),
.B2(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_198),
.B(n_174),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_143),
.A3(n_154),
.B1(n_152),
.B2(n_137),
.C1(n_159),
.C2(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_188),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_173),
.B1(n_186),
.B2(n_176),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_184),
.B(n_168),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_128),
.B1(n_98),
.B2(n_71),
.Y(n_199)
);

NOR4xp25_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_14),
.C(n_13),
.D(n_12),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_23),
.C(n_25),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_23),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_164),
.A2(n_15),
.B1(n_20),
.B2(n_29),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_128),
.C(n_64),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_163),
.C(n_172),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_29),
.B1(n_25),
.B2(n_21),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_208),
.C(n_209),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_228),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_189),
.B(n_170),
.C(n_178),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_231),
.B1(n_235),
.B2(n_29),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_23),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_207),
.B1(n_209),
.B2(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_23),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_234),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_210),
.B1(n_211),
.B2(n_193),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_14),
.B(n_13),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_214),
.B1(n_213),
.B2(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_0),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_250),
.C(n_255),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_201),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_244),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_20),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_229),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_177),
.C(n_64),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_217),
.B1(n_219),
.B2(n_223),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_29),
.C(n_25),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_21),
.C(n_20),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_219),
.C(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_259),
.A2(n_243),
.B1(n_253),
.B2(n_238),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_219),
.B(n_233),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_14),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_21),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_266),
.Y(n_277)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_21),
.B(n_20),
.C(n_15),
.D(n_12),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_15),
.C(n_1),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.C(n_256),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_0),
.C(n_1),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_254),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_275),
.B(n_283),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_282),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_246),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_270),
.C(n_260),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_241),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_238),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_240),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_279),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_293),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_292),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_270),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_295),
.B(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_276),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_257),
.A3(n_272),
.B1(n_273),
.B2(n_267),
.C1(n_5),
.C2(n_6),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_257),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_4),
.B(n_6),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_289),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_304),
.B(n_299),
.Y(n_311)
);

NAND4xp25_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_287),
.C(n_275),
.D(n_4),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_6),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_290),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.C(n_8),
.Y(n_313)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_301),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_305),
.C2(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_9),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_316),
.B(n_314),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_10),
.Y(n_318)
);


endmodule