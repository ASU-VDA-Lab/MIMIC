module fake_jpeg_12371_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_41),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_4),
.B(n_5),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_40),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_47),
.B1(n_44),
.B2(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_72),
.B1(n_78),
.B2(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_44),
.B1(n_5),
.B2(n_6),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_13),
.B(n_14),
.Y(n_83)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_10),
.B(n_12),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_80),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_76),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_88),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_90)
);

AOI211xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_92),
.B(n_29),
.C(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_27),
.Y(n_92)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_102),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_100),
.C(n_97),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_92),
.CI(n_95),
.CON(n_106),
.SN(n_106)
);

NOR2xp67_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_99),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

NAND2x1_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_104),
.Y(n_110)
);


endmodule