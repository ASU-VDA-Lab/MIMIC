module fake_jpeg_3001_n_641 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_641);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_641;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_587;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_7),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_84),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_65),
.Y(n_129)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_19),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g172 ( 
.A(n_74),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_24),
.B(n_8),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_86),
.Y(n_192)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_91),
.A2(n_26),
.B1(n_47),
.B2(n_44),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_18),
.B(n_17),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_102),
.A2(n_19),
.B(n_11),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_60),
.B(n_18),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_118),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_48),
.B(n_17),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_127),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_124),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_19),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_25),
.Y(n_126)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_61),
.Y(n_161)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_65),
.B(n_38),
.CON(n_130),
.SN(n_130)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_130),
.Y(n_276)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_73),
.B(n_38),
.CON(n_134),
.SN(n_134)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_134),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_23),
.B1(n_52),
.B2(n_37),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_137),
.A2(n_140),
.B1(n_148),
.B2(n_166),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_55),
.B1(n_52),
.B2(n_37),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_90),
.B(n_26),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_143),
.B(n_195),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_145),
.B(n_163),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_77),
.A2(n_29),
.B1(n_54),
.B2(n_53),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_146),
.A2(n_137),
.B1(n_208),
.B2(n_166),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_52),
.B1(n_54),
.B2(n_53),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_151),
.A2(n_181),
.B1(n_193),
.B2(n_200),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_29),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_125),
.A2(n_23),
.B1(n_47),
.B2(n_44),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_23),
.B1(n_40),
.B2(n_34),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_185),
.B1(n_188),
.B2(n_123),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_46),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_178),
.B(n_183),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_97),
.A2(n_46),
.B1(n_50),
.B2(n_34),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_50),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_63),
.A2(n_40),
.B1(n_36),
.B2(n_43),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_184),
.A2(n_208),
.B1(n_80),
.B2(n_75),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_78),
.A2(n_61),
.B1(n_35),
.B2(n_43),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_79),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_114),
.A2(n_45),
.B1(n_32),
.B2(n_27),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_87),
.B(n_11),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_143),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_67),
.A2(n_32),
.B1(n_27),
.B2(n_45),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_71),
.A2(n_32),
.B1(n_27),
.B2(n_45),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_213),
.Y(n_348)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_214),
.Y(n_319)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_215),
.Y(n_316)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_216),
.Y(n_327)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_218),
.A2(n_271),
.B1(n_201),
.B2(n_176),
.Y(n_320)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_167),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_220),
.B(n_247),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_221),
.Y(n_338)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_222),
.Y(n_290)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_224),
.Y(n_339)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_225),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_136),
.B(n_70),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_226),
.Y(n_307)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_240),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_110),
.C(n_113),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_234),
.B(n_269),
.C(n_226),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_235),
.B(n_248),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_139),
.Y(n_236)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_236),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_237),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_136),
.A2(n_93),
.B1(n_111),
.B2(n_108),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_238),
.B(n_244),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_239),
.Y(n_325)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_241),
.B(n_242),
.Y(n_299)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_246),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_144),
.A2(n_86),
.B1(n_106),
.B2(n_105),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_129),
.A2(n_122),
.B1(n_66),
.B2(n_99),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_245),
.A2(n_251),
.B1(n_261),
.B2(n_262),
.Y(n_335)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_130),
.B(n_45),
.CI(n_27),
.CON(n_248),
.SN(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_172),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_255),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_129),
.A2(n_100),
.B1(n_95),
.B2(n_83),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_172),
.B(n_82),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_252),
.B(n_273),
.Y(n_324)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

INVx13_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_254),
.A2(n_177),
.B1(n_202),
.B2(n_192),
.Y(n_292)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_154),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_260),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_159),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_258),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_153),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_259),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_164),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_134),
.A2(n_32),
.B1(n_27),
.B2(n_45),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_158),
.A2(n_20),
.B1(n_17),
.B2(n_16),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_142),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_263),
.B(n_266),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_158),
.A2(n_20),
.B1(n_12),
.B2(n_11),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_184),
.A2(n_20),
.B1(n_12),
.B2(n_9),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_147),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_131),
.B(n_0),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_196),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_270),
.B(n_281),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_200),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_162),
.B(n_0),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_274),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_277),
.A2(n_287),
.B1(n_4),
.B2(n_5),
.Y(n_337)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_198),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_286),
.B(n_210),
.Y(n_322)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_164),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_206),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_283),
.Y(n_298)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_285),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_138),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_175),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_292),
.A2(n_294),
.B1(n_303),
.B2(n_309),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_149),
.B1(n_212),
.B2(n_205),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_235),
.B(n_165),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_329),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_212),
.B1(n_177),
.B2(n_202),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_217),
.A2(n_185),
.B(n_188),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_306),
.A2(n_347),
.B(n_228),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_160),
.B1(n_176),
.B2(n_201),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_308),
.A2(n_255),
.B1(n_285),
.B2(n_259),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_170),
.B1(n_192),
.B2(n_191),
.Y(n_309)
);

AO22x1_ASAP7_75t_SL g315 ( 
.A1(n_254),
.A2(n_170),
.B1(n_156),
.B2(n_191),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_320),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_234),
.B(n_269),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_341),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_322),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_275),
.A2(n_169),
.B1(n_203),
.B2(n_150),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_333),
.B1(n_340),
.B2(n_344),
.Y(n_350)
);

AO22x1_ASAP7_75t_SL g332 ( 
.A1(n_217),
.A2(n_169),
.B1(n_150),
.B2(n_203),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_337),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_232),
.A2(n_190),
.B1(n_210),
.B2(n_152),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_217),
.B(n_190),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_219),
.C(n_266),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_223),
.A2(n_284),
.B1(n_253),
.B2(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_269),
.B(n_4),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_248),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_223),
.B(n_4),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_247),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_248),
.A2(n_6),
.B1(n_226),
.B2(n_244),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_346),
.A2(n_344),
.B1(n_291),
.B2(n_317),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_272),
.A2(n_6),
.B(n_249),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_328),
.A2(n_238),
.B1(n_280),
.B2(n_224),
.Y(n_351)
);

AOI22x1_ASAP7_75t_L g425 ( 
.A1(n_351),
.A2(n_360),
.B1(n_371),
.B2(n_372),
.Y(n_425)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_353),
.A2(n_391),
.B1(n_290),
.B2(n_330),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_343),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_357),
.A2(n_335),
.B(n_290),
.Y(n_409)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_359),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_328),
.A2(n_282),
.B1(n_239),
.B2(n_236),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_278),
.C(n_241),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_369),
.C(n_375),
.Y(n_404)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_366),
.B(n_382),
.Y(n_402)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_302),
.B(n_318),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_289),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_384),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_328),
.A2(n_231),
.B1(n_229),
.B2(n_243),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_331),
.A2(n_233),
.B1(n_227),
.B2(n_242),
.Y(n_372)
);

AOI22x1_ASAP7_75t_SL g373 ( 
.A1(n_317),
.A2(n_308),
.B1(n_306),
.B2(n_332),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_373),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_311),
.B(n_213),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_263),
.C(n_246),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_346),
.A2(n_216),
.B1(n_214),
.B2(n_222),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_379),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_225),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_381),
.C(n_393),
.Y(n_430)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_274),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_291),
.A2(n_258),
.B1(n_292),
.B2(n_307),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_392),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_293),
.B(n_336),
.C(n_332),
.Y(n_381)
);

BUFx2_ASAP7_75t_SL g383 ( 
.A(n_342),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_383),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_289),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_297),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_385),
.B(n_386),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_347),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_324),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_387),
.B(n_390),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_388),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_316),
.B(n_300),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_389),
.B(n_395),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_288),
.B(n_314),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_332),
.A2(n_315),
.B1(n_337),
.B2(n_320),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_326),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_310),
.C(n_299),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_288),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_394),
.B(n_301),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_338),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_410),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_310),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_401),
.C(n_420),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_299),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_357),
.A2(n_304),
.B(n_326),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_405),
.A2(n_409),
.B(n_418),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_312),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_365),
.A2(n_315),
.B1(n_320),
.B2(n_323),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_413),
.A2(n_415),
.B1(n_422),
.B2(n_423),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_365),
.A2(n_315),
.B1(n_320),
.B2(n_323),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_390),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_417),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_382),
.A2(n_363),
.B(n_365),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_419),
.A2(n_375),
.B1(n_378),
.B2(n_364),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_295),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_361),
.A2(n_367),
.B1(n_373),
.B2(n_394),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_361),
.A2(n_325),
.B1(n_305),
.B2(n_321),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_432),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_393),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_435),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_361),
.A2(n_325),
.B1(n_305),
.B2(n_321),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_377),
.B(n_295),
.C(n_296),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_296),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_371),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_402),
.A2(n_358),
.B1(n_359),
.B2(n_363),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_437),
.A2(n_461),
.B1(n_462),
.B2(n_470),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_427),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_445),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_366),
.Y(n_440)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_440),
.Y(n_482)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_381),
.B(n_392),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_444),
.A2(n_452),
.B(n_455),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_370),
.Y(n_446)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_446),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_384),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_449),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_396),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_450),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_428),
.A2(n_387),
.B(n_388),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_453),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_417),
.A2(n_391),
.B1(n_356),
.B2(n_350),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_454),
.A2(n_464),
.B1(n_425),
.B2(n_431),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_428),
.A2(n_356),
.B(n_376),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_405),
.A2(n_380),
.B(n_351),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_457),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_424),
.B(n_355),
.Y(n_458)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_459),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_416),
.B(n_379),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_460),
.B(n_465),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_402),
.A2(n_350),
.B1(n_360),
.B2(n_349),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_435),
.A2(n_349),
.B1(n_372),
.B2(n_385),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_431),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_468),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_409),
.A2(n_431),
.B(n_419),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_399),
.C(n_429),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_406),
.A2(n_368),
.B1(n_312),
.B2(n_319),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_406),
.B(n_352),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_472),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_396),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_401),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_476),
.B(n_483),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_460),
.B(n_416),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_477),
.B(n_492),
.Y(n_526)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_444),
.B(n_422),
.CI(n_430),
.CON(n_481),
.SN(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g521 ( 
.A1(n_481),
.A2(n_447),
.B(n_448),
.C(n_440),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_430),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_500),
.C(n_458),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_404),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_494),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_436),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_493),
.A2(n_451),
.B1(n_464),
.B2(n_463),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_441),
.B(n_404),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_437),
.B(n_398),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_445),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_420),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_498),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_469),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_410),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_504),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_456),
.B(n_397),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_454),
.A2(n_425),
.B1(n_408),
.B2(n_412),
.Y(n_501)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_452),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_466),
.C(n_442),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_446),
.B(n_433),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_508),
.A2(n_510),
.B1(n_512),
.B2(n_531),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_451),
.B1(n_439),
.B2(n_455),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_474),
.B(n_436),
.Y(n_513)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_513),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_475),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_515),
.B(n_517),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_486),
.Y(n_516)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_480),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_474),
.Y(n_518)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_518),
.Y(n_546)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_475),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_520),
.B(n_523),
.Y(n_557)
);

AOI21xp33_ASAP7_75t_L g560 ( 
.A1(n_521),
.A2(n_527),
.B(n_532),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_530),
.Y(n_540)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_488),
.B(n_408),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_524),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_436),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_525),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_506),
.B(n_471),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_463),
.C(n_412),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_529),
.C(n_476),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_487),
.B(n_457),
.C(n_448),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_500),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_490),
.A2(n_465),
.B(n_438),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_491),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_533),
.A2(n_534),
.B1(n_535),
.B2(n_505),
.Y(n_561)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_490),
.A2(n_438),
.B(n_413),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_536),
.B(n_499),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_537),
.B(n_542),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_497),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_538),
.B(n_550),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_484),
.C(n_498),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_539),
.B(n_544),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_509),
.A2(n_495),
.B1(n_473),
.B2(n_482),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_526),
.B(n_504),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_508),
.A2(n_479),
.B1(n_461),
.B2(n_482),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_548),
.A2(n_552),
.B1(n_559),
.B2(n_535),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_511),
.B(n_503),
.C(n_479),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_549),
.B(n_554),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_480),
.Y(n_550)
);

FAx1_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_481),
.CI(n_491),
.CON(n_551),
.SN(n_551)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_551),
.A2(n_518),
.B1(n_513),
.B2(n_515),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_SL g552 ( 
.A(n_529),
.B(n_481),
.C(n_415),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_522),
.C(n_514),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_514),
.B(n_470),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_558),
.B(n_512),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_509),
.A2(n_468),
.B1(n_467),
.B2(n_459),
.Y(n_559)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_561),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_562),
.A2(n_567),
.B1(n_547),
.B2(n_553),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_528),
.C(n_536),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_564),
.C(n_574),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_519),
.C(n_532),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_568),
.B(n_462),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_555),
.A2(n_548),
.B1(n_517),
.B2(n_551),
.Y(n_569)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_569),
.Y(n_589)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_545),
.Y(n_572)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_537),
.B(n_519),
.C(n_520),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_533),
.C(n_525),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_577),
.C(n_579),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_551),
.A2(n_527),
.B1(n_516),
.B2(n_534),
.Y(n_576)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_576),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_542),
.B(n_478),
.C(n_450),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_543),
.A2(n_531),
.B1(n_523),
.B2(n_478),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_578),
.A2(n_546),
.B1(n_559),
.B2(n_545),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_450),
.C(n_434),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_538),
.B(n_434),
.C(n_414),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_581),
.B(n_582),
.C(n_432),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_539),
.B(n_400),
.C(n_472),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_583),
.B(n_586),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_578),
.B(n_556),
.Y(n_584)
);

OAI321xp33_ASAP7_75t_L g607 ( 
.A1(n_584),
.A2(n_588),
.A3(n_595),
.B1(n_586),
.B2(n_591),
.C(n_589),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_546),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_579),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_557),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_571),
.A2(n_557),
.B1(n_425),
.B2(n_560),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_592),
.B(n_596),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_566),
.B(n_573),
.C(n_574),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_593),
.A2(n_594),
.B(n_403),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_580),
.A2(n_552),
.B(n_541),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_558),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_565),
.B(n_549),
.Y(n_596)
);

NOR2x1_ASAP7_75t_L g597 ( 
.A(n_568),
.B(n_423),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_597),
.A2(n_584),
.B(n_587),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_598),
.B(n_600),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_565),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_605),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_563),
.C(n_582),
.Y(n_605)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_606),
.Y(n_620)
);

AOI21x1_ASAP7_75t_L g619 ( 
.A1(n_607),
.A2(n_613),
.B(n_614),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_L g608 ( 
.A1(n_588),
.A2(n_597),
.B(n_594),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_609),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_590),
.B(n_581),
.C(n_570),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_570),
.C(n_564),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_610),
.B(n_609),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_595),
.B(n_449),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_611),
.B(n_612),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_453),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_617),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_602),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_600),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_621),
.B(n_603),
.C(n_608),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_605),
.B(n_586),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_622),
.A2(n_623),
.B(n_319),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_583),
.C(n_598),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_625),
.B(n_327),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g626 ( 
.A(n_618),
.B(n_403),
.C(n_330),
.Y(n_626)
);

AO21x1_ASAP7_75t_L g632 ( 
.A1(n_626),
.A2(n_627),
.B(n_628),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_619),
.A2(n_615),
.B(n_617),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_620),
.A2(n_327),
.B(n_338),
.Y(n_630)
);

AO21x1_ASAP7_75t_L g633 ( 
.A1(n_630),
.A2(n_348),
.B(n_297),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_624),
.B(n_623),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_631),
.B(n_621),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_L g636 ( 
.A1(n_633),
.A2(n_629),
.B(n_301),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_634),
.B(n_635),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_636),
.A2(n_632),
.B(n_339),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_638),
.A2(n_637),
.B(n_339),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_313),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_640),
.A2(n_313),
.B(n_639),
.Y(n_641)
);


endmodule