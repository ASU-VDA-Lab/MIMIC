module real_jpeg_7579_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_1),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_1),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_99),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_1),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_1),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_1),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_1),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_2),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_2),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_2),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_2),
.Y(n_284)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_3),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_4),
.Y(n_202)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_5),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_5),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_5),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_5),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_5),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_5),
.B(n_399),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_5),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_6),
.Y(n_504)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_8),
.B(n_16),
.Y(n_346)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_9),
.Y(n_282)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_240),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_11),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_11),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_11),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_11),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_11),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_11),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_11),
.B(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_12),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_12),
.Y(n_240)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_13),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_14),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_14),
.B(n_37),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_14),
.B(n_42),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_14),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_14),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_14),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_14),
.B(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_15),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_16),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_16),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_16),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_16),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_16),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_17),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_17),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_17),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_17),
.B(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_499),
.B(n_501),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_74),
.B(n_111),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_21),
.B(n_74),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_21),
.Y(n_507)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_62),
.CI(n_63),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_45),
.C(n_51),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_23),
.A2(n_24),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_52),
.C(n_57),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_27),
.A2(n_28),
.B1(n_52),
.B2(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_27),
.A2(n_28),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_35),
.C(n_41),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_28),
.B(n_235),
.C(n_239),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_33),
.Y(n_376)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_34),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_36),
.B1(n_66),
.B2(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_36),
.B(n_185),
.C(n_188),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_36),
.B(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_39),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_40),
.A2(n_41),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_41),
.B(n_139),
.C(n_143),
.Y(n_168)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_51),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_70),
.C(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_52),
.A2(n_105),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_52),
.A2(n_105),
.B1(n_259),
.B2(n_260),
.Y(n_299)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_55),
.Y(n_302)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_55),
.Y(n_373)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_56),
.Y(n_242)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_56),
.Y(n_396)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_56),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_58),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_57),
.A2(n_58),
.B1(n_130),
.B2(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_58),
.B(n_128),
.C(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_70),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_66),
.B(n_198),
.C(n_203),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_66),
.A2(n_69),
.B1(n_159),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_66),
.A2(n_69),
.B1(n_203),
.B2(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_69),
.B(n_150),
.C(n_159),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_70),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_167)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_106),
.C(n_107),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_75),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_91),
.C(n_102),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_76),
.B(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_87),
.C(n_89),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_79),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_78),
.B(n_122),
.C(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_78),
.A2(n_79),
.B1(n_303),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_79),
.B(n_301),
.C(n_303),
.Y(n_300)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_81),
.B(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_81),
.Y(n_422)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_81),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_91),
.B(n_102),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.C(n_98),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_147),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_92),
.Y(n_147)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_95),
.A2(n_96),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_96),
.B(n_152),
.C(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_101),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_101),
.Y(n_341)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_105),
.B(n_259),
.C(n_264),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_106),
.B(n_107),
.Y(n_497)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AO21x1_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_494),
.B(n_498),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_249),
.B(n_491),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_213),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_115),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_172),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_116),
.B(n_172),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_163),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_117),
.B(n_164),
.C(n_170),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_145),
.C(n_148),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_118),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_133),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_119),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_124),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_128),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_124),
.B(n_236),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_124),
.A2(n_128),
.B1(n_235),
.B2(n_236),
.Y(n_458)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_125),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_126),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_129),
.B(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_139),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_139),
.B(n_227),
.Y(n_257)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_226),
.C(n_228),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_150),
.A2(n_151),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_157),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_152),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_152),
.A2(n_193),
.B1(n_199),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_152),
.A2(n_193),
.B1(n_412),
.B2(n_417),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_152),
.B(n_417),
.Y(n_459)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_154),
.Y(n_410)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_154),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_155),
.B(n_273),
.C(n_276),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_155),
.A2(n_195),
.B1(n_273),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_162),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_162),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_178),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_173),
.B(n_176),
.CI(n_178),
.CON(n_248),
.SN(n_248)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_197),
.C(n_209),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_191),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_180),
.B(n_184),
.Y(n_320)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_188),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_191),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_209),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_199),
.B(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_199),
.A2(n_224),
.B1(n_307),
.B2(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_201),
.Y(n_416)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_202),
.Y(n_407)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_207),
.Y(n_304)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_208),
.Y(n_402)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_248),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_214),
.B(n_248),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_215),
.B(n_217),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_219),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.C(n_245),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_220),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.C(n_231),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_225),
.B(n_231),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_245),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.C(n_243),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_234),
.B(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_239),
.Y(n_314)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_248),
.Y(n_508)
);

AOI221xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_384),
.B1(n_484),
.B2(n_489),
.C(n_490),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_324),
.C(n_328),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_251),
.A2(n_485),
.B(n_488),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_317),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_252),
.B(n_317),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_294),
.C(n_296),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_253),
.B(n_294),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_279),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_254),
.B(n_280),
.C(n_291),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_271),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_256),
.B(n_272),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_258),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_276),
.B(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_287),
.C(n_290),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_283),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_290),
.Y(n_316)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_311),
.C(n_315),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_305),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_300),
.A2(n_305),
.B1(n_306),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_301),
.B(n_361),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_321),
.C(n_323),
.Y(n_325)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_324),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_325),
.B(n_326),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_355),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_329),
.A2(n_486),
.B(n_487),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_353),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_330),
.B(n_353),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.C(n_351),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_351),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.C(n_342),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_337),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_421),
.Y(n_420)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.C(n_347),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_343),
.A2(n_344),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_345),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_382),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_356),
.B(n_382),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.C(n_379),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_357),
.B(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_359),
.B(n_379),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.C(n_377),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_360),
.B(n_475),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_363),
.A2(n_377),
.B1(n_378),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_363),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_369),
.C(n_374),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_364),
.A2(n_365),
.B1(n_374),
.B2(n_375),
.Y(n_463)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_369),
.B(n_463),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_479),
.B(n_483),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_465),
.B(n_478),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_452),
.B(n_464),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_428),
.B(n_451),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_418),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_418),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_403),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_390),
.B(n_404),
.C(n_411),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_397),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_391),
.B(n_398),
.C(n_400),
.Y(n_461)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_411),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_408),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_406),
.Y(n_440)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_412),
.Y(n_417)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.C(n_423),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_448),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_420),
.A2(n_423),
.B1(n_424),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_445),
.B(n_450),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_438),
.B(n_444),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_437),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_437),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_435),
.Y(n_446)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_436),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_441),
.Y(n_438)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_447),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_454),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_460),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_461),
.C(n_462),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_455),
.Y(n_506)
);

FAx1_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.CI(n_459),
.CON(n_455),
.SN(n_455)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_458),
.C(n_459),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_477),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_477),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_474),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_471),
.C(n_474),
.Y(n_480)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_472),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_481),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_496),
.Y(n_498)
);

INVx8_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);


endmodule