module fake_jpeg_22110_n_182 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_12),
.B1(n_14),
.B2(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_52),
.B1(n_58),
.B2(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_14),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_53),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_27),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_1),
.C(n_2),
.Y(n_77)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_25),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_20),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_1),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_76),
.B1(n_41),
.B2(n_65),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_27),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_72),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_17),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_74),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_17),
.B1(n_2),
.B2(n_4),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_92),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_61),
.Y(n_114)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_4),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_7),
.C(n_8),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_66),
.Y(n_93)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_60),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_7),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_92),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_101),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_110),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_70),
.B1(n_77),
.B2(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_50),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_53),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_55),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_48),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_98),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_70),
.B1(n_82),
.B2(n_79),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_131),
.B(n_132),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_68),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_115),
.C(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_95),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_133),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_92),
.B1(n_68),
.B2(n_40),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_54),
.B(n_57),
.C(n_59),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_115),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_133),
.C(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_142),
.B1(n_144),
.B2(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_132),
.B1(n_125),
.B2(n_118),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_86),
.B1(n_95),
.B2(n_140),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_152),
.C(n_155),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_127),
.C(n_119),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_162),
.B(n_163),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_143),
.A3(n_144),
.B1(n_100),
.B2(n_93),
.C1(n_96),
.C2(n_53),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_129),
.B1(n_116),
.B2(n_96),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_103),
.B1(n_54),
.B2(n_44),
.Y(n_163)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_100),
.A3(n_90),
.B1(n_57),
.B2(n_51),
.C(n_112),
.Y(n_164)
);

AOI31xp67_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_100),
.A3(n_150),
.B(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_155),
.C(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_163),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_101),
.B1(n_83),
.B2(n_112),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_165),
.C(n_10),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_175),
.Y(n_182)
);


endmodule