module fake_jpeg_7925_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_52),
.B1(n_58),
.B2(n_16),
.Y(n_93)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_16),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_30),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_69),
.B(n_73),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_68),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_71),
.C(n_80),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_20),
.B1(n_25),
.B2(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_43),
.C(n_37),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_23),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_83),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_32),
.B1(n_22),
.B2(n_17),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_32),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_37),
.CI(n_44),
.CON(n_110),
.SN(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_17),
.B1(n_58),
.B2(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_101),
.B1(n_34),
.B2(n_46),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_96),
.B1(n_98),
.B2(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_0),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_15),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_27),
.B1(n_21),
.B2(n_33),
.Y(n_104)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_37),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_107),
.B1(n_120),
.B2(n_128),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_104),
.A2(n_85),
.B1(n_125),
.B2(n_94),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_12),
.C(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_84),
.B1(n_80),
.B2(n_98),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_43),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_64),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_44),
.B1(n_36),
.B2(n_57),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_11),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_36),
.B1(n_34),
.B2(n_64),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_89),
.B(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_83),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_69),
.A2(n_34),
.B1(n_46),
.B2(n_15),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_73),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_118),
.B1(n_104),
.B2(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_134),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_139),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_141),
.B1(n_103),
.B2(n_107),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_143),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_89),
.C(n_90),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_133),
.C(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_91),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_101),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_81),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_152),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_153),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_81),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_99),
.B(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_14),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_146),
.B1(n_161),
.B2(n_147),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_0),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_160),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVxp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_123),
.Y(n_168)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_172),
.B1(n_175),
.B2(n_179),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_171),
.Y(n_198)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_170),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_115),
.B1(n_112),
.B2(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_181),
.B1(n_182),
.B2(n_176),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_86),
.B1(n_87),
.B2(n_94),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_94),
.B1(n_90),
.B2(n_88),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_180),
.B(n_183),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_88),
.B1(n_97),
.B2(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_95),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_186),
.B(n_190),
.Y(n_201)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_88),
.Y(n_190)
);

INVx5_ASAP7_75t_SL g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_75),
.A3(n_97),
.B1(n_10),
.B2(n_3),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_154),
.B(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_0),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_133),
.B(n_1),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_134),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_141),
.B(n_139),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_205),
.B(n_208),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_141),
.B1(n_160),
.B2(n_138),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_166),
.B1(n_188),
.B2(n_189),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_160),
.B1(n_157),
.B2(n_149),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_213),
.A2(n_193),
.B1(n_194),
.B2(n_190),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_152),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_222),
.C(n_171),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_165),
.B(n_158),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_221),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_170),
.B(n_158),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_167),
.B(n_152),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_233),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_244),
.B1(n_199),
.B2(n_210),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_192),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_215),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_183),
.C(n_168),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_239),
.C(n_247),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_172),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_184),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_251),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_243),
.B1(n_249),
.B2(n_209),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_193),
.B1(n_182),
.B2(n_160),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_202),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_212),
.A2(n_195),
.B1(n_179),
.B2(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_177),
.C(n_162),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_164),
.C(n_75),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_202),
.C(n_204),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_201),
.A2(n_75),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_201),
.B(n_1),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_233),
.C(n_238),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_208),
.B(n_210),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_240),
.B(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_246),
.B(n_206),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_224),
.CI(n_213),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_266),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_211),
.Y(n_286)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_209),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_248),
.B1(n_230),
.B2(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_274),
.C(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_239),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_286),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_2),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_255),
.C(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_258),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_289),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_253),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_282),
.Y(n_304)
);

FAx1_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_263),
.CI(n_278),
.CON(n_293),
.SN(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_265),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_260),
.C(n_4),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_252),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_264),
.B1(n_269),
.B2(n_252),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_301),
.B1(n_5),
.B2(n_6),
.Y(n_311)
);

AOI211xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_268),
.B(n_253),
.C(n_263),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_276),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_312),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_278),
.B1(n_265),
.B2(n_272),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_304),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_311),
.B1(n_297),
.B2(n_288),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_274),
.C(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_3),
.C(n_4),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_3),
.B(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_5),
.C(n_6),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_294),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.C(n_293),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_292),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_293),
.A3(n_301),
.B1(n_297),
.B2(n_6),
.C1(n_9),
.C2(n_7),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_319),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_302),
.B1(n_7),
.B2(n_9),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_314),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_7),
.Y(n_325)
);

OAI21x1_ASAP7_75t_SL g328 ( 
.A1(n_326),
.A2(n_316),
.B(n_318),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_327),
.B1(n_323),
.B2(n_9),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_323),
.B(n_7),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule