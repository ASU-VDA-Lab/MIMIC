module fake_netlist_6_4953_n_189 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_29, n_25, n_189);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_189;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_85;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_171;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVxp33_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_3),
.C(n_4),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_45),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_62),
.Y(n_77)
);

OAI221xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_44),
.B1(n_39),
.B2(n_48),
.C(n_43),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_48),
.B1(n_43),
.B2(n_41),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_44),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_41),
.B(n_40),
.C(n_51),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_40),
.B1(n_42),
.B2(n_10),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_58),
.B1(n_57),
.B2(n_72),
.Y(n_86)
);

OAI221xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_46),
.B1(n_38),
.B2(n_32),
.C(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_71),
.B1(n_70),
.B2(n_68),
.Y(n_94)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_61),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_71),
.B1(n_70),
.B2(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_86),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_64),
.B1(n_59),
.B2(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_81),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_100),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_86),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_73),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_75),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_96),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_78),
.C(n_109),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_95),
.B(n_92),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_95),
.B(n_91),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_101),
.B(n_95),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_79),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_109),
.B(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_108),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_114),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_112),
.B(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_80),
.C(n_109),
.D(n_98),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_108),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_116),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_130),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_132),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_135),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_127),
.B1(n_84),
.B2(n_85),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_84),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_80),
.B(n_125),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_137),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_85),
.B(n_84),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_136),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_136),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_85),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

BUFx4_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_154),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_133),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_146),
.C(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_143),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_153),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_61),
.Y(n_167)
);

NAND2x1p5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_157),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_59),
.B1(n_55),
.B2(n_54),
.C(n_157),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_54),
.A3(n_85),
.B1(n_79),
.B2(n_60),
.C1(n_15),
.C2(n_16),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_161),
.C(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_79),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_128),
.C(n_88),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_7),
.Y(n_175)
);

NAND4xp25_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_160),
.C(n_163),
.D(n_108),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_163),
.B1(n_79),
.B2(n_83),
.C(n_88),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_11),
.C(n_13),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_14),
.B(n_15),
.Y(n_180)
);

NAND4xp75_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_115),
.C(n_101),
.D(n_25),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_170),
.B1(n_115),
.B2(n_73),
.Y(n_183)
);

AO22x2_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_182),
.B1(n_181),
.B2(n_176),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_73),
.B1(n_107),
.B2(n_26),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_73),
.B1(n_19),
.B2(n_27),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_102),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_186),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_184),
.B1(n_187),
.B2(n_185),
.Y(n_189)
);


endmodule