module fake_jpeg_21267_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_47),
.B1(n_50),
.B2(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_42),
.B1(n_54),
.B2(n_49),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_55),
.B1(n_59),
.B2(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_79),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_74),
.B1(n_76),
.B2(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_46),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_53),
.B(n_61),
.C(n_58),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_85),
.B1(n_88),
.B2(n_5),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_94),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_45),
.B1(n_59),
.B2(n_52),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_71),
.B1(n_57),
.B2(n_45),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_4),
.B(n_5),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_2),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_48),
.C(n_51),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_48),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_7),
.C(n_8),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_103),
.B(n_16),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_12),
.Y(n_113)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_8),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_28),
.B1(n_39),
.B2(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_13),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_111),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_116),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_95),
.B(n_121),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_116),
.B(n_115),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_110),
.B(n_99),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_97),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_96),
.A3(n_102),
.B1(n_30),
.B2(n_31),
.C1(n_34),
.C2(n_23),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_24),
.Y(n_130)
);


endmodule