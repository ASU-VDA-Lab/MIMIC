module fake_jpeg_25158_n_279 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_22),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_13),
.B(n_26),
.C(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_36),
.B1(n_31),
.B2(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_22),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_65),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_29),
.B1(n_16),
.B2(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_29),
.B1(n_16),
.B2(n_34),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_73),
.B1(n_51),
.B2(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_23),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_70)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_50),
.B(n_30),
.Y(n_80)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_71),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_16),
.B1(n_27),
.B2(n_18),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_27),
.B1(n_14),
.B2(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

AO21x1_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_50),
.B(n_14),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_26),
.B(n_25),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_80),
.B(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_85),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_96),
.B1(n_85),
.B2(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_52),
.B1(n_13),
.B2(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_94),
.B1(n_71),
.B2(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_24),
.B1(n_69),
.B2(n_28),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_98),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_52),
.B1(n_13),
.B2(n_51),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_48),
.B(n_44),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_105),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_121),
.B1(n_108),
.B2(n_104),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_64),
.CI(n_61),
.CON(n_105),
.SN(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_109),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_73),
.B1(n_74),
.B2(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_117),
.B1(n_122),
.B2(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_110),
.B(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_84),
.B1(n_79),
.B2(n_92),
.Y(n_125)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_70),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_24),
.B(n_14),
.C(n_70),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_24),
.B(n_77),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_69),
.B1(n_54),
.B2(n_48),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_60),
.C(n_30),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_78),
.B1(n_80),
.B2(n_79),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_131),
.B1(n_145),
.B2(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_133),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_80),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_149),
.B(n_102),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_78),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_17),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_142),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_98),
.B(n_1),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_19),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_12),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_114),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_93),
.B1(n_77),
.B2(n_60),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_93),
.B1(n_28),
.B2(n_21),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_20),
.B(n_21),
.C(n_17),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_18),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_136),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_20),
.B(n_19),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_112),
.Y(n_150)
);

AO32x1_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_116),
.A3(n_102),
.B1(n_104),
.B2(n_19),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_162),
.B1(n_165),
.B2(n_172),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_158),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_147),
.B(n_149),
.Y(n_182)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_100),
.B1(n_17),
.B2(n_15),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_17),
.B1(n_15),
.B2(n_19),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_169),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_15),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_15),
.B1(n_12),
.B2(n_10),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_180),
.Y(n_192)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_12),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_10),
.C(n_9),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_9),
.C(n_1),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_10),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_142),
.B1(n_151),
.B2(n_126),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_162),
.B1(n_174),
.B2(n_173),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_135),
.B(n_124),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_198),
.B1(n_159),
.B2(n_165),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_196),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_134),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_0),
.Y(n_220)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_146),
.B(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_168),
.C(n_169),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_208),
.C(n_213),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_220),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_166),
.C(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_155),
.B1(n_159),
.B2(n_153),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_188),
.B1(n_201),
.B2(n_195),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_180),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_185),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_0),
.C(n_1),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_0),
.C(n_3),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_202),
.C(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_0),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_207),
.A2(n_189),
.B1(n_196),
.B2(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_231),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_230),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_192),
.C(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_234),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_199),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_208),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_244),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_212),
.C(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_243),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_231),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_217),
.B(n_210),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_232),
.B(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_220),
.C(n_213),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_228),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_192),
.B(n_4),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_242),
.B(n_239),
.C(n_237),
.D(n_244),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_3),
.B(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_224),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_246),
.A2(n_221),
.B1(n_227),
.B2(n_229),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_221),
.B1(n_235),
.B2(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_227),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_3),
.C(n_4),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_262),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_5),
.B(n_6),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_248),
.C(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_267),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_250),
.B(n_6),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_5),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_272),
.B(n_270),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_268),
.B(n_264),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

AO21x1_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_273),
.B(n_275),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_7),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_7),
.B1(n_8),
.B2(n_246),
.Y(n_279)
);


endmodule