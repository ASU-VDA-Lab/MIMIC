module real_jpeg_18533_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_0),
.A2(n_203),
.B1(n_206),
.B2(n_209),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_0),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_2),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_2),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_3),
.A2(n_139),
.B1(n_144),
.B2(n_146),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_3),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_3),
.A2(n_146),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_3),
.A2(n_146),
.B1(n_303),
.B2(n_305),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_4),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_5),
.A2(n_64),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_6),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_6),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_7),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_7),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_153),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_77),
.B1(n_80),
.B2(n_85),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_9),
.A2(n_85),
.B1(n_218),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_9),
.A2(n_85),
.B1(n_293),
.B2(n_297),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_9),
.A2(n_85),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_26),
.Y(n_25)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_11),
.A2(n_160),
.A3(n_162),
.B1(n_163),
.B2(n_169),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_11),
.A2(n_211),
.A3(n_217),
.B1(n_221),
.B2(n_225),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_11),
.A2(n_168),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_11),
.B(n_102),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_11),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_11),
.B(n_261),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_11),
.A2(n_168),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_13),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_53),
.B2(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_15),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_267),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_266),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_190),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_20),
.B(n_190),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_120),
.C(n_157),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_21),
.A2(n_22),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_75),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_24),
.B(n_75),
.C(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OR2x6_ASAP7_75t_L g234 ( 
.A(n_26),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_26),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_29),
.Y(n_236)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_32),
.Y(n_370)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_36),
.Y(n_174)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_36),
.Y(n_216)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_41),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_58),
.Y(n_41)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_42),
.Y(n_352)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_45),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_46),
.A2(n_179),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_68),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_59),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_63),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_132)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_63),
.Y(n_304)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_63),
.Y(n_346)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_68),
.A2(n_302),
.B(n_308),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_68),
.A2(n_168),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_68),
.A2(n_325),
.B1(n_338),
.B2(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_70),
.Y(n_340)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_71),
.Y(n_307)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_72),
.Y(n_277)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_86),
.B1(n_113),
.B2(n_114),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_76),
.A2(n_86),
.B1(n_113),
.B2(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_86),
.A2(n_113),
.B1(n_114),
.B2(n_253),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_102),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_93),
.Y(n_254)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_109),
.Y(n_102)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_104),
.Y(n_291)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_106),
.Y(n_316)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_118),
.A2(n_119),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_118),
.A2(n_119),
.B1(n_286),
.B2(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_120),
.B(n_158),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_137),
.B(n_147),
.Y(n_120)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_121),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_121),
.A2(n_261),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_121),
.A2(n_261),
.B1(n_292),
.B2(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_126),
.B1(n_128),
.B2(n_131),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_131),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_132),
.A2(n_138),
.B1(n_259),
.B2(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_133),
.Y(n_279)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_135),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_145),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_148),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_178),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_159),
.B(n_178),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_168),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_168),
.B(n_281),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_SL g290 ( 
.A1(n_168),
.A2(n_280),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B(n_184),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_179),
.A2(n_324),
.B1(n_329),
.B2(n_330),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_181),
.B(n_310),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_188),
.Y(n_312)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_232),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_201),
.Y(n_337)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_231),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_251),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_241),
.B1(n_247),
.B2(n_250),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_257),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_373),
.B(n_378),
.Y(n_268)
);

OAI21x1_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_357),
.B(n_372),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_321),
.B(n_356),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_300),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_272),
.B(n_300),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_288),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_273),
.A2(n_288),
.B1(n_289),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.A3(n_278),
.B1(n_280),
.B2(n_283),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_314),
.C(n_320),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_334),
.B(n_355),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_332),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_332),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_350),
.B(n_354),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_353),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_358),
.B(n_359),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_371),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_363),
.C(n_371),
.Y(n_374)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx6_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_374),
.B(n_375),
.Y(n_378)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_376),
.Y(n_377)
);


endmodule