module fake_netlist_1_8732_n_840 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_840);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_840;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_695;
wire n_650;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_8), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_79), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_84), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_102), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_100), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_0), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_80), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_39), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_66), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_28), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_4), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_27), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_9), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_52), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_72), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_104), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_71), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_36), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_31), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_43), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_23), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_63), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_46), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_103), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_54), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_97), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_93), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_12), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_17), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_57), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_75), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_92), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_62), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_16), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_67), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_68), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_59), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_113), .B(n_0), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_113), .B(n_1), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_146), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_109), .B(n_1), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_119), .B(n_2), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_109), .B(n_2), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_119), .B(n_3), .Y(n_166) );
BUFx8_ASAP7_75t_SL g167 ( .A(n_124), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_128), .B(n_3), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_110), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_121), .B(n_4), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_128), .B(n_5), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_120), .B(n_5), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_151), .A2(n_106), .B1(n_111), .B2(n_115), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_170), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_151), .A2(n_116), .B1(n_117), .B2(n_118), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_151), .A2(n_126), .B1(n_145), .B2(n_138), .Y(n_176) );
INVxp33_ASAP7_75t_L g177 ( .A(n_167), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_165), .B(n_169), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_170), .A2(n_123), .B1(n_122), .B2(n_130), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_170), .A2(n_123), .B1(n_122), .B2(n_130), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_170), .A2(n_130), .B1(n_133), .B2(n_120), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_157), .A2(n_130), .B1(n_134), .B2(n_133), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_166), .B(n_121), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_165), .B(n_127), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_166), .B(n_121), .Y(n_187) );
INVx8_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_157), .A2(n_130), .B1(n_134), .B2(n_149), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g190 ( .A1(n_157), .A2(n_149), .B1(n_140), .B2(n_127), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_166), .B(n_143), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_168), .B(n_143), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_168), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_170), .A2(n_130), .B1(n_129), .B2(n_131), .Y(n_194) );
OAI22xp33_ASAP7_75t_SL g195 ( .A1(n_150), .A2(n_129), .B1(n_131), .B2(n_140), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_170), .A2(n_130), .B1(n_141), .B2(n_148), .Y(n_196) );
OA22x2_ASAP7_75t_L g197 ( .A1(n_168), .A2(n_141), .B1(n_125), .B2(n_112), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_150), .A2(n_125), .B1(n_107), .B2(n_144), .Y(n_199) );
NAND2xp33_ASAP7_75t_SL g200 ( .A(n_168), .B(n_108), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_156), .A2(n_136), .B1(n_132), .B2(n_135), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_165), .B(n_143), .Y(n_202) );
AO22x2_ASAP7_75t_L g203 ( .A1(n_169), .A2(n_125), .B1(n_147), .B2(n_8), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_169), .B(n_147), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_156), .A2(n_142), .B1(n_137), .B2(n_114), .Y(n_207) );
OR2x6_ASAP7_75t_L g208 ( .A(n_152), .B(n_147), .Y(n_208) );
AO22x2_ASAP7_75t_L g209 ( .A1(n_171), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_162), .B(n_164), .Y(n_210) );
OA22x2_ASAP7_75t_L g211 ( .A1(n_171), .A2(n_6), .B1(n_10), .B2(n_11), .Y(n_211) );
OA22x2_ASAP7_75t_L g212 ( .A1(n_162), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_161), .A2(n_146), .B1(n_14), .B2(n_15), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g214 ( .A1(n_161), .A2(n_172), .B1(n_167), .B2(n_164), .Y(n_214) );
OAI22xp33_ASAP7_75t_SL g215 ( .A1(n_172), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_162), .A2(n_13), .B1(n_16), .B2(n_17), .Y(n_216) );
OR2x6_ASAP7_75t_L g217 ( .A(n_164), .B(n_18), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_160), .B(n_18), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
INVxp67_ASAP7_75t_SL g220 ( .A(n_178), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_176), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_174), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_199), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_206), .B(n_19), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_174), .Y(n_225) );
INVxp33_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_183), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_198), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_205), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_203), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_203), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_181), .B(n_19), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_185), .B(n_160), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_188), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_210), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_187), .B(n_160), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_188), .A2(n_155), .B(n_160), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
BUFx6f_ASAP7_75t_SL g242 ( .A(n_217), .Y(n_242) );
XOR2xp5_ASAP7_75t_L g243 ( .A(n_214), .B(n_20), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_191), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_192), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_193), .B(n_160), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_201), .B(n_160), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_186), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_207), .B(n_160), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_200), .B(n_160), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
INVxp67_ASAP7_75t_SL g253 ( .A(n_173), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_212), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_173), .B(n_160), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_208), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_175), .B(n_160), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_217), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
INVxp33_ASAP7_75t_L g263 ( .A(n_190), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_211), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_208), .B(n_160), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_217), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_175), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_209), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_195), .B(n_153), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_20), .Y(n_270) );
XOR2xp5_ASAP7_75t_L g271 ( .A(n_197), .B(n_21), .Y(n_271) );
INVxp33_ASAP7_75t_SL g272 ( .A(n_197), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_184), .B(n_21), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_179), .B(n_155), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
NOR2xp33_ASAP7_75t_SL g276 ( .A(n_215), .B(n_155), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_180), .B(n_184), .Y(n_277) );
CKINVDCx16_ASAP7_75t_R g278 ( .A(n_216), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_209), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_219), .B(n_189), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
NOR2xp67_ASAP7_75t_SL g283 ( .A(n_238), .B(n_153), .Y(n_283) );
NOR2xp33_ASAP7_75t_R g284 ( .A(n_266), .B(n_22), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_230), .B(n_189), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_224), .B(n_213), .Y(n_286) );
AND3x1_ASAP7_75t_SL g287 ( .A(n_262), .B(n_22), .C(n_23), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_219), .B(n_24), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_227), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_220), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_224), .B(n_24), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_224), .B(n_25), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_260), .B(n_25), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_228), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_248), .B(n_155), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_248), .B(n_26), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_244), .B(n_26), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_235), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_257), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_260), .B(n_27), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_257), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_222), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_228), .Y(n_307) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_230), .B(n_163), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_229), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_279), .B(n_28), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_229), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_225), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_238), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_279), .B(n_29), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_279), .B(n_29), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_252), .B(n_30), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_270), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_225), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_234), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_237), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_252), .B(n_30), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_236), .B(n_31), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_231), .B(n_163), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_242), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_244), .B(n_32), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_279), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_270), .B(n_32), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_232), .B(n_33), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_246), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_236), .B(n_33), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_253), .B(n_34), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_326), .B(n_231), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_291), .B(n_278), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_291), .B(n_262), .Y(n_336) );
INVx5_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_294), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_324), .B(n_232), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_289), .B(n_264), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_289), .B(n_264), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_290), .Y(n_342) );
BUFx4f_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_294), .B(n_268), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_317), .B(n_278), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_289), .B(n_240), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_324), .B(n_245), .Y(n_347) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_294), .B(n_233), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_317), .B(n_267), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_289), .B(n_254), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_317), .B(n_221), .Y(n_351) );
AND2x6_ASAP7_75t_L g352 ( .A(n_294), .B(n_233), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_290), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_282), .B(n_280), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_282), .B(n_240), .Y(n_355) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_282), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_290), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_290), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_296), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_324), .B(n_245), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_281), .B(n_254), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_281), .B(n_255), .Y(n_363) );
BUFx10_ASAP7_75t_L g364 ( .A(n_352), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_343), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_334), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_353), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_337), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_353), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
INVx5_ASAP7_75t_L g374 ( .A(n_338), .Y(n_374) );
BUFx8_ASAP7_75t_L g375 ( .A(n_360), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_337), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
BUFx2_ASAP7_75t_SL g378 ( .A(n_338), .Y(n_378) );
BUFx4f_ASAP7_75t_L g379 ( .A(n_352), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_334), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
BUFx4_ASAP7_75t_SL g383 ( .A(n_357), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_342), .B(n_292), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_337), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_338), .Y(n_386) );
BUFx2_ASAP7_75t_SL g387 ( .A(n_338), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_335), .Y(n_388) );
BUFx12f_ASAP7_75t_L g389 ( .A(n_360), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
BUFx12f_ASAP7_75t_L g391 ( .A(n_352), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_378), .A2(n_242), .B1(n_284), .B2(n_348), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_383), .Y(n_395) );
INVx4_ASAP7_75t_L g396 ( .A(n_379), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_388), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_379), .A2(n_335), .B1(n_345), .B2(n_324), .Y(n_398) );
CKINVDCx6p67_ASAP7_75t_R g399 ( .A(n_374), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_388), .A2(n_349), .B1(n_294), .B2(n_271), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_383), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_383), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_378), .A2(n_242), .B1(n_284), .B2(n_348), .Y(n_403) );
CKINVDCx6p67_ASAP7_75t_R g404 ( .A(n_374), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_374), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_365), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_379), .A2(n_335), .B1(n_345), .B2(n_324), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_374), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g409 ( .A1(n_386), .A2(n_243), .B(n_271), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_367), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_379), .A2(n_345), .B1(n_324), .B2(n_344), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_365), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_367), .B(n_331), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_370), .A2(n_351), .B1(n_243), .B2(n_272), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
CKINVDCx12_ASAP7_75t_R g417 ( .A(n_384), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_369), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_370), .A2(n_327), .B1(n_286), .B2(n_361), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_366), .Y(n_424) );
BUFx12f_ASAP7_75t_L g425 ( .A(n_364), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_378), .A2(n_284), .B1(n_348), .B2(n_352), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_386), .A2(n_304), .B(n_297), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_378), .A2(n_352), .B1(n_324), .B2(n_294), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_385), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_369), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_373), .Y(n_433) );
INVx8_ASAP7_75t_L g434 ( .A(n_374), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_385), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_385), .B(n_342), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_433), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_427), .A2(n_379), .B1(n_391), .B2(n_344), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_394), .B(n_368), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_426), .A2(n_386), .B(n_292), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_398), .A2(n_375), .B1(n_370), .B2(n_371), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_397), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_409), .A2(n_331), .B1(n_268), .B2(n_263), .C1(n_297), .C2(n_304), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_435), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_433), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_407), .A2(n_375), .B1(n_377), .B2(n_370), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_400), .A2(n_276), .B(n_331), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_400), .A2(n_375), .B1(n_371), .B2(n_370), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_410), .B(n_372), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_394), .B(n_368), .Y(n_452) );
NOR2xp67_ASAP7_75t_SL g453 ( .A(n_401), .B(n_391), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_434), .A2(n_375), .B1(n_371), .B2(n_370), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_434), .A2(n_391), .B1(n_389), .B2(n_387), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_427), .A2(n_286), .B(n_322), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_434), .A2(n_391), .B1(n_389), .B2(n_387), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_434), .A2(n_375), .B1(n_377), .B2(n_371), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_434), .A2(n_375), .B1(n_377), .B2(n_371), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_399), .A2(n_375), .B1(n_377), .B2(n_371), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_399), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_393), .A2(n_379), .B1(n_391), .B2(n_374), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_404), .A2(n_375), .B1(n_377), .B2(n_389), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_436), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_415), .A2(n_331), .B1(n_297), .B2(n_304), .C1(n_325), .C2(n_301), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_401), .A2(n_389), .B1(n_387), .B2(n_377), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_394), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
CKINVDCx11_ASAP7_75t_R g471 ( .A(n_406), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_405), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_416), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_402), .A2(n_374), .B1(n_379), .B2(n_389), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_402), .A2(n_387), .B1(n_374), .B2(n_379), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_423), .A2(n_344), .B1(n_368), .B2(n_386), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_404), .A2(n_403), .B1(n_327), .B2(n_286), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_408), .A2(n_374), .B1(n_385), .B2(n_381), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_408), .A2(n_374), .B1(n_385), .B2(n_381), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_428), .A2(n_344), .B1(n_390), .B2(n_372), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_418), .Y(n_482) );
INVx6_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
BUFx12f_ASAP7_75t_L g484 ( .A(n_395), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_412), .A2(n_327), .B1(n_286), .B2(n_374), .Y(n_485) );
BUFx4f_ASAP7_75t_SL g486 ( .A(n_413), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_396), .A2(n_327), .B1(n_286), .B2(n_374), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_418), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_425), .A2(n_374), .B1(n_385), .B2(n_381), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g491 ( .A1(n_414), .A2(n_304), .B1(n_297), .B2(n_325), .C1(n_301), .C2(n_292), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_429), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_416), .B(n_380), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_429), .B(n_372), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_396), .A2(n_327), .B1(n_286), .B2(n_339), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_420), .A2(n_390), .B1(n_382), .B2(n_392), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_420), .Y(n_497) );
AOI211xp5_ASAP7_75t_L g498 ( .A1(n_422), .A2(n_327), .B(n_292), .C(n_273), .Y(n_498) );
BUFx12f_ASAP7_75t_L g499 ( .A(n_425), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_425), .A2(n_324), .B1(n_369), .B2(n_376), .Y(n_500) );
BUFx12f_ASAP7_75t_L g501 ( .A(n_396), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_417), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_420), .B(n_382), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_421), .B(n_380), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_421), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_417), .A2(n_327), .B1(n_286), .B2(n_287), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_421), .A2(n_392), .B1(n_390), .B2(n_382), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_433), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_396), .A2(n_327), .B1(n_286), .B2(n_339), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_439), .A2(n_430), .B1(n_381), .B2(n_364), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_439), .A2(n_339), .B1(n_352), .B2(n_361), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_498), .B(n_390), .C(n_382), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_449), .A2(n_339), .B1(n_352), .B2(n_361), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_440), .B(n_424), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_449), .A2(n_339), .B1(n_352), .B2(n_361), .Y(n_515) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_450), .A2(n_330), .B1(n_322), .B2(n_325), .C(n_301), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_498), .A2(n_430), .B1(n_392), .B2(n_376), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_440), .B(n_424), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_452), .B(n_424), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_441), .A2(n_456), .B1(n_458), .B2(n_478), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_444), .A2(n_287), .B1(n_328), .B2(n_346), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_465), .A2(n_392), .B1(n_432), .B2(n_381), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_457), .A2(n_352), .B1(n_347), .B2(n_361), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_452), .B(n_431), .Y(n_524) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_457), .A2(n_431), .B(n_380), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_444), .A2(n_347), .B1(n_328), .B2(n_384), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_462), .A2(n_381), .B1(n_364), .B2(n_373), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_447), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_476), .A2(n_347), .B1(n_328), .B2(n_384), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_476), .A2(n_287), .B1(n_328), .B2(n_346), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_481), .A2(n_347), .B1(n_328), .B2(n_384), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_490), .B(n_373), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_447), .B(n_454), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_506), .A2(n_381), .B1(n_328), .B2(n_419), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_481), .A2(n_347), .B1(n_328), .B2(n_384), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_485), .A2(n_328), .B1(n_329), .B2(n_346), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_454), .B(n_464), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_471), .B(n_322), .C(n_330), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_506), .A2(n_330), .B1(n_255), .B2(n_273), .C(n_321), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_468), .A2(n_419), .B1(n_223), .B2(n_332), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_467), .A2(n_332), .B1(n_364), .B2(n_316), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_487), .A2(n_329), .B1(n_295), .B2(n_364), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_467), .A2(n_329), .B1(n_295), .B2(n_364), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_469), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_495), .A2(n_295), .B1(n_364), .B2(n_315), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_479), .B(n_321), .C(n_316), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_462), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_482), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_509), .A2(n_295), .B1(n_364), .B2(n_310), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_442), .A2(n_295), .B1(n_310), .B2(n_314), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_448), .A2(n_295), .B1(n_310), .B2(n_314), .Y(n_553) );
AOI222xp33_ASAP7_75t_L g554 ( .A1(n_486), .A2(n_316), .B1(n_300), .B2(n_321), .C1(n_269), .C2(n_362), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_488), .Y(n_555) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_445), .A2(n_433), .B1(n_419), .B2(n_373), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_501), .A2(n_373), .B1(n_433), .B2(n_419), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_492), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_480), .B(n_300), .C(n_154), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_501), .A2(n_295), .B1(n_314), .B2(n_310), .Y(n_560) );
AOI21xp33_ASAP7_75t_L g561 ( .A1(n_474), .A2(n_300), .B(n_363), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_491), .A2(n_356), .B1(n_363), .B2(n_362), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_463), .A2(n_295), .B1(n_314), .B2(n_315), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_499), .A2(n_373), .B1(n_315), .B2(n_337), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_492), .B(n_342), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_455), .A2(n_295), .B1(n_315), .B2(n_303), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_438), .B(n_472), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_459), .A2(n_295), .B1(n_303), .B2(n_354), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_443), .B(n_226), .Y(n_569) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_461), .B(n_373), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_460), .A2(n_303), .B1(n_354), .B2(n_305), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_493), .B(n_373), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_491), .A2(n_305), .B1(n_373), .B2(n_355), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_475), .A2(n_373), .B1(n_358), .B2(n_356), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_470), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_502), .A2(n_305), .B1(n_355), .B2(n_341), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_483), .A2(n_355), .B1(n_341), .B2(n_340), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_493), .B(n_504), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_500), .B(n_256), .C(n_259), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_483), .A2(n_340), .B1(n_350), .B2(n_358), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_496), .B(n_358), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_483), .A2(n_285), .B1(n_319), .B2(n_320), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_453), .A2(n_241), .B1(n_336), .B2(n_319), .C(n_320), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_466), .A2(n_285), .B1(n_309), .B2(n_311), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_470), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_473), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_496), .A2(n_311), .B1(n_307), .B2(n_309), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_507), .A2(n_337), .B1(n_311), .B2(n_309), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_508), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_507), .A2(n_337), .B1(n_308), .B2(n_307), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_451), .B(n_296), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_477), .A2(n_298), .B1(n_309), .B2(n_311), .Y(n_592) );
NAND2xp33_ASAP7_75t_SL g593 ( .A(n_489), .B(n_333), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_484), .A2(n_308), .B1(n_307), .B2(n_298), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_484), .A2(n_298), .B1(n_309), .B2(n_311), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_494), .A2(n_296), .B1(n_298), .B2(n_307), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_503), .A2(n_308), .B1(n_307), .B2(n_296), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_473), .A2(n_296), .B1(n_298), .B2(n_308), .Y(n_598) );
OAI221xp5_ASAP7_75t_SL g599 ( .A1(n_504), .A2(n_299), .B1(n_277), .B2(n_250), .C(n_251), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_497), .A2(n_308), .B1(n_333), .B2(n_326), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_497), .B(n_153), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_505), .B(n_34), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_437), .A2(n_308), .B1(n_326), .B2(n_302), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_578), .B(n_505), .Y(n_604) );
OAI221xp5_ASAP7_75t_SL g605 ( .A1(n_539), .A2(n_446), .B1(n_437), .B2(n_299), .C(n_249), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_529), .B(n_508), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_550), .B(n_508), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_550), .B(n_508), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_520), .B(n_247), .C(n_299), .D(n_239), .Y(n_609) );
OA211x2_ASAP7_75t_L g610 ( .A1(n_533), .A2(n_35), .B(n_36), .C(n_37), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_512), .A2(n_326), .B1(n_313), .B2(n_302), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_555), .B(n_35), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g613 ( .A1(n_521), .A2(n_251), .B1(n_326), .B2(n_265), .C(n_306), .Y(n_613) );
NAND4xp25_ASAP7_75t_SL g614 ( .A(n_511), .B(n_37), .C(n_38), .D(n_39), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_512), .A2(n_313), .B1(n_288), .B2(n_302), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_525), .B(n_153), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_521), .A2(n_288), .B1(n_302), .B2(n_306), .C(n_293), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_554), .B(n_153), .C(n_154), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_548), .B(n_559), .C(n_531), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_531), .B(n_153), .C(n_154), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_555), .B(n_38), .Y(n_621) );
AOI21xp5_ASAP7_75t_SL g622 ( .A1(n_517), .A2(n_323), .B(n_313), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_541), .A2(n_302), .B1(n_288), .B2(n_306), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_527), .A2(n_288), .B1(n_302), .B2(n_306), .C(n_293), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_556), .B(n_153), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_558), .B(n_40), .Y(n_626) );
OA21x2_ASAP7_75t_L g627 ( .A1(n_581), .A2(n_323), .B(n_274), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_532), .A2(n_313), .B1(n_288), .B2(n_302), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_558), .B(n_40), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_534), .B(n_41), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_525), .B(n_163), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_525), .B(n_163), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_564), .B(n_153), .C(n_154), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_538), .B(n_41), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_510), .B(n_602), .C(n_567), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_514), .B(n_42), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_525), .B(n_163), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_545), .B(n_163), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_536), .A2(n_153), .B(n_154), .C(n_158), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_545), .B(n_163), .Y(n_640) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_528), .A2(n_42), .B(n_43), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_542), .B(n_153), .C(n_154), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_546), .B(n_163), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_518), .B(n_154), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_542), .A2(n_288), .B1(n_293), .B2(n_313), .C(n_312), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_519), .B(n_154), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_546), .B(n_163), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_530), .A2(n_288), .B1(n_312), .B2(n_293), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_575), .B(n_163), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_556), .B(n_154), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_524), .B(n_154), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_523), .A2(n_312), .B1(n_323), .B2(n_318), .Y(n_652) );
NAND2xp33_ASAP7_75t_L g653 ( .A(n_593), .B(n_312), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_562), .B(n_261), .C(n_258), .D(n_318), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_594), .B(n_158), .C(n_275), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_573), .A2(n_318), .B1(n_275), .B2(n_158), .Y(n_656) );
AOI222xp33_ASAP7_75t_L g657 ( .A1(n_540), .A2(n_158), .B1(n_318), .B2(n_283), .C1(n_48), .C2(n_49), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_557), .B(n_158), .C(n_318), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_544), .A2(n_158), .B1(n_318), .B2(n_283), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_561), .A2(n_158), .B1(n_318), .B2(n_283), .C(n_50), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_585), .B(n_158), .Y(n_661) );
OAI221xp5_ASAP7_75t_SL g662 ( .A1(n_562), .A2(n_44), .B1(n_45), .B2(n_47), .C(n_51), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_526), .B(n_283), .C(n_55), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_579), .A2(n_53), .B1(n_56), .B2(n_60), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_587), .B(n_61), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_535), .A2(n_64), .B1(n_65), .B2(n_69), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_549), .B(n_70), .C(n_73), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_587), .B(n_74), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_585), .B(n_76), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_586), .B(n_81), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_586), .B(n_82), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_570), .B(n_85), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_513), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_522), .B(n_90), .C(n_91), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_570), .A2(n_94), .B(n_95), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_565), .B(n_96), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g677 ( .A1(n_595), .A2(n_98), .B(n_101), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_591), .B(n_105), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_589), .B(n_601), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_589), .B(n_601), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_580), .B(n_577), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_599), .B(n_515), .C(n_590), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_584), .B(n_563), .Y(n_683) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_583), .A2(n_597), .B(n_574), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_576), .B(n_592), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_588), .B(n_582), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_593), .B(n_600), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_571), .B(n_568), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g689 ( .A(n_569), .B(n_537), .C(n_553), .D(n_552), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_596), .B(n_560), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g691 ( .A1(n_566), .A2(n_547), .B(n_551), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_543), .B(n_516), .Y(n_692) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_603), .A2(n_598), .B(n_520), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_578), .B(n_572), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_520), .B(n_539), .C(n_512), .D(n_521), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_695), .B(n_693), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_604), .B(n_694), .Y(n_697) );
AO21x2_ASAP7_75t_L g698 ( .A1(n_616), .A2(n_637), .B(n_631), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_682), .A2(n_683), .B1(n_618), .B2(n_686), .Y(n_699) );
AO21x2_ASAP7_75t_L g700 ( .A1(n_632), .A2(n_637), .B(n_650), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_635), .B(n_650), .C(n_625), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_689), .B(n_681), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_606), .B(n_607), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_679), .Y(n_704) );
NAND4xp75_ASAP7_75t_L g705 ( .A(n_610), .B(n_625), .C(n_687), .D(n_672), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_683), .A2(n_686), .B1(n_688), .B2(n_619), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_641), .B(n_614), .C(n_662), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_644), .Y(n_708) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_658), .B(n_622), .Y(n_709) );
INVx3_ASAP7_75t_L g710 ( .A(n_680), .Y(n_710) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_653), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_680), .B(n_608), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_684), .B(n_687), .C(n_634), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_646), .B(n_651), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_609), .A2(n_692), .B1(n_690), .B2(n_685), .Y(n_715) );
NAND4xp75_ASAP7_75t_L g716 ( .A(n_672), .B(n_623), .C(n_636), .D(n_630), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_638), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_638), .B(n_643), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_640), .B(n_661), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_640), .B(n_649), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_605), .B(n_675), .C(n_677), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_612), .Y(n_722) );
NOR3xp33_ASAP7_75t_L g723 ( .A(n_621), .B(n_626), .C(n_629), .Y(n_723) );
OAI211xp5_ASAP7_75t_L g724 ( .A1(n_691), .A2(n_657), .B(n_613), .C(n_617), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_643), .B(n_647), .Y(n_725) );
AND2x2_ASAP7_75t_SL g726 ( .A(n_653), .B(n_669), .Y(n_726) );
OAI211xp5_ASAP7_75t_L g727 ( .A1(n_639), .A2(n_645), .B(n_654), .C(n_633), .Y(n_727) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_642), .B(n_655), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_615), .A2(n_611), .B1(n_620), .B2(n_674), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_660), .B(n_667), .C(n_664), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_666), .B(n_665), .C(n_668), .Y(n_731) );
NAND4xp75_ASAP7_75t_L g732 ( .A(n_670), .B(n_671), .C(n_678), .D(n_676), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_627), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g734 ( .A(n_673), .B(n_656), .C(n_663), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_627), .B(n_648), .Y(n_735) );
XNOR2x1_ASAP7_75t_L g736 ( .A(n_628), .B(n_652), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_624), .B(n_659), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_695), .B(n_693), .C(n_635), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_695), .B(n_618), .C(n_641), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_695), .B(n_693), .C(n_635), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_695), .B(n_693), .C(n_635), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_695), .A2(n_682), .B1(n_520), .B2(n_683), .Y(n_742) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_625), .Y(n_743) );
NAND4xp75_ASAP7_75t_L g744 ( .A(n_610), .B(n_650), .C(n_625), .D(n_402), .Y(n_744) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_695), .B(n_693), .C(n_635), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_695), .B(n_471), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_694), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_695), .A2(n_682), .B1(n_520), .B2(n_683), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_694), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_695), .A2(n_682), .B1(n_520), .B2(n_683), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_604), .B(n_694), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_695), .B(n_693), .C(n_635), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_695), .A2(n_682), .B1(n_520), .B2(n_683), .Y(n_753) );
INVx1_ASAP7_75t_SL g754 ( .A(n_749), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_717), .Y(n_755) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_701), .B(n_705), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_697), .B(n_751), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_709), .B(n_726), .Y(n_758) );
NOR4xp25_ASAP7_75t_L g759 ( .A(n_738), .B(n_745), .C(n_741), .D(n_752), .Y(n_759) );
XNOR2x2_ASAP7_75t_L g760 ( .A(n_740), .B(n_713), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_696), .A2(n_702), .B1(n_753), .B2(n_748), .Y(n_761) );
XOR2x2_ASAP7_75t_L g762 ( .A(n_746), .B(n_742), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_750), .A2(n_724), .B1(n_739), .B2(n_699), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_706), .B(n_722), .Y(n_764) );
NAND4xp75_ASAP7_75t_L g765 ( .A(n_728), .B(n_726), .C(n_737), .D(n_735), .Y(n_765) );
INVx2_ASAP7_75t_SL g766 ( .A(n_710), .Y(n_766) );
NOR4xp25_ASAP7_75t_L g767 ( .A(n_715), .B(n_727), .C(n_743), .D(n_731), .Y(n_767) );
INVx4_ASAP7_75t_L g768 ( .A(n_700), .Y(n_768) );
AND4x2_ASAP7_75t_L g769 ( .A(n_705), .B(n_721), .C(n_716), .D(n_711), .Y(n_769) );
NOR4xp25_ASAP7_75t_L g770 ( .A(n_708), .B(n_730), .C(n_714), .D(n_747), .Y(n_770) );
INVx3_ASAP7_75t_L g771 ( .A(n_700), .Y(n_771) );
XOR2x2_ASAP7_75t_L g772 ( .A(n_707), .B(n_744), .Y(n_772) );
NAND4xp75_ASAP7_75t_SL g773 ( .A(n_736), .B(n_700), .C(n_719), .D(n_718), .Y(n_773) );
NOR3xp33_ASAP7_75t_L g774 ( .A(n_734), .B(n_723), .C(n_729), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_703), .B(n_704), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g776 ( .A(n_736), .B(n_733), .C(n_703), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_704), .B(n_710), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_764), .B(n_712), .Y(n_778) );
XNOR2xp5_ASAP7_75t_L g779 ( .A(n_772), .B(n_732), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_761), .B(n_712), .Y(n_780) );
XNOR2xp5_ASAP7_75t_L g781 ( .A(n_772), .B(n_718), .Y(n_781) );
INVxp67_ASAP7_75t_L g782 ( .A(n_756), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g783 ( .A(n_762), .B(n_719), .Y(n_783) );
XOR2x2_ASAP7_75t_L g784 ( .A(n_762), .B(n_698), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_775), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_775), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_757), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_777), .Y(n_788) );
XNOR2xp5_ASAP7_75t_L g789 ( .A(n_763), .B(n_720), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_755), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_754), .Y(n_791) );
XNOR2x2_ASAP7_75t_L g792 ( .A(n_760), .B(n_720), .Y(n_792) );
INVxp67_ASAP7_75t_L g793 ( .A(n_776), .Y(n_793) );
XOR2x2_ASAP7_75t_L g794 ( .A(n_774), .B(n_698), .Y(n_794) );
XNOR2x2_ASAP7_75t_L g795 ( .A(n_765), .B(n_725), .Y(n_795) );
OA22x2_ASAP7_75t_L g796 ( .A1(n_782), .A2(n_758), .B1(n_768), .B2(n_759), .Y(n_796) );
OA22x2_ASAP7_75t_L g797 ( .A1(n_779), .A2(n_758), .B1(n_768), .B2(n_769), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_787), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_791), .Y(n_799) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_779), .B(n_765), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_791), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_788), .Y(n_802) );
XNOR2x1_ASAP7_75t_L g803 ( .A(n_792), .B(n_773), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_781), .Y(n_804) );
AOI22x1_ASAP7_75t_L g805 ( .A1(n_792), .A2(n_768), .B1(n_769), .B2(n_767), .Y(n_805) );
OAI22x1_ASAP7_75t_L g806 ( .A1(n_793), .A2(n_766), .B1(n_770), .B2(n_771), .Y(n_806) );
INVx1_ASAP7_75t_SL g807 ( .A(n_790), .Y(n_807) );
AO22x2_ASAP7_75t_L g808 ( .A1(n_785), .A2(n_786), .B1(n_794), .B2(n_784), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_807), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_799), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_799), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_801), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_801), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_802), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_802), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_798), .Y(n_816) );
OA22x2_ASAP7_75t_L g817 ( .A1(n_809), .A2(n_804), .B1(n_806), .B2(n_781), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_809), .Y(n_818) );
AOI22x1_ASAP7_75t_L g819 ( .A1(n_815), .A2(n_808), .B1(n_804), .B2(n_806), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_814), .A2(n_800), .B1(n_808), .B2(n_784), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_814), .Y(n_821) );
AOI22x1_ASAP7_75t_SL g822 ( .A1(n_818), .A2(n_800), .B1(n_805), .B2(n_795), .Y(n_822) );
INVx4_ASAP7_75t_SL g823 ( .A(n_821), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_820), .A2(n_803), .B1(n_808), .B2(n_797), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_823), .Y(n_825) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_824), .B(n_803), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_825), .B(n_817), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_826), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_827), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_828), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_830), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_829), .Y(n_832) );
AO22x2_ASAP7_75t_L g833 ( .A1(n_832), .A2(n_822), .B1(n_816), .B2(n_810), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_833), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_834), .A2(n_832), .B1(n_819), .B2(n_831), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_835), .Y(n_836) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_836), .A2(n_819), .B1(n_797), .B2(n_796), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_837), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g839 ( .A1(n_838), .A2(n_811), .B1(n_812), .B2(n_813), .C(n_780), .Y(n_839) );
AOI211xp5_ASAP7_75t_L g840 ( .A1(n_839), .A2(n_789), .B(n_783), .C(n_778), .Y(n_840) );
endmodule