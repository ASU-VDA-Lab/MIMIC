module fake_jpeg_21003_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_19),
.B1(n_37),
.B2(n_22),
.Y(n_63)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_39),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_25),
.B1(n_31),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_19),
.B1(n_43),
.B2(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_67),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_25),
.B1(n_31),
.B2(n_47),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_96),
.B1(n_97),
.B2(n_101),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_31),
.B1(n_25),
.B2(n_27),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_49),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_84),
.C(n_93),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_95),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_92),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_35),
.B1(n_21),
.B2(n_28),
.Y(n_131)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_91),
.Y(n_130)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_49),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_41),
.B1(n_36),
.B2(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_24),
.B1(n_19),
.B2(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_56),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_37),
.B1(n_39),
.B2(n_21),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_44),
.B1(n_61),
.B2(n_54),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_103),
.B1(n_108),
.B2(n_89),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_61),
.B1(n_54),
.B2(n_35),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_84),
.B1(n_83),
.B2(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_123),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_126),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_129),
.Y(n_156)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_42),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_105),
.B1(n_129),
.B2(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_73),
.B1(n_76),
.B2(n_82),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_149),
.B1(n_155),
.B2(n_130),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_153),
.B(n_26),
.Y(n_177)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_42),
.C(n_46),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_50),
.C(n_48),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_71),
.B1(n_86),
.B2(n_90),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_114),
.B1(n_124),
.B2(n_111),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_119),
.B1(n_105),
.B2(n_102),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_154),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_103),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_92),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_86),
.B1(n_71),
.B2(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_94),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_160),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_26),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_69),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_29),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_120),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_183),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_167),
.A2(n_168),
.B1(n_179),
.B2(n_184),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_124),
.B1(n_111),
.B2(n_106),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_148),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_172),
.B(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_29),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_182),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_149),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_106),
.B1(n_104),
.B2(n_115),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_181),
.B1(n_118),
.B2(n_109),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_104),
.B1(n_115),
.B2(n_130),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_146),
.C(n_134),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_156),
.C(n_150),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_130),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_120),
.B1(n_28),
.B2(n_118),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_156),
.B1(n_154),
.B2(n_146),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_139),
.B1(n_136),
.B2(n_109),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_188),
.B(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_0),
.B(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_194),
.B(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_206),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_202),
.C(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_140),
.C(n_144),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_160),
.A3(n_135),
.B1(n_138),
.B2(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_169),
.C(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_209),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_168),
.B1(n_167),
.B2(n_184),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_38),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_118),
.B1(n_50),
.B2(n_48),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_224),
.B1(n_181),
.B2(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_38),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_34),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_221),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_162),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_163),
.B(n_182),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_225),
.A2(n_227),
.B(n_249),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_193),
.A2(n_163),
.B(n_179),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_230),
.A2(n_23),
.B1(n_18),
.B2(n_30),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_188),
.B(n_186),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_246),
.B(n_247),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_165),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_165),
.C(n_38),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_202),
.C(n_198),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_50),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_248),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_32),
.B(n_13),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_197),
.A2(n_206),
.B(n_209),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_48),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_2),
.B(n_3),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_210),
.A2(n_18),
.B1(n_23),
.B2(n_30),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_195),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_268),
.C(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_262),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_210),
.B1(n_207),
.B2(n_217),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_238),
.B1(n_230),
.B2(n_242),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_215),
.B(n_204),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_227),
.A2(n_204),
.B(n_14),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_226),
.B1(n_242),
.B2(n_233),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_243),
.C(n_245),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_32),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_271),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_255),
.B1(n_269),
.B2(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_244),
.C(n_231),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_284),
.C(n_287),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_226),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_258),
.B(n_247),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_289),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_244),
.C(n_228),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_286),
.A2(n_263),
.B1(n_258),
.B2(n_264),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_233),
.C(n_239),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_246),
.B(n_249),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_265),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_256),
.B1(n_267),
.B2(n_260),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_303),
.B1(n_58),
.B2(n_23),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_252),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_298),
.B1(n_299),
.B2(n_288),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_271),
.C(n_262),
.Y(n_297)
);

OAI321xp33_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_11),
.A3(n_16),
.B1(n_15),
.B2(n_14),
.C(n_7),
.Y(n_312)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_13),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_284),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_58),
.C(n_46),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_58),
.C(n_46),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_283),
.B1(n_288),
.B2(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_308),
.Y(n_318)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_272),
.B1(n_273),
.B2(n_276),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_304),
.B(n_296),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_312),
.B(n_291),
.Y(n_323)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_34),
.C(n_30),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_32),
.B1(n_18),
.B2(n_9),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_30),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_306),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_322),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_9),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_300),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_307),
.CI(n_314),
.CON(n_326),
.SN(n_326)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_309),
.A2(n_292),
.B1(n_302),
.B2(n_5),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_315),
.C(n_4),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_331),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_332),
.C(n_319),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_8),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_336),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_317),
.C(n_325),
.Y(n_336)
);

AOI221xp5_ASAP7_75t_SL g337 ( 
.A1(n_335),
.A2(n_329),
.B1(n_10),
.B2(n_7),
.C(n_12),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_337),
.A2(n_333),
.B(n_12),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_338),
.B(n_12),
.C(n_16),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_6),
.B(n_3),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_3),
.B(n_5),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_3),
.C(n_5),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_5),
.Y(n_345)
);


endmodule