module fake_ariane_109_n_482 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_482);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_482;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_180;
wire n_124;
wire n_119;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_34;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_133;
wire n_66;
wire n_205;
wire n_341;
wire n_71;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_319;
wire n_49;
wire n_416;
wire n_283;
wire n_50;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_36;
wire n_370;
wire n_189;
wire n_72;
wire n_286;
wire n_443;
wire n_57;
wire n_424;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_32;
wire n_410;
wire n_379;
wire n_445;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_52;
wire n_441;
wire n_385;
wire n_73;
wire n_327;
wire n_77;
wire n_372;
wire n_377;
wire n_396;
wire n_23;
wire n_399;
wire n_87;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_41;
wire n_140;
wire n_419;
wire n_151;
wire n_28;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_59;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_35;
wire n_272;
wire n_54;
wire n_339;
wire n_167;
wire n_90;
wire n_38;
wire n_422;
wire n_47;
wire n_153;
wire n_269;
wire n_75;
wire n_158;
wire n_69;
wire n_259;
wire n_95;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_320;
wire n_309;
wire n_115;
wire n_331;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_62;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_79;
wire n_271;
wire n_465;
wire n_247;
wire n_91;
wire n_369;
wire n_240;
wire n_128;
wire n_224;
wire n_44;
wire n_82;
wire n_31;
wire n_420;
wire n_439;
wire n_222;
wire n_478;
wire n_256;
wire n_326;
wire n_227;
wire n_48;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_427;
wire n_108;
wire n_303;
wire n_442;
wire n_168;
wire n_81;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_88;
wire n_141;
wire n_390;
wire n_104;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_56;
wire n_60;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_86;
wire n_361;
wire n_458;
wire n_89;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_74;
wire n_40;
wire n_181;
wire n_53;
wire n_362;
wire n_260;
wire n_310;
wire n_236;
wire n_281;
wire n_24;
wire n_461;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_464;
wire n_297;
wire n_290;
wire n_46;
wire n_84;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_452;
wire n_178;
wire n_42;
wire n_308;
wire n_417;
wire n_201;
wire n_70;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_94;
wire n_284;
wire n_448;
wire n_249;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_468;
wire n_61;
wire n_102;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_43;
wire n_407;
wire n_27;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_55;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_68;
wire n_415;
wire n_78;
wire n_63;
wire n_99;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_25;
wire n_83;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_67;
wire n_306;
wire n_313;
wire n_92;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_33;
wire n_324;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_51;
wire n_76;
wire n_342;
wire n_26;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_30;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_45;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_121;
wire n_118;
wire n_411;
wire n_353;
wire n_241;
wire n_29;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_80;
wire n_480;
wire n_211;
wire n_97;
wire n_408;
wire n_322;
wire n_251;
wire n_116;
wire n_397;
wire n_471;
wire n_351;
wire n_39;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_127;

BUFx5_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_13),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_18),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_0),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_24),
.A2(n_1),
.B(n_3),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

OR2x6_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_36),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_28),
.B1(n_38),
.B2(n_34),
.Y(n_70)
);

NOR2x1p5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_46),
.Y(n_73)
);

AND3x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_29),
.C(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_55),
.B1(n_50),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_55),
.B1(n_48),
.B2(n_47),
.Y(n_80)
);

AND2x6_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_55),
.B1(n_47),
.B2(n_27),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_62),
.Y(n_88)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_47),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_47),
.B1(n_26),
.B2(n_35),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_40),
.B1(n_30),
.B2(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_66),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_31),
.B1(n_66),
.B2(n_35),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_52),
.B(n_26),
.C(n_42),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_33),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_33),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_39),
.B1(n_52),
.B2(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_73),
.B1(n_65),
.B2(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_23),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_75),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_52),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_52),
.B1(n_59),
.B2(n_72),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_69),
.B(n_58),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_69),
.B(n_58),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_69),
.B(n_58),
.C(n_59),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_72),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_72),
.B(n_59),
.C(n_56),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_72),
.B(n_59),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_72),
.B(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

O2A1O1Ixp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_53),
.B(n_56),
.C(n_54),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_57),
.B(n_54),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_57),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_4),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_57),
.Y(n_132)
);

O2A1O1Ixp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_54),
.B(n_51),
.C(n_23),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_79),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_84),
.B(n_23),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_23),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_54),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_78),
.A2(n_51),
.B(n_23),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_83),
.A2(n_51),
.B1(n_7),
.B2(n_10),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_51),
.B(n_7),
.C(n_11),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_23),
.B(n_11),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_92),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_87),
.A2(n_5),
.B(n_15),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_16),
.B1(n_17),
.B2(n_105),
.Y(n_145)
);

OR2x6_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_17),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_84),
.A2(n_87),
.B1(n_93),
.B2(n_96),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_93),
.B(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_97),
.B(n_101),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_81),
.A2(n_88),
.B(n_89),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_90),
.A2(n_88),
.B(n_98),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_79),
.A2(n_63),
.B1(n_82),
.B2(n_70),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_90),
.A2(n_88),
.B(n_98),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_110),
.B(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_109),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_153),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_154),
.B(n_128),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_123),
.Y(n_161)
);

AOI221x1_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_142),
.B1(n_139),
.B2(n_141),
.C(n_145),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_149),
.B(n_135),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_150),
.B(n_114),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_121),
.B(n_138),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_113),
.B(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_151),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_119),
.B(n_144),
.C(n_137),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_115),
.B1(n_129),
.B2(n_140),
.Y(n_169)
);

AO31x2_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_144),
.A3(n_122),
.B(n_111),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_111),
.B1(n_118),
.B2(n_125),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_136),
.B(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

AO31x2_ASAP7_75t_L g175 ( 
.A1(n_118),
.A2(n_115),
.A3(n_117),
.B(n_153),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_130),
.B(n_70),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_148),
.B(n_110),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_153),
.B1(n_134),
.B2(n_135),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_124),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_110),
.B(n_152),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_150),
.B(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_79),
.B(n_85),
.C(n_153),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

AO31x2_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_117),
.A3(n_153),
.B(n_101),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_124),
.B(n_99),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_79),
.B1(n_134),
.B2(n_63),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_134),
.B(n_124),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_159),
.B(n_183),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_183),
.B(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_168),
.B(n_155),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_188),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_160),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_185),
.B(n_189),
.Y(n_203)
);

AO21x2_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_177),
.B(n_166),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_176),
.B1(n_171),
.B2(n_169),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_163),
.B(n_161),
.C(n_171),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_181),
.Y(n_209)
);

AO31x2_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_174),
.A3(n_190),
.B(n_175),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_173),
.B(n_174),
.Y(n_211)
);

AO31x2_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_187),
.A3(n_178),
.B(n_170),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_160),
.B1(n_186),
.B2(n_157),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_164),
.B(n_159),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_191),
.B(n_158),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_170),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_159),
.B(n_164),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_159),
.B(n_158),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_159),
.B(n_183),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_182),
.B(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_158),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g229 ( 
.A1(n_164),
.A2(n_159),
.B(n_183),
.Y(n_229)
);

AO21x2_ASAP7_75t_L g230 ( 
.A1(n_159),
.A2(n_158),
.B(n_115),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_155),
.A2(n_182),
.B(n_165),
.Y(n_231)
);

AOI21x1_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_231),
.B(n_194),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_195),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_193),
.B(n_229),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

AO21x2_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_203),
.B(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_219),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_210),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_210),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_218),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_224),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_230),
.Y(n_250)
);

AO21x2_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_204),
.B(n_217),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_224),
.Y(n_256)
);

AO31x2_ASAP7_75t_L g257 ( 
.A1(n_205),
.A2(n_228),
.A3(n_207),
.B(n_206),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_208),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

NOR2x1_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_197),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_223),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_223),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_253),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_230),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_278),
.Y(n_283)
);

BUFx2_ASAP7_75t_SL g284 ( 
.A(n_270),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_246),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_246),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_246),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_258),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_256),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_246),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_209),
.B1(n_201),
.B2(n_239),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_243),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_243),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_274),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_276),
.Y(n_301)
);

OA21x2_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_235),
.B(n_232),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_243),
.Y(n_303)
);

OR2x6_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_254),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_256),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_264),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_258),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_281),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_279),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_277),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_277),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_280),
.Y(n_326)
);

OR2x6_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_259),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_243),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_257),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_262),
.B(n_233),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_233),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_306),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_300),
.B(n_238),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_273),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_233),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_333),
.A2(n_295),
.B1(n_293),
.B2(n_215),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_289),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_SL g359 ( 
.A(n_328),
.B(n_284),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_289),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_313),
.B(n_304),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_301),
.Y(n_362)
);

AOI21xp33_ASAP7_75t_SL g363 ( 
.A1(n_333),
.A2(n_200),
.B(n_283),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_339),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_308),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_336),
.B(n_292),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_315),
.B(n_293),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_329),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_348),
.A2(n_336),
.B1(n_332),
.B2(n_327),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_366),
.A2(n_295),
.B1(n_332),
.B2(n_233),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_342),
.Y(n_371)
);

AOI221xp5_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_330),
.B1(n_317),
.B2(n_262),
.C(n_320),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_318),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_320),
.A3(n_318),
.B1(n_317),
.B2(n_326),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_366),
.A2(n_215),
.B1(n_327),
.B2(n_338),
.Y(n_375)
);

OAI322xp33_ASAP7_75t_L g376 ( 
.A1(n_355),
.A2(n_323),
.A3(n_337),
.B1(n_335),
.B2(n_324),
.C1(n_285),
.C2(n_330),
.Y(n_376)
);

AOI221xp5_ASAP7_75t_L g377 ( 
.A1(n_350),
.A2(n_301),
.B1(n_294),
.B2(n_297),
.C(n_296),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_L g378 ( 
.A1(n_364),
.A2(n_327),
.B1(n_304),
.B2(n_285),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_354),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_346),
.B(n_329),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_364),
.A2(n_313),
.B1(n_338),
.B2(n_327),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_326),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_313),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_338),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_346),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_301),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_360),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_370),
.A2(n_338),
.B1(n_327),
.B2(n_346),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_362),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_369),
.A2(n_361),
.B(n_353),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_368),
.A2(n_361),
.B1(n_359),
.B2(n_238),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_L g398 ( 
.A1(n_370),
.A2(n_374),
.B(n_368),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_361),
.B1(n_297),
.B2(n_296),
.Y(n_400)
);

AOI221xp5_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_341),
.B1(n_343),
.B2(n_357),
.C(n_356),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_296),
.B1(n_297),
.B2(n_294),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_294),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_377),
.A2(n_292),
.B1(n_284),
.B2(n_352),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_378),
.A2(n_303),
.B1(n_359),
.B2(n_354),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_378),
.A2(n_380),
.B(n_381),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g408 ( 
.A1(n_380),
.A2(n_344),
.B(n_351),
.Y(n_408)
);

OAI322xp33_ASAP7_75t_L g409 ( 
.A1(n_386),
.A2(n_324),
.A3(n_337),
.B1(n_335),
.B2(n_307),
.C1(n_249),
.C2(n_303),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_383),
.Y(n_411)
);

AOI221xp5_ASAP7_75t_L g412 ( 
.A1(n_379),
.A2(n_358),
.B1(n_237),
.B2(n_240),
.C(n_307),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_392),
.B(n_391),
.Y(n_414)
);

AOI21xp33_ASAP7_75t_L g415 ( 
.A1(n_407),
.A2(n_299),
.B(n_309),
.Y(n_415)
);

AOI221xp5_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_387),
.B1(n_358),
.B2(n_240),
.C(n_237),
.Y(n_416)
);

AOI211xp5_ASAP7_75t_L g417 ( 
.A1(n_409),
.A2(n_387),
.B(n_384),
.C(n_373),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

AOI211xp5_ASAP7_75t_L g419 ( 
.A1(n_397),
.A2(n_299),
.B(n_309),
.C(n_307),
.Y(n_419)
);

OAI311xp33_ASAP7_75t_L g420 ( 
.A1(n_400),
.A2(n_249),
.A3(n_303),
.B1(n_237),
.C1(n_240),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_214),
.Y(n_421)
);

A2O1A1O1Ixp25_ASAP7_75t_L g422 ( 
.A1(n_396),
.A2(n_257),
.B(n_284),
.C(n_273),
.D(n_304),
.Y(n_422)
);

OAI211xp5_ASAP7_75t_SL g423 ( 
.A1(n_401),
.A2(n_244),
.B(n_245),
.C(n_236),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_394),
.A2(n_340),
.B1(n_331),
.B2(n_321),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_290),
.Y(n_426)
);

AOI221xp5_ASAP7_75t_L g427 ( 
.A1(n_403),
.A2(n_340),
.B1(n_331),
.B2(n_325),
.C(n_239),
.Y(n_427)
);

OAI211xp5_ASAP7_75t_L g428 ( 
.A1(n_405),
.A2(n_302),
.B(n_238),
.C(n_232),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_302),
.B(n_310),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_340),
.B1(n_331),
.B2(n_325),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_L g431 ( 
.A1(n_412),
.A2(n_325),
.B1(n_249),
.B2(n_252),
.Y(n_431)
);

AO221x1_ASAP7_75t_L g432 ( 
.A1(n_425),
.A2(n_413),
.B1(n_410),
.B2(n_393),
.C(n_258),
.Y(n_432)
);

NOR4xp25_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_395),
.C(n_258),
.D(n_196),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_428),
.C(n_427),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_290),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_419),
.B(n_310),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_290),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_L g438 ( 
.A1(n_423),
.A2(n_310),
.B(n_290),
.Y(n_438)
);

OAI211xp5_ASAP7_75t_SL g439 ( 
.A1(n_429),
.A2(n_236),
.B(n_244),
.C(n_245),
.Y(n_439)
);

AOI211xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_310),
.B(n_201),
.C(n_290),
.Y(n_440)
);

NAND4xp25_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_238),
.C(n_310),
.D(n_244),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_L g442 ( 
.A1(n_422),
.A2(n_241),
.B1(n_252),
.B2(n_258),
.Y(n_442)
);

NAND4xp25_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_424),
.C(n_418),
.D(n_426),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_443),
.Y(n_444)
);

NAND4xp75_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_420),
.C(n_431),
.D(n_250),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_238),
.C(n_258),
.Y(n_446)
);

AND3x4_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_310),
.C(n_290),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_238),
.Y(n_448)
);

NOR2x1p5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_238),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_440),
.Y(n_450)
);

NAND4xp25_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_236),
.C(n_244),
.D(n_245),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_302),
.Y(n_452)
);

NAND4xp75_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_250),
.C(n_202),
.D(n_302),
.Y(n_453)
);

NAND4xp25_ASAP7_75t_SL g454 ( 
.A(n_439),
.B(n_257),
.C(n_236),
.D(n_244),
.Y(n_454)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_302),
.C(n_211),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_302),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_202),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_SL g458 ( 
.A(n_447),
.B(n_261),
.C(n_260),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_241),
.Y(n_459)
);

NOR3xp33_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_258),
.C(n_199),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_257),
.Y(n_461)
);

NOR4xp25_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_196),
.C(n_199),
.D(n_227),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_SL g463 ( 
.A(n_446),
.B(n_261),
.C(n_260),
.Y(n_463)
);

NAND4xp75_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_250),
.C(n_227),
.D(n_211),
.Y(n_464)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_445),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_457),
.Y(n_468)
);

AND2x2_ASAP7_75t_SL g469 ( 
.A(n_462),
.B(n_452),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_460),
.B(n_454),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_468),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_467),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_466),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_469),
.A2(n_458),
.B1(n_464),
.B2(n_457),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_471),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_474),
.A2(n_469),
.B1(n_470),
.B2(n_465),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_477),
.A2(n_476),
.B(n_475),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_476),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_478),
.A2(n_470),
.B(n_466),
.Y(n_480)
);

AO21x2_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_479),
.B(n_463),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_481),
.A2(n_453),
.B1(n_239),
.B2(n_250),
.Y(n_482)
);


endmodule