module real_jpeg_30482_n_27 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_191, n_10, n_186, n_9, n_12, n_24, n_189, n_187, n_6, n_190, n_194, n_183, n_192, n_23, n_11, n_14, n_25, n_195, n_7, n_22, n_18, n_3, n_193, n_5, n_4, n_1, n_26, n_184, n_20, n_19, n_16, n_15, n_13, n_27);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_191;
input n_10;
input n_186;
input n_9;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_194;
input n_183;
input n_192;
input n_23;
input n_11;
input n_14;
input n_25;
input n_195;
input n_7;
input n_22;
input n_18;
input n_3;
input n_193;
input n_5;
input n_4;
input n_1;
input n_26;
input n_184;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_80;
wire n_32;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_0),
.A2(n_91),
.A3(n_93),
.B1(n_99),
.B2(n_161),
.C1(n_163),
.C2(n_193),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_1),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_1),
.B(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_2),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_6),
.Y(n_172)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_38),
.B1(n_40),
.B2(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_9),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_74),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_13),
.B(n_101),
.Y(n_159)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_14),
.B(n_79),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_15),
.B(n_69),
.Y(n_178)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_16),
.A2(n_19),
.B1(n_121),
.B2(n_125),
.C(n_129),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_16),
.B(n_121),
.C(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_18),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_18),
.B(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_19),
.Y(n_131)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_123),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_36),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_34),
.Y(n_154)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_35),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_82),
.B(n_166),
.Y(n_36)
);

NAND4xp25_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_47),
.C(n_72),
.D(n_77),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_44),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_56),
.C(n_62),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_49),
.B(n_176),
.C(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_50),
.B(n_55),
.Y(n_170)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g174 ( 
.A1(n_56),
.A2(n_64),
.A3(n_175),
.B1(n_178),
.B2(n_179),
.C1(n_180),
.C2(n_195),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_57),
.Y(n_173)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_63),
.A2(n_169),
.A3(n_170),
.B1(n_171),
.B2(n_174),
.C(n_194),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_73),
.A2(n_168),
.B(n_181),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI31xp67_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_110),
.A3(n_148),
.B(n_156),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_98),
.C(n_106),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_157),
.B(n_160),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_86),
.B(n_106),
.C(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_184),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_98),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_141),
.C(n_142),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_133),
.B(n_140),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B1(n_131),
.B2(n_132),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_189),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_139),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_183),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_185),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_186),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_187),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_188),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_190),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_191),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_192),
.Y(n_151)
);


endmodule