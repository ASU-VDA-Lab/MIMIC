module fake_jpeg_28155_n_243 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx9p33_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_16),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_20),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_63),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_19),
.B(n_22),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_34),
.B1(n_27),
.B2(n_18),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_80),
.B1(n_32),
.B2(n_31),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_36),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_34),
.B1(n_19),
.B2(n_22),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx12f_ASAP7_75t_SL g85 ( 
.A(n_55),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_20),
.B(n_35),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_33),
.Y(n_133)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_20),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_28),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_28),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_65),
.B1(n_60),
.B2(n_56),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_126),
.B1(n_135),
.B2(n_97),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_65),
.B1(n_56),
.B2(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_26),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_21),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_25),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_75),
.B1(n_52),
.B2(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_25),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_128),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_75),
.B1(n_108),
.B2(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_106),
.B1(n_88),
.B2(n_94),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_135),
.B1(n_122),
.B2(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_110),
.C(n_107),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_147),
.C(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_158),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_155),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_92),
.B1(n_88),
.B2(n_85),
.Y(n_146)
);

XOR2x2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_95),
.C(n_90),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_35),
.B(n_33),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_26),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_117),
.C(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_160),
.Y(n_175)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_131),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_169),
.B(n_1),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_158),
.B1(n_160),
.B2(n_144),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_125),
.B(n_131),
.C(n_122),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_174),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_127),
.B(n_35),
.C(n_92),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_140),
.B1(n_138),
.B2(n_141),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_199),
.B(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_196),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_163),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_193),
.B1(n_172),
.B2(n_171),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_142),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_137),
.B1(n_141),
.B2(n_151),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_152),
.C(n_156),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_169),
.C(n_170),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_167),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_197),
.B(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_0),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_163),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_205),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_169),
.C(n_170),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_208),
.B(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_211),
.C(n_194),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_171),
.B(n_169),
.C(n_166),
.D(n_162),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_164),
.C(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_192),
.B(n_195),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_188),
.C(n_193),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_218),
.C(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_197),
.C(n_184),
.Y(n_218)
);

OAI21x1_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_183),
.B(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_183),
.B(n_173),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_201),
.C(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_228),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_208),
.B(n_212),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_183),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_1),
.B(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_15),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_217),
.A3(n_208),
.B1(n_15),
.B2(n_13),
.C1(n_9),
.C2(n_6),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_234),
.B(n_235),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_225),
.B1(n_224),
.B2(n_4),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_223),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_232),
.B(n_7),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_5),
.C(n_7),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_239),
.Y(n_243)
);


endmodule