module real_aes_16824_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_93;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_0), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_1), .A2(n_5), .B1(n_577), .B2(n_582), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_1), .A2(n_5), .B1(n_621), .B2(n_624), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_2), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g552 ( .A(n_2), .Y(n_552) );
INVx1_ASAP7_75t_L g505 ( .A(n_3), .Y(n_505) );
BUFx3_ASAP7_75t_L g172 ( .A(n_4), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_6), .B(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_6), .Y(n_675) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_7), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_8), .B(n_143), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_9), .B(n_107), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_10), .A2(n_64), .B1(n_140), .B2(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g469 ( .A(n_11), .Y(n_469) );
INVx1_ASAP7_75t_L g475 ( .A(n_11), .Y(n_475) );
INVx1_ASAP7_75t_L g566 ( .A(n_12), .Y(n_566) );
INVx2_ASAP7_75t_L g460 ( .A(n_13), .Y(n_460) );
OAI21x1_ASAP7_75t_L g110 ( .A1(n_14), .A2(n_34), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g470 ( .A(n_15), .Y(n_470) );
INVx1_ASAP7_75t_L g492 ( .A(n_16), .Y(n_492) );
INVx1_ASAP7_75t_L g462 ( .A(n_17), .Y(n_462) );
BUFx2_ASAP7_75t_L g672 ( .A(n_18), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_19), .B(n_116), .Y(n_196) );
OAI211xp5_ASAP7_75t_L g557 ( .A1(n_20), .A2(n_558), .B(n_559), .C(n_565), .Y(n_557) );
INVx1_ASAP7_75t_L g619 ( .A(n_20), .Y(n_619) );
INVx1_ASAP7_75t_L g478 ( .A(n_21), .Y(n_478) );
AO32x1_ASAP7_75t_L g134 ( .A1(n_22), .A2(n_135), .A3(n_136), .B1(n_144), .B2(n_146), .Y(n_134) );
AO32x2_ASAP7_75t_L g250 ( .A1(n_22), .A2(n_135), .A3(n_136), .B1(n_144), .B2(n_146), .Y(n_250) );
INVx1_ASAP7_75t_L g495 ( .A(n_23), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_24), .A2(n_38), .B1(n_116), .B2(n_117), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_25), .A2(n_69), .B1(n_140), .B2(n_141), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_26), .B(n_182), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_27), .B(n_207), .Y(n_228) );
INVx2_ASAP7_75t_L g459 ( .A(n_28), .Y(n_459) );
INVx1_ASAP7_75t_L g503 ( .A(n_28), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_29), .A2(n_52), .B1(n_141), .B2(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_30), .Y(n_666) );
INVx2_ASAP7_75t_L g649 ( .A(n_31), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_32), .B(n_230), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g585 ( .A1(n_33), .A2(n_45), .B1(n_586), .B2(n_590), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_33), .A2(n_45), .B1(n_601), .B2(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g484 ( .A(n_35), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_36), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_37), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_39), .A2(n_59), .B1(n_125), .B2(n_207), .Y(n_206) );
BUFx3_ASAP7_75t_L g467 ( .A(n_40), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_41), .A2(n_61), .B1(n_140), .B2(n_143), .Y(n_168) );
BUFx3_ASAP7_75t_L g691 ( .A(n_41), .Y(n_691) );
AND2x4_ASAP7_75t_L g85 ( .A(n_42), .B(n_86), .Y(n_85) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_42), .Y(n_635) );
INVx1_ASAP7_75t_L g111 ( .A(n_43), .Y(n_111) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_44), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_46), .B(n_140), .Y(n_178) );
INVx1_ASAP7_75t_L g86 ( .A(n_47), .Y(n_86) );
XOR2xp5_ASAP7_75t_L g448 ( .A(n_48), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_49), .B(n_146), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g121 ( .A1(n_50), .A2(n_122), .B(n_123), .C(n_126), .Y(n_121) );
NAND3xp33_ASAP7_75t_L g185 ( .A(n_51), .B(n_140), .C(n_184), .Y(n_185) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_53), .Y(n_523) );
AND2x2_ASAP7_75t_L g129 ( .A(n_54), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_55), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_56), .A2(n_73), .B1(n_125), .B2(n_143), .Y(n_209) );
INVx2_ASAP7_75t_L g95 ( .A(n_57), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_58), .B(n_199), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_60), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_62), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_62), .Y(n_661) );
BUFx3_ASAP7_75t_L g515 ( .A(n_63), .Y(n_515) );
INVx1_ASAP7_75t_L g581 ( .A(n_63), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_65), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g457 ( .A(n_66), .Y(n_457) );
INVx1_ASAP7_75t_L g502 ( .A(n_66), .Y(n_502) );
INVx2_ASAP7_75t_L g513 ( .A(n_66), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_67), .A2(n_77), .B1(n_117), .B2(n_141), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_68), .B(n_207), .Y(n_225) );
BUFx2_ASAP7_75t_L g665 ( .A(n_68), .Y(n_665) );
BUFx2_ASAP7_75t_L g677 ( .A(n_70), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_71), .B(n_107), .Y(n_231) );
INVx2_ASAP7_75t_L g660 ( .A(n_72), .Y(n_660) );
INVx1_ASAP7_75t_L g508 ( .A(n_74), .Y(n_508) );
INVx1_ASAP7_75t_L g570 ( .A(n_75), .Y(n_570) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_75), .A2(n_506), .B(n_606), .C(n_610), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_76), .Y(n_193) );
INVx1_ASAP7_75t_L g685 ( .A(n_77), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_96), .B(n_447), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_87), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
BUFx10_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g128 ( .A(n_85), .Y(n_128) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
AO31x2_ASAP7_75t_L g147 ( .A1(n_85), .A2(n_148), .A3(n_149), .B(n_155), .Y(n_147) );
BUFx10_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_86), .Y(n_637) );
AOI21xp5_ASAP7_75t_SL g693 ( .A1(n_87), .A2(n_636), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_94), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_93), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
INVx1_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
INVx1_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
INVx2_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_93), .Y(n_180) );
INVx1_ASAP7_75t_L g195 ( .A(n_93), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_94), .A2(n_137), .B1(n_139), .B2(n_142), .Y(n_136) );
INVx6_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_94), .A2(n_152), .B1(n_168), .B2(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_94), .A2(n_178), .B(n_179), .Y(n_177) );
BUFx8_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g120 ( .A(n_95), .Y(n_120) );
INVx2_ASAP7_75t_L g127 ( .A(n_95), .Y(n_127) );
INVx1_ASAP7_75t_L g138 ( .A(n_95), .Y(n_138) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND4xp75_ASAP7_75t_L g97 ( .A(n_98), .B(n_321), .C(n_375), .D(n_419), .Y(n_97) );
NOR2x1_ASAP7_75t_L g98 ( .A(n_99), .B(n_274), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_100), .B(n_240), .Y(n_99) );
O2A1O1Ixp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_157), .B(n_161), .C(n_213), .Y(n_100) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_132), .Y(n_101) );
AND2x2_ASAP7_75t_L g291 ( .A(n_102), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g280 ( .A(n_103), .B(n_216), .Y(n_280) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_104), .Y(n_246) );
AND2x2_ASAP7_75t_L g295 ( .A(n_104), .B(n_147), .Y(n_295) );
INVx1_ASAP7_75t_L g307 ( .A(n_104), .Y(n_307) );
INVx1_ASAP7_75t_L g405 ( .A(n_104), .Y(n_405) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g159 ( .A(n_105), .Y(n_159) );
AOI21x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_112), .B(n_129), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g131 ( .A(n_109), .Y(n_131) );
INVx2_ASAP7_75t_L g175 ( .A(n_109), .Y(n_175) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_121), .B(n_128), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_114), .B(n_119), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B1(n_117), .B2(n_118), .Y(n_114) );
INVx2_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx1_ASAP7_75t_L g201 ( .A(n_117), .Y(n_201) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g208 ( .A(n_120), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx2_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g200 ( .A(n_127), .Y(n_200) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_131), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g233 ( .A(n_133), .B(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_147), .Y(n_133) );
AND2x2_ASAP7_75t_L g160 ( .A(n_134), .B(n_147), .Y(n_160) );
INVx1_ASAP7_75t_L g273 ( .A(n_134), .Y(n_273) );
INVx1_ASAP7_75t_L g384 ( .A(n_134), .Y(n_384) );
INVx4_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
BUFx3_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_135), .B(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_135), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
INVx2_ASAP7_75t_SL g222 ( .A(n_135), .Y(n_222) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_137), .A2(n_193), .B(n_194), .C(n_196), .Y(n_192) );
BUFx4f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx2_ASAP7_75t_SL g207 ( .A(n_140), .Y(n_207) );
INVx2_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
INVx3_ASAP7_75t_L g230 ( .A(n_143), .Y(n_230) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_144), .A2(n_224), .B(n_227), .Y(n_223) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_SL g210 ( .A(n_145), .Y(n_210) );
INVx2_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
INVx3_ASAP7_75t_L g216 ( .A(n_147), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_147), .B(n_220), .Y(n_271) );
AND2x2_ASAP7_75t_L g306 ( .A(n_147), .B(n_307), .Y(n_306) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_148), .A2(n_205), .A3(n_210), .B(n_211), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B1(n_153), .B2(n_154), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_152), .A2(n_206), .B1(n_208), .B2(n_209), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_152), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_225), .B(n_226), .Y(n_224) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
INVx1_ASAP7_75t_L g346 ( .A(n_158), .Y(n_346) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g215 ( .A(n_159), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_159), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g248 ( .A(n_159), .Y(n_248) );
OR2x2_ASAP7_75t_L g312 ( .A(n_159), .B(n_220), .Y(n_312) );
OR2x2_ASAP7_75t_L g383 ( .A(n_159), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g320 ( .A(n_160), .Y(n_320) );
AND2x2_ASAP7_75t_L g372 ( .A(n_160), .B(n_235), .Y(n_372) );
AND2x2_ASAP7_75t_L g429 ( .A(n_160), .B(n_346), .Y(n_429) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_187), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_162), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g438 ( .A(n_162), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_173), .Y(n_162) );
INVx2_ASAP7_75t_L g239 ( .A(n_163), .Y(n_239) );
AND2x2_ASAP7_75t_L g264 ( .A(n_163), .B(n_243), .Y(n_264) );
AND2x2_ASAP7_75t_L g334 ( .A(n_163), .B(n_204), .Y(n_334) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g288 ( .A(n_164), .Y(n_288) );
AOI31xp67_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .A3(n_167), .B(n_170), .Y(n_164) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_166), .A2(n_177), .B(n_181), .Y(n_176) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_166), .A2(n_192), .B(n_197), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g242 ( .A(n_173), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g303 ( .A(n_173), .B(n_189), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_186), .Y(n_173) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_174), .A2(n_176), .B(n_186), .Y(n_259) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_185), .Y(n_181) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g310 ( .A(n_188), .B(n_287), .Y(n_310) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
INVx2_ASAP7_75t_SL g232 ( .A(n_189), .Y(n_232) );
BUFx2_ASAP7_75t_L g285 ( .A(n_189), .Y(n_285) );
INVx1_ASAP7_75t_L g357 ( .A(n_189), .Y(n_357) );
AND2x2_ASAP7_75t_L g390 ( .A(n_189), .B(n_238), .Y(n_390) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_203), .Y(n_189) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_190), .A2(n_191), .B(n_203), .Y(n_243) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_197) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g218 ( .A(n_204), .Y(n_218) );
INVx1_ASAP7_75t_L g238 ( .A(n_204), .Y(n_238) );
INVx1_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
AND2x2_ASAP7_75t_L g356 ( .A(n_204), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g397 ( .A(n_204), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g413 ( .A(n_204), .B(n_398), .Y(n_413) );
AND2x2_ASAP7_75t_L g439 ( .A(n_204), .B(n_243), .Y(n_439) );
OAI32xp33_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .A3(n_232), .B1(n_233), .B2(n_236), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_215), .B(n_380), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_215), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g249 ( .A(n_216), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g351 ( .A(n_216), .Y(n_351) );
INVx1_ASAP7_75t_L g411 ( .A(n_216), .Y(n_411) );
INVx1_ASAP7_75t_L g349 ( .A(n_217), .Y(n_349) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_SL g253 ( .A(n_218), .Y(n_253) );
AND2x2_ASAP7_75t_L g342 ( .A(n_218), .B(n_257), .Y(n_342) );
AND2x2_ASAP7_75t_L g410 ( .A(n_219), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g235 ( .A(n_220), .Y(n_235) );
AND2x2_ASAP7_75t_L g245 ( .A(n_220), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g281 ( .A(n_220), .Y(n_281) );
AND2x2_ASAP7_75t_L g292 ( .A(n_220), .B(n_250), .Y(n_292) );
AND2x2_ASAP7_75t_L g316 ( .A(n_220), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g326 ( .A(n_220), .B(n_317), .Y(n_326) );
INVxp67_ASAP7_75t_L g380 ( .A(n_220), .Y(n_380) );
BUFx2_ASAP7_75t_L g392 ( .A(n_220), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_220), .Y(n_396) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_231), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_232), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g388 ( .A(n_232), .Y(n_388) );
AND2x2_ASAP7_75t_L g296 ( .A(n_235), .B(n_273), .Y(n_296) );
AND2x2_ASAP7_75t_L g425 ( .A(n_235), .B(n_249), .Y(n_425) );
OAI22xp5_ASAP7_75t_SL g313 ( .A1(n_236), .A2(n_314), .B1(n_318), .B2(n_319), .Y(n_313) );
O2A1O1Ixp5_ASAP7_75t_R g387 ( .A1(n_236), .A2(n_388), .B(n_389), .C(n_391), .Y(n_387) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g241 ( .A(n_237), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
INVx1_ASAP7_75t_L g298 ( .A(n_239), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_239), .B(n_268), .Y(n_374) );
AND2x2_ASAP7_75t_L g386 ( .A(n_239), .B(n_257), .Y(n_386) );
AOI222xp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .B1(n_247), .B2(n_251), .C1(n_261), .C2(n_269), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_241), .A2(n_283), .B1(n_361), .B2(n_422), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_241), .A2(n_305), .B1(n_441), .B2(n_443), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_242), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_242), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g416 ( .A(n_242), .Y(n_416) );
INVx1_ASAP7_75t_L g446 ( .A(n_242), .Y(n_446) );
INVx1_ASAP7_75t_L g260 ( .A(n_243), .Y(n_260) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g315 ( .A(n_246), .Y(n_315) );
AOI321xp33_ASAP7_75t_L g393 ( .A1(n_247), .A2(n_291), .A3(n_394), .B1(n_399), .B2(n_400), .C(n_401), .Y(n_393) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
OR2x2_ASAP7_75t_L g325 ( .A(n_248), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g345 ( .A(n_249), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g317 ( .A(n_250), .Y(n_317) );
NAND2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
OR2x2_ASAP7_75t_L g318 ( .A(n_253), .B(n_287), .Y(n_318) );
AND2x2_ASAP7_75t_L g338 ( .A(n_253), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g428 ( .A(n_254), .Y(n_428) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g359 ( .A(n_256), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g268 ( .A(n_258), .Y(n_268) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g287 ( .A(n_259), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_262), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_264), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g399 ( .A(n_268), .Y(n_399) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_270), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g332 ( .A(n_271), .Y(n_332) );
INVx1_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
INVx2_ASAP7_75t_L g364 ( .A(n_273), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_299), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_283), .B(n_289), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_278), .B(n_282), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_279), .A2(n_366), .B1(n_416), .B2(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g381 ( .A(n_280), .Y(n_381) );
AND2x2_ASAP7_75t_L g305 ( .A(n_281), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g370 ( .A(n_281), .Y(n_370) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g350 ( .A(n_285), .B(n_286), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_285), .B(n_334), .Y(n_366) );
AND2x2_ASAP7_75t_L g412 ( .A(n_285), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_286), .B(n_390), .Y(n_427) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
INVx1_ASAP7_75t_L g398 ( .A(n_288), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B(n_297), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g360 ( .A(n_292), .B(n_315), .Y(n_360) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_295), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g369 ( .A(n_295), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_298), .B(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_313), .Y(n_299) );
OAI21xp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B(n_308), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_301), .A2(n_368), .B1(n_371), .B2(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AOI311xp33_ASAP7_75t_L g401 ( .A1(n_303), .A2(n_402), .A3(n_403), .B(n_406), .C(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g329 ( .A(n_306), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_306), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g400 ( .A(n_310), .Y(n_400) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g406 ( .A(n_316), .Y(n_406) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_320), .Y(n_423) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_347), .Y(n_321) );
NAND3xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .C(n_335), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AO21x1_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B(n_333), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AO221x1_ASAP7_75t_L g408 ( .A1(n_329), .A2(n_409), .B1(n_412), .B2(n_414), .C(n_415), .Y(n_408) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B(n_343), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_351), .B(n_352), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g402 ( .A(n_351), .Y(n_402) );
AOI221x1_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_360), .B1(n_361), .B2(n_365), .C(n_367), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_358), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g385 ( .A(n_356), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AO22x1_ASAP7_75t_L g432 ( .A1(n_360), .A2(n_433), .B1(n_435), .B2(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g409 ( .A(n_363), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_364), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp33_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_408), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_393), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_385), .B(n_387), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .C(n_383), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
AND2x2_ASAP7_75t_L g404 ( .A(n_384), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g414 ( .A(n_390), .B(n_399), .Y(n_414) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_396), .B(n_404), .Y(n_442) );
INVx2_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
AND2x2_ASAP7_75t_L g433 ( .A(n_413), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_430), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_426), .B1(n_428), .B2(n_429), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_440), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_633), .B1(n_638), .B2(n_686), .C(n_687), .Y(n_447) );
INVx1_ASAP7_75t_L g686 ( .A(n_449), .Y(n_686) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_556), .C(n_599), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_509), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_461), .A3(n_477), .B1(n_489), .B2(n_496), .B3(n_504), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g550 ( .A(n_455), .Y(n_550) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_455), .Y(n_632) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g598 ( .A(n_456), .Y(n_598) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g654 ( .A(n_458), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_460), .Y(n_458) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_459), .Y(n_630) );
INVx1_ASAP7_75t_L g648 ( .A(n_459), .Y(n_648) );
INVx3_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
BUFx3_ASAP7_75t_L g614 ( .A(n_460), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_470), .B2(n_471), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g516 ( .A1(n_462), .A2(n_505), .B1(n_517), .B2(n_525), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_463), .A2(n_505), .B1(n_506), .B2(n_508), .Y(n_504) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx4f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x4_ASAP7_75t_L g601 ( .A(n_466), .B(n_500), .Y(n_601) );
OR2x4_ASAP7_75t_L g623 ( .A(n_466), .B(n_604), .Y(n_623) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_467), .Y(n_476) );
INVx2_ASAP7_75t_L g483 ( .A(n_467), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_467), .B(n_475), .Y(n_488) );
AND2x4_ASAP7_75t_L g608 ( .A(n_467), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g482 ( .A(n_469), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_470), .A2(n_508), .B1(n_542), .B2(n_545), .Y(n_541) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g507 ( .A(n_473), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
BUFx2_ASAP7_75t_L g618 ( .A(n_474), .Y(n_618) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g609 ( .A(n_475), .Y(n_609) );
BUFx2_ASAP7_75t_L g615 ( .A(n_476), .Y(n_615) );
INVx2_ASAP7_75t_L g646 ( .A(n_476), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_484), .B2(n_485), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_478), .A2(n_492), .B1(n_532), .B2(n_536), .Y(n_531) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g603 ( .A(n_480), .B(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g491 ( .A(n_481), .Y(n_491) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_484), .A2(n_495), .B1(n_517), .B2(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g494 ( .A(n_487), .Y(n_494) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g626 ( .A(n_488), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_492), .B1(n_493), .B2(n_495), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND3x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .C(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g604 ( .A(n_500), .Y(n_604) );
AND2x4_ASAP7_75t_L g607 ( .A(n_500), .B(n_608), .Y(n_607) );
OR2x6_ASAP7_75t_L g625 ( .A(n_500), .B(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g647 ( .A(n_500), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI33xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_516), .A3(n_531), .B1(n_541), .B2(n_546), .B3(n_553), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g551 ( .A(n_515), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
BUFx2_ASAP7_75t_L g568 ( .A(n_515), .Y(n_568) );
AND2x4_ASAP7_75t_L g573 ( .A(n_515), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g579 ( .A(n_521), .Y(n_579) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g530 ( .A(n_523), .Y(n_530) );
INVx2_ASAP7_75t_L g535 ( .A(n_523), .Y(n_535) );
NAND2x1_ASAP7_75t_L g540 ( .A(n_523), .B(n_524), .Y(n_540) );
AND2x2_ASAP7_75t_L g564 ( .A(n_523), .B(n_524), .Y(n_564) );
INVx1_ASAP7_75t_L g575 ( .A(n_523), .Y(n_575) );
AND2x2_ASAP7_75t_L g592 ( .A(n_523), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_524), .B(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g534 ( .A(n_524), .B(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g569 ( .A(n_524), .Y(n_569) );
INVx2_ASAP7_75t_L g593 ( .A(n_524), .Y(n_593) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g555 ( .A(n_526), .Y(n_555) );
INVx4_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx8_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g584 ( .A(n_528), .B(n_568), .Y(n_584) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g544 ( .A(n_534), .Y(n_544) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx4f_ASAP7_75t_L g545 ( .A(n_539), .Y(n_545) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_539), .Y(n_558) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g596 ( .A(n_552), .Y(n_596) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI31xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_576), .A3(n_585), .B(n_594), .Y(n_556) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVxp67_ASAP7_75t_L g589 ( .A(n_562), .Y(n_589) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_570), .B2(n_571), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_566), .A2(n_611), .B1(n_616), .B2(n_619), .Y(n_610) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x6_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x6_ASAP7_75t_L g588 ( .A(n_579), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g591 ( .A(n_580), .B(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx3_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OAI31xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_605), .A3(n_620), .B(n_627), .Y(n_599) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
CKINVDCx8_ASAP7_75t_R g606 ( .A(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AND2x4_ASAP7_75t_L g617 ( .A(n_613), .B(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx4f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g656 ( .A(n_635), .Y(n_656) );
BUFx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_637), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g694 ( .A(n_637), .B(n_656), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_657), .B1(n_679), .B2(n_684), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx12f_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx3_ASAP7_75t_L g689 ( .A(n_641), .Y(n_689) );
BUFx8_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_649), .B(n_650), .C(n_655), .Y(n_642) );
AND2x2_ASAP7_75t_L g683 ( .A(n_643), .B(n_650), .Y(n_683) );
INVx4_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x6_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_645), .B(n_651), .C(n_654), .Y(n_650) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx3_ASAP7_75t_L g653 ( .A(n_649), .Y(n_653) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g682 ( .A(n_655), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_657), .A2(n_684), .B1(n_689), .B2(n_690), .Y(n_688) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_670), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_663), .B1(n_664), .B2(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g669 ( .A(n_659), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_660), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_666), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_675), .Y(n_678) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g690 ( .A(n_681), .Y(n_690) );
OR2x6_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_688), .B1(n_691), .B2(n_692), .Y(n_687) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
endmodule