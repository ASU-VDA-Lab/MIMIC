module fake_ariane_932_n_2236 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2236);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2236;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_967;
wire n_274;
wire n_437;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_439;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_94),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_103),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_17),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_34),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_126),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_125),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_18),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_52),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_96),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_85),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_90),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_82),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_6),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_139),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_89),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_141),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_35),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_140),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_37),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_100),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_81),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_158),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_67),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_164),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_108),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_93),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_222),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_62),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_114),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_132),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_147),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_178),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_107),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_197),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_171),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_37),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_43),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_23),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_119),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_137),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_55),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_0),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_86),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_150),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_130),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_131),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_199),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_151),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_162),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_128),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_28),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_30),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_149),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_98),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_179),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_156),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_214),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_204),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_75),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_201),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_29),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_117),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_143),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_64),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_124),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_161),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_198),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_11),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_170),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_31),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_180),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_73),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_76),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_72),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_26),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_174),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_67),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_167),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_136),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_55),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_19),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_16),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_6),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_207),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_175),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_97),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_11),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_78),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_123),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_41),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_138),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_166),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_44),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_25),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_79),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_58),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_0),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_14),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_92),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_194),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_46),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_189),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_228),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_193),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_88),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_106),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_219),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_2),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_74),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_15),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_3),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_154),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_95),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_51),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_217),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_22),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_80),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_185),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_43),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_115),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_34),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_15),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_66),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_3),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_187),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_112),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_48),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_17),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_72),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_210),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_153),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_24),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_122),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_26),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_28),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_33),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_35),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_9),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_127),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_46),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_144),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_205),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_208),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_29),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_7),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_45),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_220),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_61),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_118),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_49),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_102),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_69),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_25),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_213),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_116),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_18),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_48),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_73),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_227),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_64),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_195),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_33),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_8),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_27),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_172),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_49),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_83),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_23),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_16),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_71),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_56),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_110),
.Y(n_424)
);

BUFx5_ASAP7_75t_L g425 ( 
.A(n_184),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_84),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_188),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_52),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_186),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_224),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_135),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_62),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_182),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_142),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_77),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_57),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_160),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_22),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_109),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_111),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_216),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_53),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_91),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_1),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_203),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_9),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_53),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_121),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_176),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_234),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_245),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_334),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_234),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_334),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_334),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_334),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_334),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_423),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_334),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_334),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_292),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_297),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_297),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_237),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_316),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_282),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_269),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_379),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_233),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_233),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_334),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_237),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_295),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_375),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_249),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_239),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_249),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_340),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_239),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_356),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_274),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_230),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_274),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_294),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_294),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_240),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_304),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_365),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_304),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_321),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_352),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_385),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_352),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_277),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_242),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_364),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_240),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_364),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_369),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_235),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_266),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_251),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_255),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_267),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_281),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_236),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_283),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_302),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_278),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_300),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_279),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_285),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_324),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_244),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_326),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_332),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_339),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_286),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_314),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_342),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_360),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_289),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_241),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_301),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_366),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_373),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_384),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_387),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_397),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_400),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_318),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_320),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_246),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_248),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_252),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_404),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_269),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_241),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_322),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_444),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_260),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_253),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_328),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_269),
.Y(n_549)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_302),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_264),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_335),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_345),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_271),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_290),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_291),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_298),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_346),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_299),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_310),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_266),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_349),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_353),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_362),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_315),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_317),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_243),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_333),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_319),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_302),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_466),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_513),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_508),
.B(n_426),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_311),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_467),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_495),
.B(n_229),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_452),
.B(n_269),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_473),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_468),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_454),
.Y(n_581)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_455),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_481),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_493),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_467),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_465),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_467),
.Y(n_592)
);

INVxp33_ASAP7_75t_SL g593 ( 
.A(n_509),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_541),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_561),
.B(n_325),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_SL g599 ( 
.A(n_570),
.B(n_243),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_541),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_541),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_514),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_456),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_549),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_547),
.B(n_550),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_457),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_457),
.B(n_269),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_570),
.B(n_327),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_450),
.A2(n_371),
.B1(n_409),
.B2(n_350),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_472),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_549),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_461),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_459),
.B(n_357),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_549),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_459),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_460),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_469),
.B(n_311),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_460),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_471),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_471),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_462),
.B(n_329),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_476),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_478),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_521),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_482),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_537),
.B(n_236),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_463),
.B(n_336),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_482),
.Y(n_635)
);

AND2x2_ASAP7_75t_SL g636 ( 
.A(n_542),
.B(n_357),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_484),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

INVxp33_ASAP7_75t_SL g639 ( 
.A(n_526),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_485),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_508),
.B(n_337),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_508),
.B(n_341),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_L g643 ( 
.A(n_533),
.B(n_363),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_485),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_486),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_488),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_488),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_490),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_490),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_492),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_470),
.B(n_475),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_492),
.Y(n_653)
);

INVx6_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_494),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_483),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_494),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_497),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_497),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_499),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_451),
.B(n_306),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_499),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_500),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_500),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_623),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_636),
.B(n_537),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_656),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_574),
.B(n_545),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_656),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_613),
.A2(n_505),
.B1(n_542),
.B2(n_491),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_656),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_577),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_546),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_636),
.B(n_534),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_623),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_R g677 ( 
.A(n_606),
.B(n_453),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_573),
.B(n_464),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_623),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_583),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_L g681 ( 
.A(n_621),
.B(n_425),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_574),
.B(n_546),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_633),
.B(n_496),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_626),
.Y(n_684)
);

INVx8_ASAP7_75t_L g685 ( 
.A(n_633),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_621),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_583),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_626),
.Y(n_688)
);

XNOR2xp5_ASAP7_75t_L g689 ( 
.A(n_572),
.B(n_630),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_616),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_661),
.A2(n_498),
.B1(n_548),
.B2(n_544),
.Y(n_691)
);

CKINVDCx11_ASAP7_75t_R g692 ( 
.A(n_593),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_583),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_621),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_652),
.B(n_551),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_628),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_579),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_621),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_579),
.B(n_552),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_643),
.B(n_558),
.C(n_553),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_633),
.A2(n_491),
.B1(n_451),
.B2(n_622),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_632),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_599),
.B(n_563),
.C(n_562),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_581),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_632),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_581),
.B(n_564),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_584),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_SL g708 ( 
.A1(n_598),
.A2(n_569),
.B(n_554),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_584),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_596),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_632),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_628),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_622),
.A2(n_381),
.B1(n_247),
.B2(n_348),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_578),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_591),
.A2(n_510),
.B1(n_503),
.B2(n_480),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_596),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_603),
.B(n_347),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_603),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_607),
.Y(n_719)
);

NOR2x1p5_ASAP7_75t_L g720 ( 
.A(n_590),
.B(n_259),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_576),
.B(n_477),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_571),
.B(n_487),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_654),
.B(n_551),
.Y(n_723)
);

BUFx6f_ASAP7_75t_SL g724 ( 
.A(n_633),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_607),
.B(n_355),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_R g726 ( 
.A(n_586),
.B(n_479),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_654),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_654),
.B(n_554),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_602),
.B(n_567),
.C(n_525),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_654),
.B(n_555),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_654),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_629),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_608),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_608),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_620),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_641),
.B(n_555),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_620),
.B(n_358),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_629),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_631),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_631),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_652),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_637),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_637),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_588),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_632),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_642),
.B(n_556),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_612),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_644),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_644),
.Y(n_750)
);

INVx5_ASAP7_75t_L g751 ( 
.A(n_577),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_624),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_625),
.B(n_639),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_577),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_580),
.B(n_502),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_645),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_632),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_582),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_582),
.B(n_458),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_625),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_664),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_632),
.Y(n_763)
);

INVx6_ASAP7_75t_L g764 ( 
.A(n_635),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_647),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_635),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_647),
.B(n_357),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_635),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_649),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_635),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_635),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_635),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_649),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_664),
.Y(n_774)
);

BUFx6f_ASAP7_75t_SL g775 ( 
.A(n_582),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_611),
.B(n_556),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_640),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_640),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_627),
.B(n_504),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_617),
.A2(n_261),
.B1(n_416),
.B2(n_259),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_653),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_664),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_640),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_640),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_653),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_640),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_640),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_648),
.B(n_359),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_655),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_655),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_582),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_648),
.B(n_367),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_648),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_577),
.B(n_425),
.Y(n_794)
);

CKINVDCx16_ASAP7_75t_R g795 ( 
.A(n_614),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_634),
.B(n_416),
.C(n_261),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_577),
.B(n_425),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_664),
.B(n_557),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_638),
.B(n_557),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_638),
.Y(n_800)
);

INVxp33_ASAP7_75t_L g801 ( 
.A(n_648),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_648),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_577),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_648),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_658),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_638),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_658),
.Y(n_807)
);

AND2x6_ASAP7_75t_L g808 ( 
.A(n_658),
.B(n_357),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_614),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_665),
.B(n_496),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_658),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_658),
.A2(n_560),
.B1(n_565),
.B2(n_559),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_614),
.Y(n_813)
);

INVx8_ASAP7_75t_L g814 ( 
.A(n_577),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_658),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_614),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_646),
.B(n_559),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_660),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_646),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_660),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_577),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_660),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_660),
.B(n_378),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_646),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_650),
.B(n_560),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_660),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_660),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_610),
.B(n_425),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_762),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_748),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_682),
.B(n_565),
.Y(n_831)
);

BUFx5_ASAP7_75t_L g832 ( 
.A(n_803),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_762),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_727),
.B(n_663),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_782),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_669),
.B(n_489),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_697),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_782),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_682),
.B(n_566),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_714),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_669),
.B(n_568),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_727),
.B(n_663),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_669),
.B(n_678),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_742),
.B(n_566),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_816),
.B(n_506),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_707),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_707),
.Y(n_848)
);

BUFx8_ASAP7_75t_L g849 ( 
.A(n_775),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_727),
.B(n_663),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_697),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_755),
.B(n_511),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_667),
.B(n_569),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_704),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_674),
.B(n_650),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_709),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_755),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_710),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_704),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_675),
.A2(n_535),
.B1(n_536),
.B2(n_516),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_695),
.B(n_650),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_675),
.B(n_663),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_708),
.A2(n_657),
.B(n_659),
.C(n_651),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_748),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_753),
.A2(n_354),
.B1(n_231),
.B2(n_238),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_695),
.B(n_651),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_731),
.B(n_663),
.Y(n_868)
);

BUFx6f_ASAP7_75t_SL g869 ( 
.A(n_748),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_691),
.B(n_229),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_716),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_799),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_799),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_753),
.B(n_663),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_718),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_718),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_668),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_722),
.Y(n_878)
);

AO221x1_ASAP7_75t_L g879 ( 
.A1(n_671),
.A2(n_715),
.B1(n_780),
.B2(n_791),
.C(n_759),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_736),
.B(n_651),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_731),
.B(n_231),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_714),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_775),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_699),
.B(n_657),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_747),
.B(n_657),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_699),
.A2(n_518),
.B(n_519),
.C(n_517),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_670),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_745),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_745),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_719),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_689),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_706),
.B(n_665),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_776),
.B(n_659),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_726),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_706),
.B(n_665),
.Y(n_895)
);

BUFx5_ASAP7_75t_L g896 ( 
.A(n_803),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_779),
.B(n_659),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_731),
.B(n_238),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_722),
.B(n_690),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_779),
.B(n_662),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_719),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_774),
.B(n_662),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_724),
.A2(n_354),
.B1(n_250),
.B2(n_256),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_686),
.B(n_662),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_694),
.B(n_250),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_693),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_721),
.B(n_516),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_824),
.B(n_535),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_685),
.B(n_536),
.Y(n_909)
);

NAND2xp33_ASAP7_75t_L g910 ( 
.A(n_693),
.B(n_610),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_694),
.A2(n_698),
.B(n_734),
.C(n_733),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_685),
.B(n_684),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_796),
.B(n_420),
.C(n_418),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_729),
.B(n_420),
.C(n_418),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_685),
.B(n_501),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_816),
.B(n_512),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_672),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_688),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_685),
.B(n_696),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_698),
.B(n_693),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_712),
.B(n_501),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_L g922 ( 
.A(n_733),
.B(n_734),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_735),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_732),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_723),
.A2(n_432),
.B1(n_436),
.B2(n_421),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_692),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_814),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_738),
.B(n_740),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_741),
.B(n_232),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_702),
.B(n_254),
.Y(n_930)
);

BUFx5_ASAP7_75t_L g931 ( 
.A(n_803),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_743),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_700),
.B(n_368),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_735),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_SL g935 ( 
.A(n_677),
.B(n_421),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_744),
.B(n_258),
.Y(n_936)
);

AO22x2_ASAP7_75t_L g937 ( 
.A1(n_717),
.A2(n_528),
.B1(n_540),
.B2(n_517),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_724),
.B(n_374),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_749),
.B(n_750),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_702),
.B(n_254),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_756),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_728),
.A2(n_587),
.B(n_575),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_739),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_758),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_702),
.B(n_256),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_765),
.B(n_272),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_739),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_683),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_724),
.B(n_376),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_769),
.B(n_312),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_773),
.B(n_313),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_703),
.B(n_380),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_713),
.B(n_515),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_752),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_702),
.B(n_257),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_781),
.B(n_394),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_683),
.B(n_386),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_763),
.B(n_257),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_752),
.A2(n_311),
.B1(n_527),
.B2(n_528),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_785),
.B(n_399),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_789),
.B(n_262),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_763),
.B(n_262),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_790),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_817),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_825),
.Y(n_965)
);

AND2x2_ASAP7_75t_SL g966 ( 
.A(n_795),
.B(n_382),
.Y(n_966)
);

AND2x6_ASAP7_75t_L g967 ( 
.A(n_666),
.B(n_357),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_683),
.B(n_388),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_761),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_763),
.B(n_263),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_761),
.Y(n_971)
);

BUFx10_ASAP7_75t_L g972 ( 
.A(n_775),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_701),
.B(n_263),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_763),
.B(n_265),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_814),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_680),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_798),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_810),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_810),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_683),
.B(n_389),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_810),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_801),
.B(n_390),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_810),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_730),
.B(n_265),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_766),
.B(n_268),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_809),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_687),
.B(n_812),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_717),
.B(n_268),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_813),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_725),
.B(n_436),
.C(n_432),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_800),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_725),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_666),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_737),
.A2(n_427),
.B1(n_417),
.B2(n_429),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_720),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_737),
.B(n_417),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_766),
.B(n_427),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_806),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_676),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_918),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_SL g1001 ( 
.A1(n_966),
.A2(n_760),
.B1(n_442),
.B2(n_446),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_844),
.B(n_676),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_L g1003 ( 
.A(n_864),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_986),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_927),
.B(n_978),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_964),
.B(n_679),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_976),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_SL g1008 ( 
.A1(n_966),
.A2(n_442),
.B1(n_446),
.B2(n_438),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_927),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_836),
.A2(n_681),
.B1(n_805),
.B2(n_820),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_SL g1011 ( 
.A1(n_879),
.A2(n_447),
.B1(n_438),
.B2(n_396),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_899),
.B(n_766),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_883),
.B(n_814),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_927),
.Y(n_1014)
);

OAI21xp33_ASAP7_75t_SL g1015 ( 
.A1(n_928),
.A2(n_819),
.B(n_679),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_882),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_849),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_L g1018 ( 
.A(n_927),
.B(n_766),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_924),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_841),
.Y(n_1020)
);

BUFx8_ASAP7_75t_L g1021 ( 
.A(n_869),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_857),
.B(n_836),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_965),
.B(n_705),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_977),
.B(n_705),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_857),
.B(n_787),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_990),
.A2(n_792),
.B1(n_823),
.B2(n_788),
.Y(n_1026)
);

NAND2x2_ASAP7_75t_L g1027 ( 
.A(n_926),
.B(n_447),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_837),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_SL g1029 ( 
.A1(n_888),
.A2(n_398),
.B1(n_402),
.B2(n_392),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_932),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_883),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_831),
.A2(n_681),
.B(n_792),
.C(n_788),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_853),
.B(n_705),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_889),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_907),
.B(n_711),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_846),
.B(n_787),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_907),
.B(n_711),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_941),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_948),
.B(n_711),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_975),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_948),
.B(n_746),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_846),
.B(n_787),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_920),
.A2(n_826),
.B(n_820),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_855),
.B(n_746),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_916),
.B(n_746),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_944),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_884),
.B(n_757),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_920),
.A2(n_827),
.B(n_826),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_884),
.B(n_757),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_892),
.B(n_757),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_993),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_892),
.B(n_770),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_878),
.B(n_801),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_963),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_874),
.A2(n_827),
.B1(n_764),
.B2(n_784),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_842),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_916),
.B(n_770),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_894),
.B(n_770),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_975),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_999),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_847),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_848),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_861),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_867),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_895),
.B(n_897),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_939),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_912),
.B(n_787),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_969),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_877),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_891),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_979),
.B(n_784),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_922),
.A2(n_802),
.B(n_784),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_895),
.B(n_802),
.Y(n_1073)
);

NAND2x1_ASAP7_75t_L g1074 ( 
.A(n_906),
.B(n_764),
.Y(n_1074)
);

INVx5_ASAP7_75t_L g1075 ( 
.A(n_883),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_900),
.B(n_802),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_967),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_967),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_856),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_887),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_981),
.B(n_518),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_953),
.B(n_519),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_972),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_894),
.B(n_992),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_992),
.B(n_764),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_852),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_874),
.A2(n_957),
.B1(n_980),
.B2(n_968),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_981),
.B(n_522),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_917),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_849),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_830),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_972),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_990),
.A2(n_823),
.B1(n_768),
.B2(n_822),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_880),
.B(n_768),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_829),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_919),
.B(n_793),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_885),
.B(n_771),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_870),
.B(n_771),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_937),
.A2(n_772),
.B1(n_822),
.B2(n_777),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_865),
.B(n_793),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_957),
.A2(n_980),
.B1(n_968),
.B2(n_933),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_982),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_983),
.B(n_522),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_989),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_991),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_872),
.A2(n_410),
.B1(n_415),
.B2(n_405),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_913),
.B(n_935),
.C(n_952),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_998),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_952),
.B(n_933),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_873),
.B(n_772),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_866),
.A2(n_408),
.B1(n_414),
.B2(n_532),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_893),
.B(n_777),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_858),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_911),
.A2(n_904),
.B(n_843),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_845),
.B(n_871),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_909),
.A2(n_783),
.B1(n_818),
.B2(n_815),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_903),
.B(n_793),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_833),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_938),
.B(n_778),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_SL g1120 ( 
.A1(n_995),
.A2(n_538),
.B1(n_523),
.B2(n_527),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_982),
.A2(n_783),
.B1(n_818),
.B2(n_815),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_875),
.B(n_778),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_876),
.B(n_786),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_906),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_890),
.B(n_786),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_901),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_835),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_838),
.B(n_793),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_923),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_934),
.B(n_807),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_943),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_947),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_938),
.B(n_523),
.Y(n_1133)
);

OR2x2_ASAP7_75t_SL g1134 ( 
.A(n_973),
.B(n_529),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_937),
.A2(n_811),
.B1(n_807),
.B2(n_814),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_937),
.A2(n_811),
.B1(n_804),
.B2(n_828),
.Y(n_1136)
);

AND2x6_ASAP7_75t_SL g1137 ( 
.A(n_949),
.B(n_529),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_954),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_L g1139 ( 
.A(n_851),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_840),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_971),
.A2(n_804),
.B1(n_794),
.B2(n_797),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_862),
.A2(n_828),
.B(n_794),
.C(n_797),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_854),
.B(n_474),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_914),
.A2(n_804),
.B1(n_530),
.B2(n_532),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_914),
.A2(n_804),
.B1(n_530),
.B2(n_531),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_949),
.B(n_531),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_859),
.B(n_610),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_839),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_921),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_902),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_908),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_863),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_929),
.B(n_936),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_915),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_946),
.B(n_538),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_987),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_950),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_951),
.B(n_429),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_834),
.A2(n_587),
.B(n_575),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_869),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_959),
.A2(n_539),
.B1(n_540),
.B2(n_543),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_886),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_956),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_860),
.B(n_610),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_960),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_862),
.A2(n_435),
.B1(n_440),
.B2(n_441),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_961),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_905),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_994),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_988),
.B(n_539),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_959),
.A2(n_543),
.B1(n_401),
.B2(n_403),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_905),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_996),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_860),
.B(n_474),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_925),
.A2(n_437),
.B1(n_440),
.B2(n_441),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_942),
.A2(n_618),
.B(n_610),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_832),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_967),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_984),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_834),
.B(n_821),
.Y(n_1180)
);

OR2x2_ASAP7_75t_SL g1181 ( 
.A(n_930),
.B(n_395),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_930),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_832),
.B(n_610),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_832),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_997),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_967),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_881),
.B(n_431),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_997),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_940),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1065),
.A2(n_850),
.B(n_843),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1061),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1065),
.A2(n_868),
.B(n_850),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1109),
.A2(n_985),
.B1(n_974),
.B2(n_970),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1034),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1017),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1044),
.A2(n_868),
.B(n_881),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_L g1197 ( 
.A(n_1059),
.B(n_832),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1044),
.A2(n_898),
.B(n_910),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1086),
.Y(n_1199)
);

OR2x6_ASAP7_75t_L g1200 ( 
.A(n_1004),
.B(n_940),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1133),
.B(n_1146),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1101),
.A2(n_898),
.B1(n_974),
.B2(n_970),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1087),
.A2(n_985),
.B1(n_962),
.B2(n_958),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1090),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1021),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1094),
.A2(n_955),
.B(n_945),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1062),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1169),
.A2(n_945),
.B1(n_962),
.B2(n_958),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1102),
.B(n_955),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1013),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1094),
.A2(n_896),
.B(n_832),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1153),
.A2(n_424),
.B(n_430),
.C(n_448),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1079),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1111),
.A2(n_439),
.B(n_592),
.C(n_585),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1021),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1140),
.B(n_431),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1000),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_L g1218 ( 
.A1(n_1187),
.A2(n_597),
.B(n_585),
.C(n_592),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1028),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1075),
.Y(n_1220)
);

INVx3_ASAP7_75t_SL g1221 ( 
.A(n_1104),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1019),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1022),
.A2(n_434),
.B1(n_435),
.B2(n_437),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1097),
.A2(n_896),
.B(n_832),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1066),
.A2(n_1064),
.B1(n_1063),
.B2(n_1038),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1120),
.B(n_896),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1075),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1083),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1008),
.A2(n_1001),
.B1(n_1020),
.B2(n_1084),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1167),
.A2(n_597),
.B(n_585),
.C(n_592),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1132),
.Y(n_1231)
);

BUFx4f_ASAP7_75t_SL g1232 ( 
.A(n_1016),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_1056),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1155),
.B(n_434),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1114),
.A2(n_575),
.B(n_594),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1157),
.B(n_443),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1030),
.A2(n_1),
.B(n_2),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1046),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1075),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1001),
.B(n_896),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1097),
.A2(n_931),
.B(n_896),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1082),
.B(n_4),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1165),
.B(n_443),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1163),
.B(n_445),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1054),
.Y(n_1245)
);

OAI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1081),
.A2(n_445),
.B1(n_351),
.B2(n_344),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1081),
.B(n_896),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1031),
.B(n_1075),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1088),
.B(n_931),
.Y(n_1249)
);

OR2x6_ASAP7_75t_SL g1250 ( 
.A(n_1171),
.B(n_270),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1137),
.B(n_273),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1069),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1107),
.A2(n_585),
.B(n_597),
.C(n_592),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1105),
.A2(n_597),
.B1(n_370),
.B2(n_361),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1080),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1112),
.A2(n_931),
.B(n_673),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1088),
.B(n_931),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1045),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1114),
.A2(n_618),
.B(n_610),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1170),
.B(n_931),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1051),
.Y(n_1261)
);

NAND2x2_ASAP7_75t_L g1262 ( 
.A(n_1091),
.B(n_4),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1003),
.Y(n_1263)
);

INVx3_ASAP7_75t_SL g1264 ( 
.A(n_1083),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1139),
.B(n_931),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1179),
.B(n_275),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1139),
.B(n_673),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1173),
.B(n_276),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1031),
.B(n_673),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1060),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1112),
.A2(n_1049),
.B(n_1047),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1108),
.A2(n_338),
.B1(n_331),
.B2(n_330),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1150),
.B(n_610),
.Y(n_1273)
);

INVx5_ASAP7_75t_L g1274 ( 
.A(n_1013),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1013),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1149),
.B(n_808),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1119),
.A2(n_600),
.B(n_587),
.C(n_589),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1002),
.A2(n_309),
.B1(n_308),
.B2(n_307),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1011),
.A2(n_323),
.B1(n_305),
.B2(n_303),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1068),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1053),
.B(n_280),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1151),
.B(n_808),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1045),
.B(n_673),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1011),
.A2(n_767),
.B1(n_967),
.B2(n_808),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1089),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1047),
.A2(n_618),
.B(n_808),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1106),
.A2(n_605),
.B(n_600),
.C(n_595),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1181),
.B(n_284),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1083),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1057),
.B(n_673),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1143),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1057),
.B(n_751),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1154),
.B(n_821),
.Y(n_1293)
);

AOI33xp33_ASAP7_75t_L g1294 ( 
.A1(n_1175),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.B3(n_12),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_L g1295 ( 
.A1(n_1100),
.A2(n_589),
.B(n_594),
.C(n_595),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1070),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1007),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1003),
.B(n_808),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1113),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1106),
.A2(n_605),
.B(n_600),
.C(n_595),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1002),
.B(n_808),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1059),
.B(n_1039),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1160),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1166),
.B(n_413),
.C(n_288),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1177),
.A2(n_605),
.B(n_589),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1103),
.B(n_5),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1059),
.B(n_821),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1103),
.B(n_1143),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1126),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1115),
.B(n_10),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_SL g1311 ( 
.A(n_1059),
.B(n_751),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1156),
.B(n_1115),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1158),
.A2(n_594),
.B(n_13),
.C(n_14),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1006),
.B(n_618),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1127),
.B(n_287),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_R g1316 ( 
.A(n_1092),
.B(n_767),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1032),
.A2(n_293),
.B(n_296),
.C(n_343),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1049),
.A2(n_821),
.B(n_751),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1129),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1131),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1138),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1148),
.B(n_372),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1152),
.B(n_618),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1143),
.B(n_419),
.Y(n_1325)
);

INVx4_ASAP7_75t_SL g1326 ( 
.A(n_1005),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1161),
.B(n_12),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1134),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1076),
.A2(n_1145),
.B1(n_1144),
.B2(n_1162),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1122),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1050),
.A2(n_821),
.B(n_751),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1039),
.B(n_751),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1092),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1050),
.A2(n_754),
.B(n_377),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1041),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1174),
.B(n_13),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1110),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1110),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1041),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1023),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1076),
.A2(n_1033),
.B1(n_1035),
.B2(n_1037),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1023),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1005),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1024),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1025),
.A2(n_20),
.B(n_21),
.C(n_27),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1124),
.B(n_383),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1012),
.B(n_20),
.Y(n_1347)
);

CKINVDCx16_ASAP7_75t_R g1348 ( 
.A(n_1029),
.Y(n_1348)
);

BUFx2_ASAP7_75t_SL g1349 ( 
.A(n_1092),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1171),
.B(n_754),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1095),
.B(n_754),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1033),
.B(n_618),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1326),
.B(n_1036),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1232),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1250),
.B(n_1095),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1305),
.A2(n_1159),
.B(n_1184),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1234),
.A2(n_1024),
.B(n_1037),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_SL g1358 ( 
.A1(n_1317),
.A2(n_1074),
.B(n_1067),
.C(n_1096),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1201),
.B(n_1168),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1211),
.A2(n_1184),
.B(n_1072),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1212),
.A2(n_1209),
.B(n_1208),
.C(n_1202),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1224),
.A2(n_1072),
.B(n_1048),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1241),
.A2(n_1048),
.B(n_1043),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1229),
.A2(n_1035),
.B1(n_1026),
.B2(n_1182),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1242),
.B(n_1172),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1217),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1271),
.A2(n_1052),
.B(n_1073),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1222),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1312),
.B(n_1337),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1312),
.B(n_1189),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1335),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1303),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1338),
.B(n_1124),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1193),
.A2(n_1142),
.B1(n_1136),
.B2(n_1073),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1247),
.B(n_1095),
.Y(n_1375)
);

NAND2x1_ASAP7_75t_L g1376 ( 
.A(n_1343),
.B(n_1009),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1341),
.A2(n_1052),
.B(n_1117),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1219),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1202),
.A2(n_1042),
.B(n_1185),
.C(n_1015),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1238),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1348),
.B(n_1308),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1225),
.B(n_1058),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1259),
.A2(n_1043),
.B(n_1176),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1225),
.B(n_1085),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1325),
.A2(n_1010),
.B1(n_1093),
.B2(n_1135),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1219),
.B(n_1118),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1325),
.A2(n_1099),
.B1(n_1032),
.B2(n_1055),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1190),
.A2(n_1121),
.B(n_1098),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1260),
.A2(n_1018),
.B(n_1183),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1328),
.B(n_1118),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1296),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1245),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1203),
.B(n_1294),
.C(n_1281),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1341),
.A2(n_1183),
.B(n_1040),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1279),
.A2(n_1005),
.B1(n_1118),
.B2(n_1071),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1220),
.Y(n_1396)
);

AO32x2_ASAP7_75t_L g1397 ( 
.A1(n_1203),
.A2(n_1027),
.A3(n_1071),
.B1(n_1128),
.B2(n_1123),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1206),
.A2(n_1122),
.A3(n_1123),
.B(n_1125),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1345),
.A2(n_1147),
.B1(n_1130),
.B2(n_1125),
.C(n_1164),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1192),
.A2(n_1176),
.B(n_1116),
.Y(n_1400)
);

BUFx10_ASAP7_75t_L g1401 ( 
.A(n_1194),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1199),
.B(n_21),
.Y(n_1402)
);

OAI22x1_ASAP7_75t_L g1403 ( 
.A1(n_1288),
.A2(n_1186),
.B1(n_1130),
.B2(n_1180),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1280),
.Y(n_1404)
);

INVxp67_ASAP7_75t_SL g1405 ( 
.A(n_1233),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1259),
.A2(n_1147),
.B(n_1014),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1313),
.A2(n_1141),
.B(n_1180),
.C(n_1009),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1258),
.B(n_1339),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1196),
.A2(n_1240),
.B(n_1198),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1277),
.A2(n_1164),
.B(n_391),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1220),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1249),
.B(n_1014),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1197),
.A2(n_1040),
.B(n_1078),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1256),
.A2(n_1078),
.B(n_1077),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1324),
.A2(n_1005),
.B(n_1078),
.Y(n_1415)
);

BUFx5_ASAP7_75t_L g1416 ( 
.A(n_1340),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1342),
.B(n_1178),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1257),
.B(n_1078),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1324),
.A2(n_1077),
.B(n_425),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1339),
.B(n_36),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1236),
.B(n_36),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1205),
.Y(n_1422)
);

NOR2xp67_ASAP7_75t_L g1423 ( 
.A(n_1289),
.B(n_1077),
.Y(n_1423)
);

O2A1O1Ixp5_ASAP7_75t_SL g1424 ( 
.A1(n_1319),
.A2(n_1299),
.B(n_1321),
.C(n_1320),
.Y(n_1424)
);

AO21x1_ASAP7_75t_L g1425 ( 
.A1(n_1329),
.A2(n_425),
.B(n_767),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1266),
.B(n_1336),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1291),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1227),
.B(n_1239),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1251),
.B(n_38),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1191),
.Y(n_1430)
);

NAND2x1p5_ASAP7_75t_L g1431 ( 
.A(n_1210),
.B(n_754),
.Y(n_1431)
);

AO32x2_ASAP7_75t_L g1432 ( 
.A1(n_1329),
.A2(n_767),
.A3(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1252),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1221),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1350),
.A2(n_754),
.B(n_419),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1295),
.A2(n_425),
.B(n_767),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1350),
.A2(n_419),
.B(n_433),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1344),
.A2(n_419),
.B(n_433),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1214),
.A2(n_1310),
.B(n_1327),
.C(n_1304),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_L g1440 ( 
.A(n_1228),
.B(n_155),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1352),
.A2(n_419),
.B(n_433),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1253),
.A2(n_425),
.B(n_767),
.Y(n_1442)
);

AO31x2_ASAP7_75t_L g1443 ( 
.A1(n_1330),
.A2(n_618),
.A3(n_433),
.B(n_615),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1255),
.B(n_1285),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1200),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1226),
.A2(n_449),
.B(n_406),
.C(n_407),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1352),
.A2(n_433),
.B(n_393),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1230),
.A2(n_38),
.B(n_39),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1334),
.A2(n_1265),
.B(n_1286),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1286),
.A2(n_411),
.B(n_619),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1314),
.A2(n_619),
.B(n_615),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1227),
.B(n_619),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1272),
.A2(n_40),
.B(n_42),
.C(n_45),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1207),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1268),
.B(n_47),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1314),
.A2(n_619),
.B(n_615),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1326),
.B(n_145),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1287),
.A2(n_619),
.B(n_615),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1315),
.B(n_47),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1267),
.A2(n_50),
.B(n_51),
.C(n_54),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1227),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1239),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1300),
.A2(n_609),
.B(n_604),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1301),
.A2(n_609),
.A3(n_604),
.B(n_601),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1216),
.B(n_1323),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1243),
.B(n_50),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1309),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1218),
.A2(n_609),
.B(n_604),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_609),
.B(n_604),
.Y(n_1469)
);

AND2x6_ASAP7_75t_SL g1470 ( 
.A(n_1200),
.B(n_54),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1322),
.B(n_56),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1331),
.A2(n_609),
.B(n_604),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_SL g1473 ( 
.A1(n_1306),
.A2(n_57),
.B(n_59),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1311),
.A2(n_604),
.B(n_601),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1311),
.A2(n_601),
.B(n_152),
.Y(n_1475)
);

BUFx8_ASAP7_75t_L g1476 ( 
.A(n_1215),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1264),
.Y(n_1477)
);

AO22x1_ASAP7_75t_L g1478 ( 
.A1(n_1333),
.A2(n_1263),
.B1(n_1248),
.B2(n_1346),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1223),
.B(n_1244),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1343),
.A2(n_601),
.B(n_148),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1239),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1273),
.A2(n_601),
.B(n_157),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1200),
.B(n_59),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1213),
.B(n_60),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1231),
.B(n_60),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1261),
.B(n_63),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1325),
.A2(n_601),
.B(n_159),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1270),
.B(n_63),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1282),
.A2(n_163),
.B(n_221),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1273),
.A2(n_134),
.B(n_218),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1349),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1293),
.A2(n_133),
.B(n_212),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1276),
.A2(n_129),
.B(n_202),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1297),
.B(n_65),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1272),
.B(n_65),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1326),
.B(n_225),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1351),
.A2(n_120),
.B(n_196),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1284),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1248),
.B(n_70),
.Y(n_1499)
);

AO32x2_ASAP7_75t_L g1500 ( 
.A1(n_1254),
.A2(n_1278),
.A3(n_1237),
.B1(n_1262),
.B2(n_1347),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1292),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1302),
.B(n_71),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1298),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1246),
.B(n_87),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1302),
.A2(n_99),
.B(n_101),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1278),
.A2(n_104),
.B(n_105),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1307),
.A2(n_168),
.B(n_173),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1210),
.B(n_200),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1332),
.A2(n_177),
.B(n_183),
.Y(n_1509)
);

AOI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1254),
.A2(n_190),
.B(n_192),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1275),
.B(n_1292),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1283),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1210),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1210),
.A2(n_1274),
.B(n_1269),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1274),
.A2(n_1275),
.B(n_1316),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1274),
.A2(n_1275),
.B(n_1195),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1204),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1274),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1220),
.Y(n_1519)
);

AO31x2_ASAP7_75t_L g1520 ( 
.A1(n_1341),
.A2(n_1271),
.A3(n_1206),
.B(n_1203),
.Y(n_1520)
);

OAI21xp33_ASAP7_75t_L g1521 ( 
.A1(n_1201),
.A2(n_678),
.B(n_1109),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1235),
.A2(n_1305),
.B(n_1224),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1201),
.B(n_1086),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1199),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1271),
.A2(n_1109),
.B(n_1190),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1260),
.A2(n_1341),
.B(n_1271),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1201),
.A2(n_1109),
.B1(n_678),
.B2(n_1169),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1235),
.A2(n_1305),
.B(n_1224),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_SL g1529 ( 
.A1(n_1382),
.A2(n_1384),
.B(n_1448),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1525),
.A2(n_1362),
.B(n_1526),
.Y(n_1530)
);

OAI222xp33_ASAP7_75t_L g1531 ( 
.A1(n_1527),
.A2(n_1364),
.B1(n_1385),
.B2(n_1426),
.C1(n_1495),
.C2(n_1498),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1444),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1366),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1477),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1361),
.A2(n_1521),
.B(n_1393),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1393),
.A2(n_1521),
.B(n_1453),
.C(n_1439),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1476),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1514),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1528),
.A2(n_1363),
.B(n_1360),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1364),
.A2(n_1385),
.B1(n_1387),
.B2(n_1498),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1378),
.B(n_1523),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1515),
.B(n_1503),
.Y(n_1542)
);

OAI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1502),
.A2(n_1421),
.B1(n_1455),
.B2(n_1479),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1458),
.A2(n_1419),
.B(n_1356),
.Y(n_1544)
);

CKINVDCx14_ASAP7_75t_R g1545 ( 
.A(n_1422),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1459),
.A2(n_1429),
.B1(n_1483),
.B2(n_1387),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1354),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1430),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1437),
.A2(n_1379),
.B(n_1374),
.C(n_1506),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1504),
.A2(n_1466),
.B1(n_1365),
.B2(n_1374),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1454),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1369),
.B(n_1370),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1427),
.B(n_1368),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1367),
.A2(n_1383),
.B(n_1449),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1369),
.B(n_1370),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1434),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1415),
.A2(n_1441),
.B(n_1482),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1401),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1380),
.Y(n_1560)
);

AO31x2_ASAP7_75t_L g1561 ( 
.A1(n_1425),
.A2(n_1403),
.A3(n_1438),
.B(n_1447),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1525),
.A2(n_1388),
.B(n_1400),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1514),
.B(n_1353),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1435),
.A2(n_1388),
.B(n_1400),
.C(n_1496),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1503),
.B(n_1518),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1394),
.A2(n_1414),
.B(n_1480),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_R g1567 ( 
.A(n_1513),
.B(n_1381),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1399),
.A2(n_1463),
.B(n_1468),
.Y(n_1568)
);

AOI22x1_ASAP7_75t_L g1569 ( 
.A1(n_1372),
.A2(n_1473),
.B1(n_1405),
.B2(n_1391),
.Y(n_1569)
);

BUFx4f_ASAP7_75t_L g1570 ( 
.A(n_1457),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1371),
.B(n_1359),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1389),
.A2(n_1456),
.B(n_1451),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1353),
.B(n_1516),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1451),
.A2(n_1456),
.B(n_1357),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1399),
.A2(n_1463),
.B(n_1468),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1377),
.A2(n_1406),
.B(n_1490),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1442),
.A2(n_1436),
.B(n_1450),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1392),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1493),
.A2(n_1474),
.B(n_1510),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1402),
.B(n_1390),
.Y(n_1580)
);

BUFx4f_ASAP7_75t_SL g1581 ( 
.A(n_1401),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1467),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1416),
.B(n_1433),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1410),
.A2(n_1507),
.B(n_1413),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1410),
.A2(n_1505),
.B(n_1489),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1489),
.A2(n_1475),
.B(n_1492),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1478),
.Y(n_1587)
);

A2O1A1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1457),
.A2(n_1496),
.B(n_1471),
.C(n_1407),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1373),
.A2(n_1424),
.B(n_1497),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1471),
.A2(n_1373),
.B(n_1508),
.C(n_1417),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1502),
.A2(n_1355),
.B1(n_1445),
.B2(n_1524),
.Y(n_1591)
);

AOI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1418),
.A2(n_1375),
.B(n_1452),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1386),
.B(n_1502),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1408),
.B(n_1511),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1358),
.A2(n_1409),
.B(n_1417),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1446),
.A2(n_1420),
.B(n_1509),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1491),
.B(n_1500),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1487),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1520),
.A2(n_1376),
.B(n_1508),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1470),
.B(n_1499),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1470),
.A2(n_1488),
.B1(n_1484),
.B2(n_1485),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1517),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1486),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1494),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1512),
.A2(n_1395),
.B(n_1520),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1432),
.A2(n_1500),
.B(n_1440),
.C(n_1520),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1411),
.Y(n_1607)
);

AO21x2_ASAP7_75t_L g1608 ( 
.A1(n_1428),
.A2(n_1423),
.B(n_1464),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1396),
.B(n_1481),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1411),
.Y(n_1610)
);

AOI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1432),
.A2(n_1519),
.B(n_1462),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1431),
.A2(n_1464),
.B(n_1398),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1431),
.A2(n_1464),
.B(n_1416),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1461),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1461),
.A2(n_1462),
.B1(n_1519),
.B2(n_1397),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1460),
.A2(n_1432),
.B1(n_1397),
.B2(n_1519),
.C(n_1416),
.Y(n_1616)
);

NAND2x1_ASAP7_75t_L g1617 ( 
.A(n_1443),
.B(n_1384),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1443),
.A2(n_613),
.B1(n_1393),
.B2(n_1201),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1443),
.A2(n_1472),
.B(n_1469),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1501),
.B(n_1514),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1444),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1444),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1525),
.A2(n_1362),
.B(n_1526),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1527),
.B(n_1402),
.Y(n_1624)
);

AO31x2_ASAP7_75t_L g1625 ( 
.A1(n_1425),
.A2(n_1341),
.A3(n_1526),
.B(n_1271),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1361),
.A2(n_1521),
.B(n_1109),
.C(n_678),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1444),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1527),
.B(n_1109),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1371),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_SL g1630 ( 
.A1(n_1361),
.A2(n_1382),
.B(n_1393),
.C(n_1109),
.Y(n_1630)
);

NAND2x1_ASAP7_75t_L g1631 ( 
.A(n_1384),
.B(n_1382),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_SL g1633 ( 
.A1(n_1382),
.A2(n_1384),
.B(n_1448),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1520),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1444),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1469),
.A2(n_1472),
.B(n_1522),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1444),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1469),
.A2(n_1472),
.B(n_1522),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1477),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1393),
.A2(n_1109),
.B1(n_1201),
.B2(n_1521),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1444),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1469),
.A2(n_1472),
.B(n_1522),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1527),
.A2(n_1109),
.B1(n_678),
.B2(n_1101),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1393),
.A2(n_1109),
.B1(n_1201),
.B2(n_1521),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1527),
.A2(n_1348),
.B1(n_1001),
.B2(n_1008),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1527),
.A2(n_1109),
.B(n_678),
.Y(n_1646)
);

NOR3xp33_ASAP7_75t_L g1647 ( 
.A(n_1393),
.B(n_1109),
.C(n_1361),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1527),
.B(n_1402),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1527),
.B(n_1402),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1477),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1444),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1444),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1444),
.Y(n_1654)
);

AND2x2_ASAP7_75t_SL g1655 ( 
.A(n_1382),
.B(n_1109),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1469),
.A2(n_1472),
.B(n_1522),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1477),
.Y(n_1657)
);

AO31x2_ASAP7_75t_L g1658 ( 
.A1(n_1425),
.A2(n_1341),
.A3(n_1526),
.B(n_1271),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1477),
.Y(n_1659)
);

AND2x4_ASAP7_75t_SL g1660 ( 
.A(n_1354),
.B(n_1401),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1444),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1527),
.B(n_1109),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1501),
.B(n_1514),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1444),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1393),
.A2(n_1109),
.B1(n_1201),
.B2(n_1521),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1393),
.A2(n_1109),
.B1(n_1201),
.B2(n_1521),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1444),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1371),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1501),
.B(n_1514),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1502),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1361),
.A2(n_1109),
.B(n_1393),
.C(n_1521),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1525),
.A2(n_1362),
.B(n_1526),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1477),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1361),
.A2(n_1109),
.B(n_1393),
.C(n_1521),
.Y(n_1674)
);

AO21x2_ASAP7_75t_L g1675 ( 
.A1(n_1526),
.A2(n_1367),
.B(n_1271),
.Y(n_1675)
);

AO22x1_ASAP7_75t_L g1676 ( 
.A1(n_1495),
.A2(n_1109),
.B1(n_582),
.B2(n_614),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1371),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1526),
.A2(n_1525),
.B(n_1382),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1469),
.A2(n_1472),
.B(n_1522),
.Y(n_1679)
);

AOI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1393),
.A2(n_1109),
.B(n_1361),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1527),
.B(n_1109),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1469),
.A2(n_1472),
.B(n_1522),
.Y(n_1682)
);

BUFx2_ASAP7_75t_R g1683 ( 
.A(n_1422),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1525),
.A2(n_1362),
.B(n_1526),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1372),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1404),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1525),
.A2(n_1362),
.B(n_1526),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1527),
.B(n_1109),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1527),
.A2(n_1109),
.B(n_678),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1371),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1361),
.B(n_1109),
.C(n_1393),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1393),
.A2(n_613),
.B1(n_1201),
.B2(n_966),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1476),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1527),
.A2(n_1109),
.B(n_678),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1527),
.A2(n_1101),
.B1(n_1393),
.B2(n_1250),
.Y(n_1695)
);

OAI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1527),
.A2(n_1101),
.B1(n_1393),
.B2(n_1250),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1477),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1526),
.A2(n_1525),
.B(n_1382),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1444),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1605),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1685),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1646),
.A2(n_1689),
.B(n_1694),
.C(n_1626),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1599),
.B(n_1563),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1626),
.A2(n_1662),
.B(n_1681),
.C(n_1628),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1678),
.A2(n_1698),
.B(n_1539),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1634),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1678),
.A2(n_1698),
.B(n_1606),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1634),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1649),
.B(n_1650),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1532),
.B(n_1621),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1541),
.B(n_1554),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1622),
.B(n_1627),
.Y(n_1714)
);

NOR2xp67_ASAP7_75t_L g1715 ( 
.A(n_1559),
.B(n_1670),
.Y(n_1715)
);

NAND2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1631),
.B(n_1547),
.Y(n_1716)
);

INVxp33_ASAP7_75t_L g1717 ( 
.A(n_1549),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1588),
.A2(n_1674),
.B(n_1671),
.Y(n_1718)
);

OA21x2_ASAP7_75t_L g1719 ( 
.A1(n_1606),
.A2(n_1555),
.B(n_1595),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1693),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1670),
.B(n_1573),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1645),
.A2(n_1681),
.B1(n_1662),
.B2(n_1628),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1723)
);

AND2x4_ASAP7_75t_SL g1724 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1641),
.B(n_1652),
.Y(n_1725)
);

CKINVDCx16_ASAP7_75t_R g1726 ( 
.A(n_1602),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1605),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1588),
.A2(n_1674),
.B(n_1671),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1653),
.B(n_1654),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1570),
.B(n_1587),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1688),
.A2(n_1692),
.B1(n_1643),
.B2(n_1546),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1536),
.A2(n_1590),
.B(n_1564),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1538),
.B(n_1620),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1661),
.B(n_1664),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1540),
.A2(n_1691),
.B(n_1688),
.C(n_1647),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1663),
.B(n_1669),
.Y(n_1736)
);

AND2x6_ASAP7_75t_L g1737 ( 
.A(n_1663),
.B(n_1669),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1583),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1667),
.B(n_1699),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1571),
.B(n_1597),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1533),
.Y(n_1741)
);

O2A1O1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1695),
.A2(n_1696),
.B(n_1680),
.C(n_1647),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1582),
.B(n_1629),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1571),
.B(n_1668),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1677),
.B(n_1690),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1695),
.A2(n_1696),
.B(n_1680),
.C(n_1630),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1550),
.A2(n_1648),
.B(n_1632),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1560),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1578),
.B(n_1610),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1593),
.B(n_1546),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1686),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1540),
.A2(n_1692),
.B1(n_1666),
.B2(n_1644),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1553),
.B(n_1556),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1535),
.A2(n_1616),
.B(n_1611),
.C(n_1666),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1594),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1548),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1552),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1600),
.B(n_1551),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1551),
.B(n_1614),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1640),
.A2(n_1644),
.B1(n_1665),
.B2(n_1543),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1632),
.B(n_1648),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1640),
.A2(n_1665),
.B1(n_1543),
.B2(n_1601),
.Y(n_1765)
);

O2A1O1Ixp5_ASAP7_75t_L g1766 ( 
.A1(n_1531),
.A2(n_1595),
.B(n_1599),
.C(n_1598),
.Y(n_1766)
);

O2A1O1Ixp5_ASAP7_75t_L g1767 ( 
.A1(n_1531),
.A2(n_1598),
.B(n_1601),
.C(n_1596),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1553),
.B(n_1556),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1534),
.B(n_1639),
.Y(n_1769)
);

O2A1O1Ixp33_ASAP7_75t_L g1770 ( 
.A1(n_1529),
.A2(n_1633),
.B(n_1590),
.C(n_1562),
.Y(n_1770)
);

INVx3_ASAP7_75t_SL g1771 ( 
.A(n_1537),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1618),
.A2(n_1562),
.B1(n_1569),
.B2(n_1616),
.Y(n_1772)
);

O2A1O1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1611),
.A2(n_1603),
.B(n_1604),
.C(n_1615),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_L g1774 ( 
.A(n_1676),
.B(n_1618),
.C(n_1589),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1581),
.A2(n_1607),
.B1(n_1534),
.B2(n_1697),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1609),
.B(n_1639),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1530),
.Y(n_1777)
);

O2A1O1Ixp5_ASAP7_75t_L g1778 ( 
.A1(n_1617),
.A2(n_1592),
.B(n_1658),
.C(n_1625),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1542),
.A2(n_1608),
.B(n_1568),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1639),
.B(n_1651),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1530),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1651),
.B(n_1673),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1581),
.A2(n_1673),
.B1(n_1697),
.B2(n_1651),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1657),
.B(n_1697),
.Y(n_1784)
);

AOI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1567),
.A2(n_1673),
.B(n_1657),
.C(n_1586),
.Y(n_1785)
);

O2A1O1Ixp5_ASAP7_75t_L g1786 ( 
.A1(n_1625),
.A2(n_1658),
.B(n_1575),
.C(n_1568),
.Y(n_1786)
);

AOI21x1_ASAP7_75t_SL g1787 ( 
.A1(n_1675),
.A2(n_1687),
.B(n_1684),
.Y(n_1787)
);

AOI21x1_ASAP7_75t_SL g1788 ( 
.A1(n_1675),
.A2(n_1687),
.B(n_1684),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1623),
.A2(n_1672),
.B(n_1579),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1660),
.B(n_1613),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1545),
.B(n_1683),
.Y(n_1791)
);

OA21x2_ASAP7_75t_L g1792 ( 
.A1(n_1585),
.A2(n_1612),
.B(n_1576),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1575),
.A2(n_1672),
.B(n_1623),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1577),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1561),
.B(n_1574),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1572),
.A2(n_1584),
.B(n_1566),
.C(n_1558),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1561),
.Y(n_1797)
);

AOI21x1_ASAP7_75t_SL g1798 ( 
.A1(n_1544),
.A2(n_1656),
.B(n_1682),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1577),
.B(n_1619),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1636),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1638),
.B(n_1642),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1679),
.A2(n_1643),
.B1(n_1662),
.B2(n_1628),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1634),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1646),
.A2(n_1689),
.B(n_1694),
.C(n_1626),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1634),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1643),
.A2(n_1662),
.B1(n_1681),
.B2(n_1628),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1565),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1626),
.A2(n_1588),
.B(n_1109),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1659),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1570),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1541),
.B(n_1554),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1646),
.A2(n_1689),
.B(n_1694),
.C(n_1626),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1646),
.A2(n_1689),
.B(n_1694),
.C(n_1626),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1643),
.A2(n_1662),
.B1(n_1681),
.B2(n_1628),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1659),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1659),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1824)
);

OA21x2_ASAP7_75t_L g1825 ( 
.A1(n_1678),
.A2(n_1698),
.B(n_1539),
.Y(n_1825)
);

A2O1A1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1626),
.A2(n_1109),
.B(n_1643),
.C(n_1540),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1643),
.A2(n_1662),
.B1(n_1681),
.B2(n_1628),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1626),
.A2(n_1588),
.B(n_1109),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1643),
.A2(n_1662),
.B1(n_1681),
.B2(n_1628),
.Y(n_1830)
);

INVx3_ASAP7_75t_SL g1831 ( 
.A(n_1537),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1629),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1580),
.B(n_1624),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_L g1835 ( 
.A1(n_1695),
.A2(n_1696),
.B(n_1543),
.C(n_1645),
.Y(n_1835)
);

OA21x2_ASAP7_75t_L g1836 ( 
.A1(n_1678),
.A2(n_1698),
.B(n_1539),
.Y(n_1836)
);

O2A1O1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1646),
.A2(n_1689),
.B(n_1694),
.C(n_1626),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1685),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1646),
.A2(n_1689),
.B(n_1694),
.C(n_1626),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1626),
.A2(n_1588),
.B(n_1109),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1655),
.B(n_1549),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1749),
.Y(n_1843)
);

AO21x2_ASAP7_75t_L g1844 ( 
.A1(n_1789),
.A2(n_1774),
.B(n_1754),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1712),
.B(n_1812),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1738),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1708),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1741),
.Y(n_1848)
);

AO21x2_ASAP7_75t_L g1849 ( 
.A1(n_1774),
.A2(n_1754),
.B(n_1793),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1704),
.B(n_1732),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1738),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1748),
.Y(n_1852)
);

OA21x2_ASAP7_75t_L g1853 ( 
.A1(n_1786),
.A2(n_1766),
.B(n_1778),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1743),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1763),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1740),
.B(n_1708),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1794),
.Y(n_1857)
);

CKINVDCx20_ASAP7_75t_R g1858 ( 
.A(n_1726),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1707),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1753),
.B(n_1768),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1713),
.B(n_1813),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1800),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1814),
.B(n_1817),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1787),
.A2(n_1788),
.B(n_1798),
.Y(n_1864)
);

AO21x2_ASAP7_75t_L g1865 ( 
.A1(n_1797),
.A2(n_1772),
.B(n_1796),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1819),
.B(n_1838),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1709),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1803),
.B(n_1805),
.Y(n_1868)
);

OA21x2_ASAP7_75t_L g1869 ( 
.A1(n_1786),
.A2(n_1766),
.B(n_1778),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1703),
.B(n_1807),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1815),
.B(n_1822),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1704),
.B(n_1790),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1722),
.B(n_1806),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1799),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1704),
.B(n_1721),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1718),
.B(n_1728),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1842),
.B(n_1820),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1710),
.B(n_1824),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1777),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1781),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1751),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1757),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1827),
.B(n_1832),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1781),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1833),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1834),
.B(n_1744),
.Y(n_1886)
);

OA21x2_ASAP7_75t_L g1887 ( 
.A1(n_1700),
.A2(n_1727),
.B(n_1767),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1752),
.A2(n_1731),
.B1(n_1759),
.B2(n_1765),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1750),
.B(n_1755),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1758),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1714),
.Y(n_1891)
);

OA21x2_ASAP7_75t_L g1892 ( 
.A1(n_1727),
.A2(n_1767),
.B(n_1747),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1711),
.B(n_1729),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1745),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1723),
.Y(n_1895)
);

OA21x2_ASAP7_75t_L g1896 ( 
.A1(n_1747),
.A2(n_1795),
.B(n_1826),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1734),
.B(n_1739),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1792),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1792),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1828),
.B(n_1830),
.Y(n_1900)
);

AOI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1801),
.A2(n_1802),
.B(n_1761),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1719),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1725),
.Y(n_1903)
);

OAI21xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1809),
.A2(n_1841),
.B(n_1829),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1773),
.Y(n_1905)
);

AO21x2_ASAP7_75t_L g1906 ( 
.A1(n_1779),
.A2(n_1773),
.B(n_1826),
.Y(n_1906)
);

AO21x2_ASAP7_75t_L g1907 ( 
.A1(n_1742),
.A2(n_1746),
.B(n_1735),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1770),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1706),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1735),
.A2(n_1742),
.B(n_1705),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1770),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1733),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1736),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1756),
.Y(n_1914)
);

AO21x2_ASAP7_75t_L g1915 ( 
.A1(n_1746),
.A2(n_1762),
.B(n_1764),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1760),
.B(n_1776),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1737),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1717),
.B(n_1701),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1825),
.B(n_1836),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1825),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1839),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1859),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1859),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1856),
.B(n_1836),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1902),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1860),
.B(n_1782),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1877),
.B(n_1855),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1862),
.Y(n_1928)
);

INVxp67_ASAP7_75t_SL g1929 ( 
.A(n_1846),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1851),
.B(n_1705),
.Y(n_1930)
);

OAI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1864),
.A2(n_1787),
.B(n_1788),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1868),
.Y(n_1932)
);

OAI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1910),
.A2(n_1835),
.B(n_1840),
.C(n_1702),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1868),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1857),
.B(n_1785),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1867),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1857),
.B(n_1808),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_1889),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1872),
.B(n_1715),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1879),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1893),
.B(n_1897),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1893),
.B(n_1808),
.Y(n_1942)
);

INVx5_ASAP7_75t_L g1943 ( 
.A(n_1876),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1907),
.A2(n_1888),
.B1(n_1876),
.B2(n_1873),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1897),
.B(n_1724),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1860),
.B(n_1784),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1889),
.B(n_1702),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1874),
.B(n_1769),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1870),
.B(n_1780),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1848),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1870),
.B(n_1821),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1907),
.A2(n_1737),
.B1(n_1716),
.B2(n_1811),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1872),
.B(n_1737),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1852),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1854),
.B(n_1823),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1876),
.A2(n_1904),
.B1(n_1849),
.B2(n_1844),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1861),
.B(n_1863),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1878),
.B(n_1810),
.Y(n_1958)
);

INVx4_ASAP7_75t_L g1959 ( 
.A(n_1876),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1866),
.B(n_1840),
.Y(n_1960)
);

OAI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1956),
.A2(n_1904),
.B1(n_1905),
.B2(n_1901),
.C(n_1908),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1955),
.Y(n_1962)
);

OAI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1956),
.A2(n_1850),
.B1(n_1901),
.B2(n_1896),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1941),
.B(n_1894),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1950),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1933),
.A2(n_1906),
.B1(n_1844),
.B2(n_1915),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1944),
.A2(n_1906),
.B1(n_1905),
.B2(n_1896),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_R g1968 ( 
.A(n_1930),
.B(n_1858),
.Y(n_1968)
);

OAI222xp33_ASAP7_75t_L g1969 ( 
.A1(n_1947),
.A2(n_1850),
.B1(n_1908),
.B2(n_1911),
.C1(n_1845),
.C2(n_1883),
.Y(n_1969)
);

AND4x1_ASAP7_75t_L g1970 ( 
.A(n_1952),
.B(n_1791),
.C(n_1804),
.D(n_1816),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1935),
.A2(n_1906),
.B1(n_1850),
.B2(n_1911),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1960),
.A2(n_1804),
.B1(n_1816),
.B2(n_1818),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1927),
.B(n_1871),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1929),
.B(n_1938),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1949),
.B(n_1886),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1949),
.B(n_1886),
.Y(n_1976)
);

OAI211xp5_ASAP7_75t_L g1977 ( 
.A1(n_1924),
.A2(n_1818),
.B(n_1837),
.C(n_1896),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1959),
.A2(n_1837),
.B1(n_1892),
.B2(n_1843),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1926),
.B(n_1891),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1959),
.A2(n_1892),
.B1(n_1730),
.B2(n_1885),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1932),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_R g1982 ( 
.A(n_1943),
.B(n_1720),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1934),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1954),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1953),
.B(n_1875),
.Y(n_1985)
);

AO21x2_ASAP7_75t_L g1986 ( 
.A1(n_1931),
.A2(n_1898),
.B(n_1899),
.Y(n_1986)
);

AOI221xp5_ASAP7_75t_L g1987 ( 
.A1(n_1957),
.A2(n_1914),
.B1(n_1903),
.B2(n_1895),
.C(n_1891),
.Y(n_1987)
);

INVx1_ASAP7_75t_SL g1988 ( 
.A(n_1958),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1937),
.Y(n_1989)
);

NAND3xp33_ASAP7_75t_L g1990 ( 
.A(n_1936),
.B(n_1887),
.C(n_1869),
.Y(n_1990)
);

INVxp67_ASAP7_75t_SL g1991 ( 
.A(n_1940),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1951),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1953),
.B(n_1875),
.Y(n_1993)
);

AOI211xp5_ASAP7_75t_SL g1994 ( 
.A1(n_1925),
.A2(n_1775),
.B(n_1783),
.C(n_1902),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1948),
.A2(n_1865),
.B1(n_1912),
.B2(n_1913),
.Y(n_1995)
);

OAI31xp33_ASAP7_75t_L g1996 ( 
.A1(n_1939),
.A2(n_1917),
.A3(n_1881),
.B(n_1882),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1946),
.B(n_1916),
.Y(n_1997)
);

AOI33xp33_ASAP7_75t_L g1998 ( 
.A1(n_1922),
.A2(n_1919),
.A3(n_1884),
.B1(n_1880),
.B2(n_1847),
.B3(n_1909),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1942),
.B(n_1921),
.Y(n_1999)
);

OAI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1928),
.A2(n_1887),
.B1(n_1918),
.B2(n_1881),
.C(n_1890),
.Y(n_2000)
);

INVx4_ASAP7_75t_SL g2001 ( 
.A(n_1985),
.Y(n_2001)
);

AND4x1_ASAP7_75t_L g2002 ( 
.A(n_1966),
.B(n_1951),
.C(n_1945),
.D(n_1831),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1965),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1972),
.B(n_1958),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1968),
.B(n_1943),
.Y(n_2005)
);

BUFx2_ASAP7_75t_L g2006 ( 
.A(n_1990),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1986),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1981),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1986),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1968),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1984),
.Y(n_2011)
);

INVx4_ASAP7_75t_L g2012 ( 
.A(n_1962),
.Y(n_2012)
);

INVx4_ASAP7_75t_SL g2013 ( 
.A(n_1985),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1983),
.Y(n_2014)
);

BUFx2_ASAP7_75t_L g2015 ( 
.A(n_1991),
.Y(n_2015)
);

OA21x2_ASAP7_75t_L g2016 ( 
.A1(n_1967),
.A2(n_1920),
.B(n_1919),
.Y(n_2016)
);

INVx4_ASAP7_75t_SL g2017 ( 
.A(n_1985),
.Y(n_2017)
);

AND4x1_ASAP7_75t_L g2018 ( 
.A(n_1994),
.B(n_1945),
.C(n_1831),
.D(n_1771),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1998),
.B(n_1922),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1961),
.Y(n_2020)
);

INVx2_ASAP7_75t_SL g2021 ( 
.A(n_1989),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1979),
.Y(n_2022)
);

BUFx2_ASAP7_75t_L g2023 ( 
.A(n_1989),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1975),
.B(n_1942),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1998),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_2000),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_1977),
.B(n_1959),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1963),
.A2(n_1887),
.B(n_1853),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1997),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1974),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2003),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_2001),
.B(n_1975),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2001),
.B(n_1976),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2003),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2001),
.B(n_1976),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_2001),
.B(n_2013),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2025),
.B(n_1987),
.Y(n_2037)
);

INVxp67_ASAP7_75t_SL g2038 ( 
.A(n_2006),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2025),
.B(n_1923),
.Y(n_2039)
);

NAND2x1p5_ASAP7_75t_L g2040 ( 
.A(n_2002),
.B(n_1943),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2001),
.B(n_1992),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2006),
.B(n_1923),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2001),
.B(n_1992),
.Y(n_2043)
);

INVxp67_ASAP7_75t_SL g2044 ( 
.A(n_2006),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2016),
.Y(n_2045)
);

NAND3xp33_ASAP7_75t_L g2046 ( 
.A(n_2020),
.B(n_1970),
.C(n_1978),
.Y(n_2046)
);

OAI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_2020),
.A2(n_1971),
.B1(n_1995),
.B2(n_1980),
.C(n_1996),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_2013),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_2019),
.B(n_1973),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_2013),
.B(n_1993),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2003),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2019),
.B(n_1988),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2011),
.Y(n_2053)
);

NOR2x1_ASAP7_75t_L g2054 ( 
.A(n_2005),
.B(n_2012),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_2008),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2023),
.B(n_1964),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2013),
.B(n_2017),
.Y(n_2057)
);

INVxp67_ASAP7_75t_SL g2058 ( 
.A(n_2007),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_SL g2059 ( 
.A(n_2010),
.B(n_1969),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2016),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_2010),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_SL g2062 ( 
.A1(n_2020),
.A2(n_1943),
.B1(n_1982),
.B2(n_1959),
.Y(n_2062)
);

INVx1_ASAP7_75t_SL g2063 ( 
.A(n_2014),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_2012),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_2016),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2024),
.B(n_1999),
.Y(n_2066)
);

BUFx2_ASAP7_75t_SL g2067 ( 
.A(n_2018),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_L g2068 ( 
.A(n_2020),
.B(n_1869),
.C(n_1853),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2038),
.B(n_2030),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2031),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2067),
.B(n_2018),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_2061),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2031),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2061),
.B(n_2004),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2037),
.B(n_2004),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_2040),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2037),
.B(n_2030),
.Y(n_2077)
);

AND2x2_ASAP7_75t_SL g2078 ( 
.A(n_2059),
.B(n_2002),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2038),
.B(n_2029),
.Y(n_2079)
);

OAI21xp33_ASAP7_75t_SL g2080 ( 
.A1(n_2044),
.A2(n_2021),
.B(n_2027),
.Y(n_2080)
);

NOR2x1_ASAP7_75t_L g2081 ( 
.A(n_2067),
.B(n_2012),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2044),
.B(n_2008),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2039),
.B(n_2029),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2034),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2036),
.B(n_2021),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2063),
.B(n_2014),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2045),
.Y(n_2087)
);

NAND3xp33_ASAP7_75t_L g2088 ( 
.A(n_2046),
.B(n_2028),
.C(n_2026),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2039),
.B(n_2029),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2036),
.B(n_2021),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2034),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2055),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2051),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2057),
.B(n_2014),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2045),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2063),
.B(n_2046),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2051),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2055),
.B(n_2015),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2049),
.B(n_2052),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2057),
.B(n_2012),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2053),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2045),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2060),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2053),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2041),
.B(n_2012),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2060),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2041),
.B(n_2043),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2043),
.B(n_2024),
.Y(n_2108)
);

AOI21xp33_ASAP7_75t_SL g2109 ( 
.A1(n_2068),
.A2(n_1771),
.B(n_2015),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2050),
.B(n_2024),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2049),
.B(n_2022),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_2072),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2078),
.B(n_2080),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_2092),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2078),
.B(n_2032),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2078),
.B(n_2032),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2070),
.Y(n_2117)
);

NOR3xp33_ASAP7_75t_L g2118 ( 
.A(n_2088),
.B(n_2068),
.C(n_2047),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2070),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2071),
.B(n_2107),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_2081),
.Y(n_2121)
);

CKINVDCx16_ASAP7_75t_R g2122 ( 
.A(n_2071),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_2081),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2073),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2075),
.B(n_2042),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_2074),
.B(n_2064),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2073),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_2080),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2096),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_2088),
.A2(n_2047),
.B1(n_2027),
.B2(n_2040),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2084),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2110),
.B(n_2033),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_2082),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_2076),
.Y(n_2134)
);

INVx1_ASAP7_75t_SL g2135 ( 
.A(n_2086),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2110),
.B(n_2033),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2087),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2084),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2087),
.A2(n_2059),
.B1(n_2016),
.B2(n_2026),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2108),
.B(n_2035),
.Y(n_2140)
);

HB1xp67_ASAP7_75t_L g2141 ( 
.A(n_2079),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_2128),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_2128),
.A2(n_2077),
.B(n_2098),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2113),
.A2(n_2099),
.B1(n_2109),
.B2(n_2054),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2114),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2112),
.B(n_2056),
.Y(n_2146)
);

OAI21xp33_ASAP7_75t_L g2147 ( 
.A1(n_2118),
.A2(n_2094),
.B(n_2099),
.Y(n_2147)
);

NAND4xp25_ASAP7_75t_L g2148 ( 
.A(n_2118),
.B(n_2054),
.C(n_2100),
.D(n_2105),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2140),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2117),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2129),
.A2(n_2060),
.B1(n_2065),
.B2(n_2109),
.C(n_2028),
.Y(n_2151)
);

INVxp67_ASAP7_75t_SL g2152 ( 
.A(n_2113),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2112),
.B(n_2056),
.Y(n_2153)
);

OAI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2113),
.A2(n_2040),
.B1(n_2052),
.B2(n_2069),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2129),
.B(n_2056),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2122),
.B(n_2100),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_2120),
.Y(n_2157)
);

OAI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_2130),
.A2(n_2040),
.B1(n_2069),
.B2(n_2079),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_2120),
.Y(n_2159)
);

NAND3xp33_ASAP7_75t_L g2160 ( 
.A(n_2130),
.B(n_2064),
.C(n_2065),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2133),
.B(n_2066),
.Y(n_2161)
);

OAI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2139),
.A2(n_2065),
.B1(n_2016),
.B2(n_2076),
.C(n_2062),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2140),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2122),
.B(n_2107),
.Y(n_2164)
);

INVx2_ASAP7_75t_SL g2165 ( 
.A(n_2156),
.Y(n_2165)
);

OR2x2_ASAP7_75t_L g2166 ( 
.A(n_2149),
.B(n_2125),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2142),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_2164),
.B(n_2125),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2157),
.B(n_2132),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2152),
.B(n_2147),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2163),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_L g2172 ( 
.A(n_2148),
.B(n_2133),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2159),
.B(n_2141),
.Y(n_2173)
);

NAND2x1_ASAP7_75t_L g2174 ( 
.A(n_2154),
.B(n_2115),
.Y(n_2174)
);

NOR2x1_ASAP7_75t_L g2175 ( 
.A(n_2145),
.B(n_2133),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_2146),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_2150),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2143),
.B(n_2135),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2153),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2155),
.B(n_2135),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2161),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_2170),
.A2(n_2162),
.B1(n_2137),
.B2(n_2087),
.Y(n_2182)
);

AOI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_2178),
.A2(n_2158),
.B(n_2144),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2174),
.A2(n_2116),
.B1(n_2115),
.B2(n_2160),
.Y(n_2184)
);

NAND3xp33_ASAP7_75t_SL g2185 ( 
.A(n_2172),
.B(n_2123),
.C(n_2121),
.Y(n_2185)
);

XOR2xp5_ASAP7_75t_L g2186 ( 
.A(n_2167),
.B(n_2165),
.Y(n_2186)
);

A2O1A1Ixp33_ASAP7_75t_L g2187 ( 
.A1(n_2168),
.A2(n_2151),
.B(n_2116),
.C(n_2115),
.Y(n_2187)
);

NAND4xp25_ASAP7_75t_L g2188 ( 
.A(n_2175),
.B(n_2126),
.C(n_2121),
.D(n_2123),
.Y(n_2188)
);

AOI221x1_ASAP7_75t_L g2189 ( 
.A1(n_2171),
.A2(n_2158),
.B1(n_2144),
.B2(n_2154),
.C(n_2131),
.Y(n_2189)
);

AOI211xp5_ASAP7_75t_L g2190 ( 
.A1(n_2180),
.A2(n_2116),
.B(n_2076),
.C(n_2134),
.Y(n_2190)
);

AOI22xp33_ASAP7_75t_L g2191 ( 
.A1(n_2180),
.A2(n_2137),
.B1(n_2095),
.B2(n_2103),
.Y(n_2191)
);

NAND4xp25_ASAP7_75t_L g2192 ( 
.A(n_2169),
.B(n_2132),
.C(n_2136),
.D(n_2140),
.Y(n_2192)
);

NAND3x1_ASAP7_75t_L g2193 ( 
.A(n_2173),
.B(n_2076),
.C(n_2094),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2176),
.A2(n_2137),
.B1(n_2095),
.B2(n_2103),
.C(n_2106),
.Y(n_2194)
);

OAI21xp33_ASAP7_75t_L g2195 ( 
.A1(n_2173),
.A2(n_2136),
.B(n_2132),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2186),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2184),
.Y(n_2197)
);

AOI221xp5_ASAP7_75t_L g2198 ( 
.A1(n_2182),
.A2(n_2179),
.B1(n_2177),
.B2(n_2181),
.C(n_2095),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2192),
.Y(n_2199)
);

AOI211xp5_ASAP7_75t_L g2200 ( 
.A1(n_2183),
.A2(n_2166),
.B(n_2134),
.C(n_2177),
.Y(n_2200)
);

OAI32xp33_ASAP7_75t_L g2201 ( 
.A1(n_2188),
.A2(n_2138),
.A3(n_2117),
.B1(n_2119),
.B2(n_2124),
.Y(n_2201)
);

AOI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_2194),
.A2(n_2102),
.B1(n_2106),
.B2(n_2134),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2187),
.B(n_2136),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2196),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2197),
.Y(n_2205)
);

NAND2xp33_ASAP7_75t_L g2206 ( 
.A(n_2203),
.B(n_2193),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2200),
.B(n_2195),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2201),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2199),
.B(n_2185),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2202),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2198),
.A2(n_2189),
.B(n_2190),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2205),
.Y(n_2212)
);

O2A1O1Ixp33_ASAP7_75t_L g2213 ( 
.A1(n_2211),
.A2(n_2191),
.B(n_2138),
.C(n_2131),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2204),
.B(n_2105),
.Y(n_2214)
);

OAI322xp33_ASAP7_75t_L g2215 ( 
.A1(n_2208),
.A2(n_2127),
.A3(n_2124),
.B1(n_2119),
.B2(n_2102),
.C1(n_2058),
.C2(n_2083),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2207),
.B(n_2085),
.Y(n_2216)
);

HB1xp67_ASAP7_75t_L g2217 ( 
.A(n_2210),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2206),
.A2(n_2127),
.B1(n_2058),
.B2(n_2104),
.C(n_2097),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2212),
.Y(n_2219)
);

AOI221x1_ASAP7_75t_L g2220 ( 
.A1(n_2216),
.A2(n_2209),
.B1(n_2101),
.B2(n_2104),
.C(n_2097),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2214),
.B(n_2209),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2217),
.Y(n_2222)
);

NOR3xp33_ASAP7_75t_SL g2223 ( 
.A(n_2219),
.B(n_2222),
.C(n_2215),
.Y(n_2223)
);

OAI211xp5_ASAP7_75t_SL g2224 ( 
.A1(n_2223),
.A2(n_2213),
.B(n_2218),
.C(n_2221),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2224),
.Y(n_2225)
);

NAND4xp25_ASAP7_75t_L g2226 ( 
.A(n_2224),
.B(n_2221),
.C(n_2220),
.D(n_2062),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_2225),
.Y(n_2227)
);

AOI21xp33_ASAP7_75t_L g2228 ( 
.A1(n_2226),
.A2(n_2009),
.B(n_2007),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_2227),
.Y(n_2229)
);

AOI22x1_ASAP7_75t_L g2230 ( 
.A1(n_2228),
.A2(n_2085),
.B1(n_2090),
.B2(n_2093),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2229),
.A2(n_2048),
.B1(n_2083),
.B2(n_2089),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2231),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_R g2233 ( 
.A1(n_2232),
.A2(n_2230),
.B1(n_2091),
.B2(n_2101),
.Y(n_2233)
);

O2A1O1Ixp33_ASAP7_75t_L g2234 ( 
.A1(n_2233),
.A2(n_2093),
.B(n_2091),
.C(n_2048),
.Y(n_2234)
);

AOI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2234),
.A2(n_2090),
.B1(n_2048),
.B2(n_2009),
.C(n_2007),
.Y(n_2235)
);

AOI211xp5_ASAP7_75t_L g2236 ( 
.A1(n_2235),
.A2(n_2089),
.B(n_2111),
.C(n_2108),
.Y(n_2236)
);


endmodule