module fake_jpeg_7179_n_116 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_28),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_27),
.B1(n_16),
.B2(n_26),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_43),
.B1(n_18),
.B2(n_21),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_46),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_25),
.B1(n_26),
.B2(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_33),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_62),
.Y(n_68)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_59),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_0),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_34),
.B1(n_26),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_18),
.B1(n_12),
.B2(n_37),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_40),
.B(n_21),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_25),
.C(n_24),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_24),
.B1(n_15),
.B2(n_14),
.Y(n_64)
);

XNOR2x1_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_41),
.Y(n_72)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_76),
.B1(n_60),
.B2(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_10),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_54),
.C(n_65),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_86),
.C(n_89),
.Y(n_92)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_54),
.B(n_59),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_58),
.Y(n_94)
);

OAI322xp33_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_73),
.A3(n_62),
.B1(n_19),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_80),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g99 ( 
.A(n_95),
.B(n_86),
.C(n_83),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_88),
.B1(n_87),
.B2(n_89),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_83),
.C(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_97),
.C(n_100),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g104 ( 
.A(n_99),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_9),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_2),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_107),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

OAI221xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_4),
.B1(n_5),
.B2(n_32),
.C(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_111),
.B(n_5),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_113),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_110),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_112),
.Y(n_116)
);


endmodule