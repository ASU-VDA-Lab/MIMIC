module fake_jpeg_1420_n_226 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g55 ( 
.A(n_14),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

INVx11_ASAP7_75t_SL g84 ( 
.A(n_68),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_66),
.B1(n_59),
.B2(n_55),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_96),
.B1(n_76),
.B2(n_63),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_57),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_66),
.B1(n_59),
.B2(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_79),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_55),
.B1(n_63),
.B2(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_70),
.B1(n_86),
.B2(n_67),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_88),
.B(n_56),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_112),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_111),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_88),
.B1(n_70),
.B2(n_79),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_109),
.B1(n_113),
.B2(n_117),
.Y(n_127)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_118),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_88),
.B1(n_56),
.B2(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_73),
.Y(n_111)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_120),
.Y(n_140)
);

CKINVDCx12_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_98),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_98),
.B1(n_99),
.B2(n_94),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_77),
.B1(n_60),
.B2(n_81),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_95),
.B1(n_98),
.B2(n_65),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_143),
.B1(n_146),
.B2(n_49),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_129),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_0),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2x1p5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_54),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_78),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_61),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_44),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_77),
.B1(n_81),
.B2(n_60),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_114),
.C(n_60),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_171),
.C(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_61),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_156),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_164),
.B(n_158),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_169),
.B(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_162),
.B1(n_153),
.B2(n_164),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_141),
.B1(n_135),
.B2(n_8),
.Y(n_176)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_162)
);

CKINVDCx6p67_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_2),
.B(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_38),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_4),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_5),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_35),
.C(n_32),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_173),
.B(n_17),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_182),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_140),
.B(n_135),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_179),
.B(n_150),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_184),
.B1(n_174),
.B2(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_154),
.B1(n_12),
.B2(n_13),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_31),
.C(n_29),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_180),
.C(n_187),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_28),
.B(n_27),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_26),
.C(n_24),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_22),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_171),
.B(n_165),
.C(n_150),
.D(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_195),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

NAND5xp2_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_11),
.C(n_14),
.D(n_15),
.E(n_16),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_15),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_182),
.C(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_199),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_193),
.C(n_200),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_213),
.B1(n_205),
.B2(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_193),
.C(n_172),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_206),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_204),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_192),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_215),
.C(n_183),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_181),
.B1(n_190),
.B2(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_184),
.C(n_18),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_17),
.B(n_18),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.C(n_161),
.Y(n_225)
);

XNOR2x2_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_19),
.Y(n_226)
);


endmodule