module real_jpeg_27522_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_343, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_343;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_23),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_49),
.B1(n_58),
.B2(n_60),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_1),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_117),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_3),
.A2(n_58),
.B1(n_60),
.B2(n_117),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_117),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_4),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_28),
.B1(n_32),
.B2(n_122),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_122),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_4),
.A2(n_58),
.B1(n_60),
.B2(n_122),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_23),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_38),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_38),
.B1(n_58),
.B2(n_60),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_28),
.B1(n_32),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_8),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_115),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_115),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_115),
.Y(n_206)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_9),
.B(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_9),
.B(n_32),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_32),
.B(n_164),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_120),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_9),
.A2(n_58),
.B(n_61),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_9),
.B(n_78),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_9),
.A2(n_98),
.B1(n_106),
.B2(n_214),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_10),
.A2(n_47),
.B1(n_58),
.B2(n_60),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_47),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_12),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_12),
.A2(n_25),
.B1(n_58),
.B2(n_60),
.Y(n_161)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_341),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_83),
.B(n_339),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_20),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_21),
.A2(n_45),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_22),
.A2(n_34),
.B(n_82),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_22),
.A2(n_27),
.B(n_34),
.Y(n_341)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_27),
.B(n_30),
.C(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_30),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g119 ( 
.A(n_23),
.B(n_120),
.CON(n_119),
.SN(n_119)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_27),
.A2(n_34),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_28),
.A2(n_32),
.B1(n_67),
.B2(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_28),
.A2(n_35),
.B1(n_119),
.B2(n_134),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_28),
.A2(n_54),
.A3(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_30),
.B(n_32),
.Y(n_134)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_33),
.A2(n_46),
.B(n_50),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_34),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_40),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_75),
.C(n_80),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_41),
.A2(n_42),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.C(n_64),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_43),
.A2(n_44),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_45),
.A2(n_50),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_45),
.A2(n_50),
.B1(n_128),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_51),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_51),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_51),
.A2(n_64),
.B1(n_307),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_62),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_52),
.A2(n_62),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_52),
.A2(n_57),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_52),
.A2(n_172),
.B(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_52),
.A2(n_57),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_52),
.A2(n_57),
.B1(n_171),
.B2(n_190),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_52),
.A2(n_57),
.B1(n_93),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_52),
.A2(n_110),
.B(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_55),
.B(n_73),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_55),
.A2(n_56),
.B(n_120),
.C(n_192),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_57),
.B(n_120),
.Y(n_212)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_60),
.B(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_63),
.B(n_111),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_64),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_77),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_71),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_71),
.B1(n_114),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_66),
.A2(n_71),
.B1(n_147),
.B2(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_66),
.B(n_70),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_66),
.A2(n_71),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_69),
.A2(n_78),
.B(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_77),
.A2(n_79),
.B(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_77),
.A2(n_257),
.B(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_80),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_332),
.B(n_338),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_302),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_343),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_283),
.B(n_301),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_261),
.B(n_282),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_153),
.B(n_238),
.C(n_260),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_139),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_89),
.B(n_139),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_123),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_107),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_91),
.B(n_107),
.C(n_123),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_92),
.B(n_97),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_94),
.B(n_182),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B(n_103),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_102),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_98),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_98),
.A2(n_206),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_98),
.A2(n_137),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_99),
.A2(n_104),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_99),
.A2(n_138),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_136),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_106),
.B(n_120),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_118),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_132),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_125),
.B(n_130),
.C(n_132),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.Y(n_144)
);

INVx5_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_138),
.B(n_161),
.Y(n_201)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_140),
.A2(n_141),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_151),
.B(n_201),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_237),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_230),
.B(n_236),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_183),
.B(n_229),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_173),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_157),
.B(n_173),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.C(n_169),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_158),
.A2(n_159),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_162),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_161),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_180),
.C(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_223),
.B(n_228),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_202),
.B(n_222),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_186),
.B(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_210),
.B(n_221),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_208),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_216),
.B(n_220),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_240),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_258),
.B2(n_259),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_249),
.C(n_259),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_281),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_275),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_270),
.C(n_272),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_277),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_295),
.B(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_285),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_299),
.B2(n_300),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_294),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_294),
.C(n_300),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_293),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_292),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_304),
.C(n_314),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_304),
.B1(n_305),
.B2(n_329),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_293),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_313),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_322),
.C(n_323),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_315),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);


endmodule