module fake_jpeg_7252_n_56 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_56);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_56;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx6_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_31),
.B1(n_13),
.B2(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_15),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_6),
.B(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_10),
.B1(n_18),
.B2(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_5),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.C(n_39),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_16),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_52),
.B(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

AOI322xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_44),
.A3(n_39),
.B1(n_37),
.B2(n_47),
.C1(n_17),
.C2(n_22),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_49),
.Y(n_56)
);


endmodule