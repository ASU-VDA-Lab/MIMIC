module fake_jpeg_28833_n_150 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_2),
.Y(n_89)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_1),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_2),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_60),
.Y(n_79)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_87),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_49),
.B1(n_62),
.B2(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_83),
.B1(n_66),
.B2(n_57),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_59),
.B1(n_68),
.B2(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_56),
.B1(n_69),
.B2(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_65),
.B1(n_68),
.B2(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_9),
.B1(n_15),
.B2(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_55),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_4),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_5),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_54),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_6),
.B(n_8),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_28),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_117),
.B1(n_40),
.B2(n_42),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_97),
.C(n_104),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_32),
.C(n_36),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_34),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_43),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_124)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_132),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_124),
.C(n_122),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_37),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_111),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_38),
.B(n_39),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_130),
.A2(n_135),
.B(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_44),
.B1(n_46),
.B2(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_141),
.B(n_135),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

BUFx4f_ASAP7_75t_SL g145 ( 
.A(n_142),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_144),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_136),
.B(n_134),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_143),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_129),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_128),
.Y(n_150)
);


endmodule