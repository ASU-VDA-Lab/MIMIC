module fake_netlist_1_6716_n_755 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_755);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_755;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_476;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g82 ( .A(n_33), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_42), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_73), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_5), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_69), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_41), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_52), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_0), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_48), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_80), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_79), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_27), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_31), .Y(n_98) );
NOR2xp33_ASAP7_75t_L g99 ( .A(n_3), .B(n_14), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_57), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_54), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_75), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_23), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_12), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_53), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_18), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_77), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_70), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_61), .Y(n_110) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_0), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_35), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_60), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_45), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_66), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_20), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_26), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_38), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_17), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_44), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_4), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_63), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_16), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_74), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_43), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_62), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_28), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_72), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_130), .B(n_30), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_124), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_84), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_130), .Y(n_139) );
INVxp67_ASAP7_75t_SL g140 ( .A(n_85), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_100), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_118), .B(n_1), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_126), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_118), .B(n_2), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_94), .B(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_88), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_123), .B(n_5), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_111), .B(n_6), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_84), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_123), .B(n_6), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_91), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_103), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_92), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_103), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
XNOR2xp5_ASAP7_75t_L g165 ( .A(n_86), .B(n_7), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_102), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_95), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_90), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_96), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_96), .B(n_8), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_125), .B(n_9), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_109), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_109), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_97), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_125), .B(n_9), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_121), .A2(n_104), .B1(n_119), .B2(n_122), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_104), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_133), .B(n_131), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_141), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_133), .B(n_114), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_140), .B(n_122), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_141), .Y(n_189) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_152), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_157), .B(n_107), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_149), .A2(n_176), .B1(n_137), .B2(n_164), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_157), .B(n_129), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_157), .B(n_129), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_162), .B(n_106), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_143), .B(n_119), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_135), .B(n_128), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_171), .B(n_128), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_164), .B(n_143), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_132), .B(n_108), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_146), .B(n_117), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_146), .B(n_105), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_134), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_147), .B(n_113), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_134), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_138), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_145), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_150), .A2(n_99), .B1(n_97), .B2(n_116), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_132), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_150), .B(n_110), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_138), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_138), .Y(n_228) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_170), .A2(n_105), .B(n_110), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_151), .A2(n_101), .B1(n_116), .B2(n_115), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_151), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_145), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_171), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_159), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_161), .B(n_115), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_167), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_175), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_139), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_175), .B(n_101), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_163), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_174), .B(n_113), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_155), .A2(n_112), .B1(n_127), .B2(n_120), .Y(n_246) );
BUFx4f_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_233), .A2(n_155), .B1(n_160), .B2(n_136), .Y(n_248) );
AOI21xp33_ASAP7_75t_L g249 ( .A1(n_214), .A2(n_154), .B(n_174), .Y(n_249) );
INVx8_ASAP7_75t_L g250 ( .A(n_178), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_246), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_204), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_185), .A2(n_153), .B(n_142), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_190), .B(n_156), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_204), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_178), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_235), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
OR2x2_ASAP7_75t_SL g260 ( .A(n_208), .B(n_160), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_211), .A2(n_166), .B1(n_177), .B2(n_148), .Y(n_261) );
NOR2x2_ASAP7_75t_L g262 ( .A(n_211), .B(n_165), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_231), .B(n_166), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_234), .Y(n_264) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_240), .A2(n_165), .B1(n_172), .B2(n_173), .C(n_144), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_236), .Y(n_266) );
AND2x4_ASAP7_75t_SL g267 ( .A(n_182), .B(n_168), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_236), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_231), .B(n_168), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_212), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_238), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_194), .B(n_168), .Y(n_274) );
OAI21xp33_ASAP7_75t_L g275 ( .A1(n_243), .A2(n_139), .B(n_93), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_182), .A2(n_87), .B1(n_82), .B2(n_139), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_242), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_243), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_202), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_208), .B(n_219), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_219), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_186), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_239), .B(n_139), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_239), .B(n_139), .Y(n_284) );
CKINVDCx6p67_ASAP7_75t_R g285 ( .A(n_186), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_241), .B(n_40), .Y(n_286) );
NOR3xp33_ASAP7_75t_SL g287 ( .A(n_196), .B(n_10), .C(n_11), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_241), .B(n_49), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_186), .B(n_14), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_244), .B(n_50), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_186), .B(n_15), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_217), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_217), .B(n_15), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_203), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_185), .A2(n_51), .B(n_78), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_191), .B(n_16), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_195), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_185), .B(n_47), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_242), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_191), .B(n_17), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_203), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_244), .B(n_19), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_235), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_217), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_245), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_235), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_225), .B(n_22), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_218), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_191), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_193), .B(n_24), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_225), .B(n_25), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_225), .B(n_29), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_229), .B(n_32), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_245), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_218), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_229), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_193), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_193), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_242), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_280), .B(n_229), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_315), .B(n_255), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_251), .A2(n_224), .B1(n_205), .B2(n_210), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_252), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_316), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_257), .Y(n_327) );
AND2x2_ASAP7_75t_SL g328 ( .A(n_247), .B(n_205), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_247), .A2(n_224), .B1(n_205), .B2(n_230), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_259), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_253), .A2(n_224), .B(n_200), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_264), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_273), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_288), .A2(n_198), .B(n_237), .C(n_232), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_254), .A2(n_200), .B(n_179), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_266), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_268), .Y(n_337) );
NAND2x1_ASAP7_75t_SL g338 ( .A(n_290), .B(n_232), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_293), .A2(n_210), .B1(n_179), .B2(n_216), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_270), .B(n_223), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_254), .B(n_222), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_295), .A2(n_222), .B(n_220), .C(n_210), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_258), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_258), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_281), .B(n_210), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_187), .B(n_183), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_258), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_272), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_278), .B(n_220), .Y(n_350) );
BUFx4_ASAP7_75t_SL g351 ( .A(n_297), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_318), .A2(n_184), .B(n_215), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_285), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_273), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_302), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_314), .A2(n_184), .B(n_215), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_278), .B(n_206), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_256), .A2(n_206), .B(n_213), .C(n_209), .Y(n_360) );
INVx3_ASAP7_75t_SL g361 ( .A(n_297), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_311), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_305), .B(n_206), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_311), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_269), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_282), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_267), .B(n_183), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_314), .A2(n_207), .B(n_188), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_290), .B(n_207), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_263), .B(n_227), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_292), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_277), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_283), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_292), .B(n_227), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_250), .B(n_209), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_306), .B(n_187), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_301), .A2(n_213), .B1(n_197), .B2(n_188), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_283), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_334), .A2(n_249), .B(n_275), .C(n_294), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_321), .B(n_298), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_358), .A2(n_291), .B(n_286), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_368), .A2(n_291), .B(n_286), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
CKINVDCx6p67_ASAP7_75t_R g385 ( .A(n_361), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_354), .B(n_250), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_330), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
OAI21x1_ASAP7_75t_SL g389 ( .A1(n_330), .A2(n_296), .B(n_303), .Y(n_389) );
O2A1O1Ixp5_ASAP7_75t_L g390 ( .A1(n_370), .A2(n_299), .B(n_303), .C(n_289), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
AO31x2_ASAP7_75t_L g393 ( .A1(n_343), .A2(n_317), .A3(n_289), .B(n_284), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_321), .B(n_301), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_332), .Y(n_395) );
CKINVDCx11_ASAP7_75t_R g396 ( .A(n_361), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_340), .A2(n_248), .B1(n_265), .B2(n_250), .C(n_261), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_332), .A2(n_313), .B(n_312), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_331), .A2(n_308), .B(n_284), .Y(n_400) );
AOI21x1_ASAP7_75t_L g401 ( .A1(n_377), .A2(n_221), .B(n_228), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g402 ( .A1(n_365), .A2(n_249), .B(n_287), .C(n_274), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_362), .A2(n_221), .B(n_228), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_350), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_354), .Y(n_405) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_362), .A2(n_226), .B(n_201), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_362), .A2(n_226), .B(n_201), .Y(n_407) );
OR2x6_ASAP7_75t_L g408 ( .A(n_354), .B(n_301), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_336), .Y(n_409) );
OAI21x1_ASAP7_75t_L g410 ( .A1(n_364), .A2(n_307), .B(n_304), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_344), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_364), .A2(n_180), .B(n_189), .Y(n_412) );
BUFx2_ASAP7_75t_SL g413 ( .A(n_351), .Y(n_413) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_325), .Y(n_414) );
OR2x6_ASAP7_75t_L g415 ( .A(n_408), .B(n_355), .Y(n_415) );
INVx4_ASAP7_75t_SL g416 ( .A(n_408), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_381), .B(n_260), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_400), .A2(n_364), .B(n_335), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_380), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_413), .A2(n_355), .B1(n_353), .B2(n_322), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_398), .A2(n_348), .B(n_344), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_413), .Y(n_422) );
OAI222xp33_ASAP7_75t_L g423 ( .A1(n_408), .A2(n_350), .B1(n_371), .B2(n_353), .C1(n_276), .C2(n_322), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_405), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_374), .B(n_342), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_405), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_404), .A2(n_337), .B1(n_341), .B2(n_349), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g428 ( .A1(n_397), .A2(n_376), .B(n_322), .C(n_262), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_387), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_394), .B(n_376), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_396), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g432 ( .A1(n_397), .A2(n_338), .B(n_366), .C(n_367), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_379), .B(n_360), .C(n_346), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_394), .B(n_365), .Y(n_434) );
OAI21x1_ASAP7_75t_L g435 ( .A1(n_400), .A2(n_336), .B(n_341), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_398), .A2(n_345), .B(n_348), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_398), .A2(n_345), .B(n_348), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_381), .B(n_327), .Y(n_438) );
OAI22xp5_ASAP7_75t_SL g439 ( .A1(n_414), .A2(n_279), .B1(n_328), .B2(n_327), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_387), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_380), .A2(n_338), .B1(n_357), .B2(n_324), .C(n_333), .Y(n_441) );
AO31x2_ASAP7_75t_L g442 ( .A1(n_395), .A2(n_349), .A3(n_337), .B(n_339), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_408), .B(n_323), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_419), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_429), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_432), .A2(n_408), .B(n_389), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_429), .B(n_395), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_435), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_416), .B(n_405), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_435), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_440), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_434), .B(n_409), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_443), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_421), .A2(n_389), .B(n_401), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_417), .B(n_414), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_427), .B(n_409), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_393), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_442), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_438), .B(n_388), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_426), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_388), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_442), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_444), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_415), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_415), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_417), .B(n_385), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_442), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_442), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_439), .B(n_414), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_415), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_446), .B(n_393), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_457), .B(n_425), .C(n_420), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_446), .B(n_393), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_476), .A2(n_462), .B1(n_445), .B2(n_441), .C(n_480), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_464), .A2(n_433), .B(n_423), .Y(n_486) );
INVx5_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_450), .Y(n_488) );
OAI31xp33_ASAP7_75t_L g489 ( .A1(n_471), .A2(n_386), .A3(n_329), .B(n_392), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_465), .B(n_393), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_448), .B(n_393), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_448), .B(n_393), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_481), .B(n_388), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_455), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_466), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_471), .A2(n_422), .B1(n_385), .B2(n_431), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_455), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_465), .B(n_375), .C(n_363), .D(n_197), .Y(n_499) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_464), .Y(n_500) );
AO31x2_ASAP7_75t_L g501 ( .A1(n_466), .A2(n_437), .A3(n_436), .B(n_384), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_452), .B(n_388), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_452), .Y(n_503) );
AND3x1_ASAP7_75t_L g504 ( .A(n_469), .B(n_431), .C(n_422), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_467), .B(n_392), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_481), .B(n_392), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_467), .B(n_392), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_481), .B(n_410), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_466), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_453), .B(n_410), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_479), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_472), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_453), .B(n_373), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_450), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_479), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_472), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_454), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_469), .B(n_357), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_470), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_472), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_474), .B(n_403), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_477), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_474), .B(n_378), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_477), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_470), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_456), .B(n_373), .Y(n_529) );
OAI31xp33_ASAP7_75t_L g530 ( .A1(n_447), .A2(n_323), .A3(n_326), .B(n_333), .Y(n_530) );
AOI31xp33_ASAP7_75t_L g531 ( .A1(n_473), .A2(n_326), .A3(n_359), .B(n_378), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_478), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_482), .B(n_478), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_531), .B(n_447), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_494), .B(n_475), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_498), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_482), .B(n_468), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_505), .B(n_475), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_505), .B(n_468), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_507), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_483), .B(n_463), .C(n_460), .Y(n_544) );
NOR2xp33_ASAP7_75t_R g545 ( .A(n_487), .B(n_463), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_487), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_507), .B(n_502), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_484), .B(n_460), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_484), .B(n_458), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_497), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_485), .B(n_458), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_491), .B(n_456), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_516), .Y(n_554) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_507), .B(n_451), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_491), .B(n_451), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_496), .B(n_227), .C(n_454), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_502), .B(n_459), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_503), .B(n_449), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_487), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_487), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_515), .B(n_459), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_515), .B(n_459), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_496), .B(n_459), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_499), .B(n_461), .Y(n_566) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_486), .B(n_461), .C(n_454), .D(n_390), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_492), .B(n_461), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_514), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_525), .B(n_490), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_492), .B(n_449), .Y(n_572) );
OR2x6_ASAP7_75t_L g573 ( .A(n_523), .B(n_449), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_525), .B(n_399), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_489), .B(n_390), .C(n_189), .D(n_181), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_529), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_490), .B(n_399), .Y(n_577) );
OR2x6_ASAP7_75t_L g578 ( .A(n_523), .B(n_403), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_529), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_487), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_527), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_527), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_508), .B(n_399), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_500), .B(n_398), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_487), .B(n_407), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_488), .B(n_407), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_495), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_530), .B(n_227), .C(n_199), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_495), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_488), .B(n_411), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_488), .B(n_411), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_512), .B(n_406), .Y(n_592) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_518), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_513), .B(n_406), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_506), .B(n_411), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_519), .B(n_323), .C(n_372), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_552), .B(n_520), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_538), .B(n_520), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_547), .B(n_528), .Y(n_600) );
INVx6_ASAP7_75t_L g601 ( .A(n_585), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_569), .B(n_520), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_541), .B(n_528), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_550), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_571), .B(n_513), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_551), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_587), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_558), .B(n_509), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_556), .B(n_517), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_568), .B(n_509), .Y(n_610) );
INVx5_ASAP7_75t_L g611 ( .A(n_578), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_556), .B(n_524), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_563), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_576), .B(n_524), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_579), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_570), .B(n_517), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_553), .B(n_521), .Y(n_617) );
INVx2_ASAP7_75t_SL g618 ( .A(n_545), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_553), .B(n_521), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_584), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_566), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_554), .B(n_533), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_557), .A2(n_504), .B(n_493), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_554), .B(n_522), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_537), .B(n_533), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_540), .B(n_522), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_540), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_548), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_548), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_562), .B(n_526), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_549), .B(n_526), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_572), .B(n_534), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_549), .B(n_511), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_552), .B(n_533), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_581), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_589), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_542), .B(n_511), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_543), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_535), .B(n_534), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_535), .B(n_532), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_559), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_564), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_572), .B(n_565), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_577), .B(n_532), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_582), .B(n_510), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_544), .A2(n_493), .B(n_506), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_596), .B(n_510), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_555), .B(n_493), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_583), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_594), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_628), .B(n_584), .Y(n_652) );
NOR2xp33_ASAP7_75t_SL g653 ( .A(n_618), .B(n_546), .Y(n_653) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_619), .A2(n_536), .B1(n_561), .B2(n_580), .C1(n_560), .C2(n_588), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_619), .A2(n_596), .B1(n_567), .B2(n_573), .Y(n_655) );
OAI32xp33_ASAP7_75t_L g656 ( .A1(n_639), .A2(n_592), .A3(n_574), .B1(n_575), .B2(n_594), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_622), .B(n_573), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_597), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_629), .B(n_595), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_604), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_600), .B(n_573), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_630), .B(n_591), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_644), .B(n_592), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_622), .A2(n_578), .B(n_585), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_618), .B(n_586), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_625), .Y(n_666) );
NOR2xp67_ASAP7_75t_SL g667 ( .A(n_611), .B(n_590), .Y(n_667) );
NAND3xp33_ASAP7_75t_SL g668 ( .A(n_624), .B(n_578), .C(n_523), .Y(n_668) );
OAI32xp33_ASAP7_75t_L g669 ( .A1(n_598), .A2(n_523), .A3(n_586), .B1(n_391), .B2(n_384), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_621), .B(n_493), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_635), .A2(n_593), .B1(n_518), .B2(n_412), .Y(n_671) );
OAI32xp33_ASAP7_75t_L g672 ( .A1(n_598), .A2(n_384), .A3(n_391), .B1(n_593), .B2(n_181), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_621), .A2(n_227), .B1(n_518), .B2(n_199), .C(n_192), .Y(n_673) );
OAI32xp33_ASAP7_75t_SL g674 ( .A1(n_634), .A2(n_501), .A3(n_36), .B1(n_37), .B2(n_55), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_599), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_635), .A2(n_518), .B1(n_391), .B2(n_401), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_606), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_608), .B(n_501), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_608), .A2(n_518), .B(n_180), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_611), .B(n_34), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_650), .B(n_501), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_613), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_636), .Y(n_683) );
AOI22xp5_ASAP7_75t_SL g684 ( .A1(n_649), .A2(n_501), .B1(n_333), .B2(n_372), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_610), .B(n_501), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_615), .B(n_199), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_610), .B(n_412), .Y(n_687) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_611), .B(n_56), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_626), .A2(n_372), .B1(n_199), .B2(n_192), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_609), .B(n_58), .Y(n_690) );
CKINVDCx16_ASAP7_75t_R g691 ( .A(n_653), .Y(n_691) );
INVx3_ASAP7_75t_L g692 ( .A(n_685), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_675), .A2(n_648), .B(n_647), .Y(n_693) );
AO22x2_ASAP7_75t_L g694 ( .A1(n_668), .A2(n_623), .B1(n_602), .B2(n_642), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_681), .B(n_643), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_660), .Y(n_696) );
OAI22x1_ASAP7_75t_L g697 ( .A1(n_675), .A2(n_611), .B1(n_603), .B2(n_642), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_655), .A2(n_601), .B1(n_638), .B2(n_605), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_661), .B(n_643), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_652), .B(n_631), .Y(n_700) );
AOI321xp33_ASAP7_75t_L g701 ( .A1(n_655), .A2(n_656), .A3(n_657), .B1(n_665), .B2(n_669), .C(n_690), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_677), .Y(n_702) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_668), .B(n_612), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_682), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_683), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_666), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_654), .A2(n_601), .B1(n_631), .B2(n_617), .Y(n_707) );
AOI222xp33_ASAP7_75t_L g708 ( .A1(n_678), .A2(n_620), .B1(n_627), .B2(n_632), .C1(n_641), .C2(n_640), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_663), .B(n_651), .Y(n_709) );
XNOR2xp5_ASAP7_75t_L g710 ( .A(n_662), .B(n_633), .Y(n_710) );
AOI31xp33_ASAP7_75t_L g711 ( .A1(n_664), .A2(n_614), .A3(n_616), .B(n_645), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_658), .A2(n_601), .B1(n_651), .B2(n_646), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_670), .B(n_637), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_686), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_659), .B(n_637), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_698), .A2(n_690), .B1(n_687), .B2(n_671), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_715), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_691), .Y(n_718) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_701), .A2(n_679), .B(n_673), .C(n_672), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_706), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_708), .B(n_684), .Y(n_721) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_703), .B(n_667), .Y(n_722) );
AOI322xp5_ASAP7_75t_L g723 ( .A1(n_707), .A2(n_674), .A3(n_673), .B1(n_607), .B2(n_689), .C1(n_680), .C2(n_688), .Y(n_723) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_693), .B(n_676), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_696), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_694), .A2(n_607), .B1(n_192), .B2(n_199), .C(n_369), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_702), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_711), .A2(n_328), .B(n_382), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_704), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_697), .A2(n_383), .B(n_382), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g731 ( .A1(n_718), .A2(n_694), .B1(n_697), .B2(n_705), .C1(n_712), .C2(n_692), .Y(n_731) );
XNOR2x1_ASAP7_75t_L g732 ( .A(n_720), .B(n_694), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_722), .A2(n_712), .B1(n_692), .B2(n_710), .C(n_695), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_720), .A2(n_692), .B(n_700), .Y(n_734) );
OAI211xp5_ASAP7_75t_L g735 ( .A1(n_723), .A2(n_714), .B(n_713), .C(n_709), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_717), .B(n_714), .Y(n_736) );
AO22x1_ASAP7_75t_L g737 ( .A1(n_721), .A2(n_709), .B1(n_699), .B2(n_356), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_719), .B(n_356), .C(n_383), .Y(n_738) );
O2A1O1Ixp33_ASAP7_75t_L g739 ( .A1(n_724), .A2(n_319), .B(n_347), .C(n_352), .Y(n_739) );
NAND5xp2_ASAP7_75t_L g740 ( .A(n_731), .B(n_726), .C(n_728), .D(n_716), .E(n_730), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_732), .A2(n_729), .B1(n_727), .B2(n_725), .Y(n_741) );
AO22x2_ASAP7_75t_L g742 ( .A1(n_735), .A2(n_59), .B1(n_64), .B2(n_65), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g743 ( .A(n_734), .B(n_348), .Y(n_743) );
NAND4xp75_ASAP7_75t_L g744 ( .A(n_736), .B(n_67), .C(n_68), .D(n_71), .Y(n_744) );
AND3x4_ASAP7_75t_L g745 ( .A(n_740), .B(n_738), .C(n_733), .Y(n_745) );
NAND3xp33_ASAP7_75t_SL g746 ( .A(n_741), .B(n_739), .C(n_737), .Y(n_746) );
AOI22xp5_ASAP7_75t_SL g747 ( .A1(n_743), .A2(n_81), .B1(n_192), .B2(n_345), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_747), .Y(n_748) );
OR3x1_ASAP7_75t_L g749 ( .A(n_746), .B(n_742), .C(n_744), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_748), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_749), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_750), .Y(n_752) );
BUFx4_ASAP7_75t_R g753 ( .A(n_752), .Y(n_753) );
OA22x2_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_751), .B1(n_745), .B2(n_320), .Y(n_754) );
OAI321xp33_ASAP7_75t_L g755 ( .A1(n_754), .A2(n_192), .A3(n_300), .B1(n_345), .B2(n_348), .C(n_751), .Y(n_755) );
endmodule