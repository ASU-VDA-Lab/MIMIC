module fake_jpeg_4877_n_261 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_36),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_41),
.B1(n_25),
.B2(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_43),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_26),
.C(n_22),
.Y(n_56)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_25),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_47),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_51),
.Y(n_115)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_24),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_56),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_62),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_71),
.B(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_69),
.Y(n_117)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_70),
.Y(n_101)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_35),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_32),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_82),
.Y(n_96)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_34),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_32),
.B(n_24),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_89),
.B1(n_26),
.B2(n_27),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_40),
.B(n_16),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_88),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_28),
.B(n_15),
.C(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_104),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_28),
.B(n_15),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_28),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_28),
.B(n_15),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_75),
.A2(n_28),
.B1(n_15),
.B2(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_119),
.B1(n_61),
.B2(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_53),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_120),
.B(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_124),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_147),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_55),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_76),
.B1(n_80),
.B2(n_57),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_86),
.B1(n_63),
.B2(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_144),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

HAxp5_ASAP7_75t_SL g141 ( 
.A(n_97),
.B(n_28),
.CON(n_141),
.SN(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_83),
.C(n_63),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_83),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_91),
.A2(n_114),
.B1(n_106),
.B2(n_102),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_91),
.A2(n_99),
.B1(n_106),
.B2(n_114),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_15),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_169),
.Y(n_196)
);

BUFx12f_ASAP7_75t_SL g163 ( 
.A(n_139),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_134),
.B(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_172),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_107),
.B1(n_93),
.B2(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_107),
.B1(n_108),
.B2(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_178),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_103),
.B1(n_81),
.B2(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_143),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_187),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_193),
.B(n_153),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_121),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_126),
.A3(n_138),
.B1(n_123),
.B2(n_99),
.C1(n_146),
.C2(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_150),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_116),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_189),
.B(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_140),
.B(n_27),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_12),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_2),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_12),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_178),
.B(n_155),
.C(n_176),
.D(n_153),
.Y(n_210)
);

BUFx12f_ASAP7_75t_SL g199 ( 
.A(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_209),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_156),
.B(n_157),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_213),
.B1(n_171),
.B2(n_198),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_167),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_212),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_175),
.B(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_160),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_215),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_198),
.C(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_222),
.C(n_226),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_154),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_181),
.C(n_158),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_158),
.C(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_230),
.B(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_200),
.B1(n_204),
.B2(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_222),
.C(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_242),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_226),
.B1(n_211),
.B2(n_210),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_208),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_229),
.B1(n_232),
.B2(n_230),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_246),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_203),
.B(n_231),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_185),
.B(n_165),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_208),
.A3(n_201),
.B1(n_221),
.B2(n_185),
.C1(n_165),
.C2(n_11),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_238),
.C(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_248),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_247),
.C(n_255),
.Y(n_258)
);

AOI321xp33_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_259),
.A3(n_249),
.B1(n_11),
.B2(n_9),
.C(n_5),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_2),
.Y(n_261)
);


endmodule