module real_jpeg_24415_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_16;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_3),
.A2(n_29),
.B1(n_38),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_15),
.B1(n_19),
.B2(n_46),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_20),
.B1(n_29),
.B2(n_38),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_6),
.A2(n_15),
.B1(n_19),
.B2(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_15),
.C(n_32),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_7),
.A2(n_29),
.B1(n_38),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_7),
.A2(n_14),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_68),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_47),
.B(n_67),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_26),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_12),
.B(n_26),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_24),
.B(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_15),
.A2(n_19),
.B1(n_32),
.B2(n_39),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_18),
.A2(n_51),
.B(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_28),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_29),
.A2(n_38),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_41),
.B(n_43),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_36),
.B(n_45),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_40),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_56),
.B(n_66),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_50),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_84),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);


endmodule