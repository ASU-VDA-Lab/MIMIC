module fake_jpeg_30971_n_436 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_436);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_436;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_79),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_47),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g82 ( 
.A(n_50),
.Y(n_82)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_60),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_57),
.Y(n_113)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_73),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_17),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_91),
.B1(n_54),
.B2(n_43),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_37),
.B(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_88),
.B(n_17),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_50),
.B(n_40),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

NAND2x1p5_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_59),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_77),
.B1(n_57),
.B2(n_67),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_40),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_48),
.A2(n_39),
.B(n_2),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_80),
.B(n_2),
.Y(n_131)
);

HAxp5_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_21),
.CON(n_126),
.SN(n_126)
);

BUFx12f_ASAP7_75t_SL g155 ( 
.A(n_126),
.Y(n_155)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_139),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_144),
.B(n_151),
.Y(n_178)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_63),
.B1(n_69),
.B2(n_68),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_146),
.B1(n_148),
.B2(n_156),
.Y(n_172)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_20),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_24),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_24),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_149),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_1),
.B(n_2),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_65),
.B1(n_62),
.B2(n_53),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_86),
.B1(n_93),
.B2(n_110),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_57),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_24),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_24),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_16),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_158),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_86),
.A2(n_103),
.B1(n_99),
.B2(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_84),
.B(n_16),
.Y(n_158)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_160),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_103),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_90),
.B1(n_121),
.B2(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_84),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_143),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_180),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_130),
.B1(n_121),
.B2(n_90),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_189),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_98),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_206),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_155),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_127),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_207),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_201),
.B1(n_215),
.B2(n_204),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_131),
.B1(n_144),
.B2(n_172),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_151),
.B(n_147),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_208),
.B(n_214),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_139),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_165),
.B(n_127),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_139),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_213),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_169),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_158),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_139),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_146),
.B1(n_139),
.B2(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_224),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_230),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_236),
.B1(n_199),
.B2(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_171),
.B1(n_177),
.B2(n_152),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_149),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_159),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_128),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_159),
.C(n_150),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_193),
.C(n_206),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_156),
.B1(n_161),
.B2(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_179),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_174),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_208),
.B(n_205),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_247),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_208),
.B(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_252),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_245),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_199),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_232),
.B1(n_219),
.B2(n_234),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_200),
.B1(n_213),
.B2(n_202),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_202),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_194),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_251),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_211),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_207),
.B(n_180),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_257),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_254),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_258),
.Y(n_270)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_174),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_128),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_229),
.B1(n_236),
.B2(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_235),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_275),
.C(n_281),
.Y(n_310)
);

XOR2x2_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_232),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_263),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_224),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_279),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_232),
.B(n_234),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_253),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_232),
.C(n_225),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_228),
.C(n_150),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_228),
.B1(n_188),
.B2(n_190),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_256),
.B1(n_248),
.B2(n_254),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_244),
.A2(n_188),
.B1(n_190),
.B2(n_210),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_290),
.B1(n_182),
.B2(n_168),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_287),
.C(n_246),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_195),
.C(n_176),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_247),
.A2(n_190),
.B1(n_210),
.B2(n_157),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_259),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_258),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_313),
.Y(n_329)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_241),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_307),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_300),
.B1(n_303),
.B2(n_317),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_276),
.B1(n_285),
.B2(n_280),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_248),
.B1(n_250),
.B2(n_254),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_245),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_311),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_272),
.A2(n_246),
.B1(n_257),
.B2(n_251),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_268),
.A2(n_238),
.B(n_243),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_292),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_195),
.Y(n_306)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_238),
.Y(n_308)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_182),
.Y(n_309)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_245),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_182),
.C(n_184),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_319),
.C(n_288),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_264),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_281),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_278),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_276),
.A2(n_110),
.B1(n_118),
.B2(n_122),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_289),
.A2(n_277),
.B1(n_267),
.B2(n_282),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_318),
.A2(n_290),
.B1(n_304),
.B2(n_277),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_186),
.C(n_176),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_293),
.B1(n_292),
.B2(n_274),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_327),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_332),
.Y(n_357)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_283),
.C(n_293),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_330),
.C(n_339),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_313),
.C(n_314),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_294),
.B(n_278),
.CI(n_283),
.CON(n_333),
.SN(n_333)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_287),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_334),
.B(n_336),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_135),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_264),
.Y(n_336)
);

FAx1_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_267),
.CI(n_168),
.CON(n_338),
.SN(n_338)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_338),
.A2(n_315),
.B(n_137),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_175),
.C(n_166),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_95),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_341),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_97),
.Y(n_342)
);

BUFx12_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_175),
.B1(n_166),
.B2(n_164),
.Y(n_347)
);

AO221x1_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_312),
.B1(n_295),
.B2(n_317),
.C(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_345),
.Y(n_373)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_321),
.B(n_339),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_355),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_337),
.A2(n_160),
.B1(n_118),
.B2(n_122),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_353),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_117),
.B1(n_116),
.B2(n_164),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_337),
.A2(n_133),
.B(n_107),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_354),
.A2(n_365),
.B(n_89),
.Y(n_381)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_160),
.B1(n_112),
.B2(n_117),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_116),
.B1(n_97),
.B2(n_112),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_364),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_93),
.B1(n_100),
.B2(n_133),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_363),
.B(n_136),
.Y(n_376)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_137),
.B(n_85),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_333),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_330),
.C(n_329),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_367),
.A2(n_374),
.B(n_357),
.Y(n_389)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_369),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_366),
.A2(n_338),
.B1(n_329),
.B2(n_324),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_370),
.A2(n_378),
.B1(n_365),
.B2(n_348),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_360),
.B(n_346),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_328),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_379),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_324),
.C(n_145),
.Y(n_374)
);

NOR2x1_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_140),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_376),
.A2(n_381),
.B1(n_375),
.B2(n_380),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_107),
.B1(n_101),
.B2(n_85),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_120),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_358),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_392),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_349),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_377),
.C(n_383),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_390),
.B(n_381),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_357),
.B(n_361),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_349),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_391),
.B(n_393),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_364),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_352),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_382),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_393),
.Y(n_404)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_400),
.B(n_406),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_401),
.B(n_405),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_106),
.C(n_89),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_378),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_404),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_383),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_387),
.B(n_356),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_358),
.B(n_377),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g410 ( 
.A1(n_407),
.A2(n_395),
.A3(n_391),
.B1(n_101),
.B2(n_113),
.C1(n_136),
.C2(n_124),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_385),
.A2(n_354),
.B1(n_358),
.B2(n_120),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

AOI21x1_ASAP7_75t_L g420 ( 
.A1(n_410),
.A2(n_15),
.B(n_3),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_106),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_412),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_399),
.A2(n_89),
.B(n_113),
.Y(n_413)
);

A2O1A1O1Ixp25_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_397),
.B(n_399),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_416),
.B(n_418),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g428 ( 
.A1(n_420),
.A2(n_423),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_428)
);

AOI21xp33_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_1),
.B(n_3),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g429 ( 
.A1(n_422),
.A2(n_425),
.B(n_8),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_414),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_5),
.C(n_6),
.Y(n_427)
);

A2O1A1O1Ixp25_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_417),
.B(n_409),
.C(n_415),
.D(n_7),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_4),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_427),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_428),
.Y(n_432)
);

OAI311xp33_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_419),
.A3(n_9),
.B1(n_10),
.C1(n_11),
.Y(n_430)
);

AOI322xp5_ASAP7_75t_L g433 ( 
.A1(n_430),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_433),
.Y(n_434)
);

OAI31xp33_ASAP7_75t_L g435 ( 
.A1(n_434),
.A2(n_431),
.A3(n_432),
.B(n_12),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_12),
.C(n_13),
.Y(n_436)
);


endmodule