module real_jpeg_23805_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_286;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_293;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_0),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_160)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_66),
.B1(n_74),
.B2(n_111),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_66),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_66),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_3),
.B(n_82),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_44),
.C(n_58),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_155),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_184),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_3),
.B(n_28),
.C(n_49),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_3),
.A2(n_30),
.B(n_245),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_72),
.B1(n_74),
.B2(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_6),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_136),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_136),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_136),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_8),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_71),
.Y(n_244)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_12),
.A2(n_72),
.B1(n_74),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_12),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_86),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_86),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_14),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_15),
.A2(n_29),
.B1(n_43),
.B2(n_44),
.Y(n_95)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_20),
.B(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_116),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.C(n_68),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_23),
.A2(n_24),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_25),
.A2(n_39),
.B1(n_40),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_25),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_26),
.A2(n_30),
.B1(n_102),
.B2(n_125),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_28),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_27),
.B(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_30),
.A2(n_34),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_30),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_30),
.A2(n_160),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_30),
.B(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_30),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_38),
.B(n_184),
.Y(n_270)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_42),
.A2(n_51),
.B1(n_93),
.B2(n_128),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_44),
.B(n_252),
.Y(n_251)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_47),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_47),
.A2(n_54),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_51),
.A2(n_128),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_51),
.A2(n_180),
.B(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_51),
.B(n_184),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_54),
.B(n_181),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_55),
.B(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_67),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_57),
.B1(n_67),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_56),
.A2(n_152),
.B(n_154),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_56),
.A2(n_154),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_65),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_57),
.A2(n_131),
.B(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_62),
.B1(n_79),
.B2(n_80),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_61),
.A2(n_72),
.A3(n_80),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_62),
.B(n_79),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_62),
.B(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_76),
.B(n_83),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_70),
.A2(n_77),
.B1(n_82),
.B2(n_135),
.Y(n_134)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_77),
.A2(n_84),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_110),
.B(n_114),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_81),
.A2(n_114),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_97),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_93),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_93),
.A2(n_233),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_121)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_103),
.B(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_111),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.C(n_134),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_124),
.B(n_127),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_153),
.B1(n_155),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_169),
.B(n_294),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_167),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_141),
.B(n_167),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_148),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_146),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_148),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_156),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_151),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_158),
.A2(n_256),
.B1(n_258),
.B2(n_260),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_201),
.B(n_288),
.C(n_293),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_195),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.C(n_187),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_172),
.A2(n_173),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_186),
.B(n_187),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_192),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_194),
.A2(n_257),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_196),
.B(n_199),
.C(n_200),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_282),
.B(n_287),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_234),
.B(n_281),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_223),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_206),
.B(n_223),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_216),
.C(n_220),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_210),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B(n_214),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_216),
.A2(n_220),
.B1(n_221),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_230),
.C(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_275),
.B(n_280),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_253),
.B(n_274),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_247),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_247),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_244),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_263),
.B(n_273),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_261),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_268),
.B(n_272),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);


endmodule