module fake_jpeg_3053_n_389 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_59),
.Y(n_115)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2x1p5_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_8),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_60),
.B(n_15),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_90),
.Y(n_119)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_88),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx2_ASAP7_75t_R g74 ( 
.A(n_27),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_39),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_43),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_85),
.Y(n_170)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_18),
.B(n_9),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_5),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_92),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_42),
.B(n_7),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_7),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx16f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_11),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_105),
.Y(n_127)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx12f_ASAP7_75t_SL g101 ( 
.A(n_27),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_106),
.B(n_110),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_53),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_13),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_13),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_111),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_49),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_60),
.A2(n_109),
.B(n_38),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_113),
.A2(n_127),
.B(n_120),
.C(n_118),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_48),
.C(n_51),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_121),
.B(n_156),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_131),
.B(n_153),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_52),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_133),
.B(n_163),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_67),
.A2(n_19),
.B1(n_50),
.B2(n_23),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_137),
.A2(n_62),
.B1(n_81),
.B2(n_93),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_55),
.B(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_141),
.B(n_147),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_66),
.A2(n_28),
.B1(n_47),
.B2(n_52),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_142),
.A2(n_144),
.B1(n_150),
.B2(n_114),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_57),
.A2(n_68),
.B1(n_84),
.B2(n_65),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_23),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_94),
.A2(n_47),
.B1(n_49),
.B2(n_37),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_95),
.A2(n_36),
.B1(n_37),
.B2(n_19),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_32),
.C(n_17),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_32),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_76),
.C(n_80),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_106),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_86),
.B(n_17),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_97),
.Y(n_176)
);

OR2x2_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_81),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_22),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_176),
.B(n_181),
.Y(n_267)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_177),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_72),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_178),
.B(n_212),
.Y(n_249)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_73),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_119),
.B(n_87),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_184),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_79),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_186),
.B(n_189),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_79),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_192),
.Y(n_232)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_188),
.Y(n_265)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_115),
.B(n_22),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_15),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_205),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_75),
.B1(n_64),
.B2(n_58),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_155),
.B1(n_158),
.B2(n_157),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_208),
.Y(n_230)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_128),
.B(n_138),
.C(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_204),
.B(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_41),
.B1(n_2),
.B2(n_1),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_41),
.B1(n_1),
.B2(n_15),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_167),
.A2(n_1),
.B1(n_114),
.B2(n_169),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_145),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_146),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_140),
.B(n_145),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_225),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_216),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_125),
.B(n_140),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_223),
.Y(n_257)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_175),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_222),
.Y(n_256)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_130),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_154),
.B(n_166),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_116),
.B(n_172),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_227),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_122),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_142),
.A2(n_150),
.B1(n_144),
.B2(n_148),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_229),
.Y(n_258)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_122),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_154),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_166),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_237),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_172),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_129),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_254),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_178),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_173),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_194),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_173),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_259),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_196),
.A2(n_129),
.B1(n_158),
.B2(n_197),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_185),
.B(n_180),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_177),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_204),
.B(n_186),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_189),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_272),
.B(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_235),
.B(n_225),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_251),
.B(n_255),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_277),
.A2(n_290),
.B(n_231),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_228),
.B1(n_224),
.B2(n_202),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_285),
.B1(n_295),
.B2(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_234),
.B(n_202),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_294),
.Y(n_306)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_280),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_245),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_286),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_234),
.A2(n_228),
.B1(n_224),
.B2(n_207),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_292),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_258),
.A2(n_224),
.B(n_228),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

CKINVDCx12_ASAP7_75t_R g293 ( 
.A(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_190),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_258),
.A2(n_208),
.B1(n_199),
.B2(n_182),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_201),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_259),
.C(n_260),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_247),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_236),
.A2(n_216),
.B1(n_221),
.B2(n_218),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_179),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_230),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_300),
.B1(n_282),
.B2(n_291),
.C(n_296),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_268),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_294),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_277),
.A2(n_250),
.B(n_253),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_305),
.A2(n_292),
.B(n_281),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_243),
.B1(n_254),
.B2(n_237),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_307),
.A2(n_315),
.B1(n_319),
.B2(n_301),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_313),
.B(n_270),
.Y(n_329)
);

NAND2x1_ASAP7_75t_SL g313 ( 
.A(n_278),
.B(n_230),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_276),
.A2(n_230),
.B1(n_259),
.B2(n_257),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.C(n_275),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_232),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_275),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_271),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_285),
.A2(n_299),
.B1(n_295),
.B2(n_271),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_314),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_330),
.Y(n_353)
);

OAI22x1_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_287),
.B1(n_286),
.B2(n_284),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_328),
.B1(n_307),
.B2(n_304),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_326),
.B(n_327),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_332),
.B(n_333),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_241),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_273),
.C(n_244),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_334),
.C(n_335),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_310),
.A2(n_289),
.B(n_299),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_248),
.C(n_298),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_248),
.C(n_239),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_320),
.B(n_239),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_306),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_305),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_264),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_313),
.B(n_312),
.Y(n_342)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_340),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_347),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_342),
.A2(n_344),
.B(n_339),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_312),
.B(n_314),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_348),
.A2(n_328),
.B1(n_304),
.B2(n_339),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_306),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_354),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_314),
.C(n_315),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_351),
.B(n_321),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_355),
.B(n_358),
.Y(n_367)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_345),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_361),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_309),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_359),
.A2(n_363),
.B1(n_364),
.B2(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_338),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_362),
.Y(n_370)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_350),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_322),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_366),
.A2(n_369),
.B1(n_371),
.B2(n_372),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_359),
.A2(n_348),
.B1(n_343),
.B2(n_325),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_363),
.A2(n_341),
.B1(n_354),
.B2(n_334),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_364),
.A2(n_360),
.B1(n_349),
.B2(n_347),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_365),
.A2(n_346),
.B(n_311),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_373),
.A2(n_346),
.B(n_356),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_372),
.B(n_365),
.C(n_349),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_374),
.B(n_379),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_370),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_L g377 ( 
.A1(n_366),
.A2(n_322),
.A3(n_356),
.B1(n_308),
.B2(n_331),
.C1(n_311),
.C2(n_326),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_367),
.A2(n_308),
.B(n_264),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_266),
.C(n_265),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_269),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_371),
.C(n_369),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_381),
.B(n_377),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_252),
.C(n_203),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

AOI322xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_280),
.A3(n_193),
.B1(n_382),
.B2(n_380),
.C1(n_229),
.C2(n_188),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_387),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_388),
.Y(n_389)
);


endmodule