module fake_jpeg_31878_n_438 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_438);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_43),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_56),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_68),
.Y(n_118)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_9),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_92),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_122),
.B1(n_30),
.B2(n_32),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_43),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_58),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_44),
.B(n_40),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_113),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_39),
.B1(n_28),
.B2(n_29),
.Y(n_122)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_30),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_148),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_144),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_73),
.B1(n_49),
.B2(n_45),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_138),
.B(n_146),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_51),
.B1(n_76),
.B2(n_52),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_147),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_79),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_31),
.B(n_40),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_48),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_32),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_152),
.Y(n_188)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_42),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_25),
.B1(n_36),
.B2(n_39),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_71),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_162),
.B(n_100),
.Y(n_173)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_25),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_160),
.Y(n_192)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_105),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_163),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_42),
.B(n_36),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_86),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_112),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_185),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_100),
.B(n_106),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_147),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_152),
.B1(n_149),
.B2(n_131),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_183),
.B1(n_135),
.B2(n_93),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_161),
.B1(n_159),
.B2(n_94),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_140),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_157),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_155),
.B1(n_147),
.B2(n_137),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_194),
.A2(n_201),
.B1(n_218),
.B2(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_137),
.C(n_140),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_196),
.B(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_176),
.B(n_173),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_155),
.B1(n_138),
.B2(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g231 ( 
.A(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_158),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_85),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_210),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_188),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_169),
.A2(n_135),
.B1(n_136),
.B2(n_129),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_172),
.B1(n_175),
.B2(n_178),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_144),
.B(n_154),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_133),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_175),
.B1(n_178),
.B2(n_169),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_219),
.A2(n_226),
.B1(n_164),
.B2(n_160),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_233),
.B(n_200),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_207),
.B(n_194),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_188),
.B1(n_182),
.B2(n_172),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_182),
.A3(n_185),
.B1(n_125),
.B2(n_115),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_232),
.A2(n_230),
.B1(n_220),
.B2(n_241),
.Y(n_268)
);

AO22x1_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_160),
.B1(n_166),
.B2(n_190),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_214),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_186),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

NAND2x1p5_ASAP7_75t_R g293 ( 
.A(n_248),
.B(n_253),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_186),
.B(n_168),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_218),
.B1(n_207),
.B2(n_215),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_254),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_240),
.B1(n_219),
.B2(n_221),
.Y(n_254)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_257),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_201),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_190),
.Y(n_276)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_195),
.B(n_197),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_262),
.Y(n_280)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_260),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_217),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_213),
.B1(n_204),
.B2(n_205),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_268),
.B1(n_229),
.B2(n_222),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_266),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_143),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_171),
.B(n_189),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_171),
.B1(n_166),
.B2(n_89),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_231),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_296),
.B1(n_265),
.B2(n_266),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_229),
.C(n_222),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_277),
.C(n_287),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_112),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_170),
.C(n_189),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_285),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_170),
.Y(n_286)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_168),
.C(n_165),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_245),
.A2(n_231),
.B1(n_235),
.B2(n_198),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_250),
.B1(n_242),
.B2(n_258),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_165),
.C(n_134),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_291),
.C(n_129),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_163),
.C(n_156),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_245),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_106),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_143),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_242),
.A2(n_231),
.B1(n_235),
.B2(n_198),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_296),
.B1(n_294),
.B2(n_281),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_302),
.A2(n_316),
.B1(n_307),
.B2(n_300),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_264),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_322),
.C(n_287),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_248),
.B(n_257),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_306),
.A2(n_139),
.B(n_142),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_308),
.B(n_142),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_272),
.B(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_313),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_255),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_321),
.Y(n_332)
);

AO22x1_ASAP7_75t_SL g315 ( 
.A1(n_269),
.A2(n_97),
.B1(n_89),
.B2(n_126),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_318),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_116),
.B1(n_97),
.B2(n_126),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_283),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_290),
.B(n_16),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_320),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_123),
.C(n_121),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_324),
.A2(n_329),
.B1(n_339),
.B2(n_136),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_68),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_275),
.C(n_289),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_291),
.C(n_280),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_269),
.C(n_295),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_301),
.A2(n_314),
.B1(n_305),
.B2(n_319),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_283),
.C(n_271),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_342),
.C(n_343),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_335),
.B(n_344),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_337),
.Y(n_369)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_278),
.B1(n_116),
.B2(n_108),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_108),
.B1(n_119),
.B2(n_105),
.Y(n_341)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_125),
.C(n_119),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_50),
.C(n_54),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_310),
.B(n_323),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_345),
.B(n_14),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_316),
.A2(n_94),
.B1(n_25),
.B2(n_95),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

OAI321xp33_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_311),
.A3(n_303),
.B1(n_309),
.B2(n_315),
.C(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_315),
.B1(n_120),
.B2(n_59),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_351),
.A2(n_69),
.B1(n_7),
.B2(n_10),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_327),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_363),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_142),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_359),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_139),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_326),
.A2(n_14),
.B(n_16),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_366),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_334),
.A2(n_139),
.B(n_13),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_37),
.Y(n_385)
);

AOI21xp33_ASAP7_75t_L g365 ( 
.A1(n_333),
.A2(n_11),
.B(n_15),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_365),
.Y(n_384)
);

BUFx12f_ASAP7_75t_SL g367 ( 
.A(n_342),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_7),
.Y(n_380)
);

BUFx12_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_335),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_358),
.A2(n_324),
.B1(n_325),
.B2(n_330),
.Y(n_372)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_376),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_353),
.A2(n_328),
.B(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_374),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_47),
.C(n_46),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_120),
.C(n_10),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_379),
.Y(n_396)
);

XOR2x2_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_357),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_378),
.B(n_380),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_6),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_10),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_369),
.B1(n_356),
.B2(n_380),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_360),
.C(n_348),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_390),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_361),
.C(n_364),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_363),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_349),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_397),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_386),
.A2(n_361),
.B(n_366),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_12),
.B(n_11),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_368),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_398),
.B(n_399),
.Y(n_400)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_387),
.A2(n_372),
.B1(n_368),
.B2(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_405),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_391),
.A2(n_381),
.B(n_375),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_407),
.B(n_408),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_388),
.A2(n_36),
.B(n_6),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_393),
.C(n_399),
.Y(n_408)
);

OAI21x1_ASAP7_75t_SL g409 ( 
.A1(n_393),
.A2(n_6),
.B(n_15),
.Y(n_409)
);

AOI221xp5_ASAP7_75t_L g417 ( 
.A1(n_409),
.A2(n_410),
.B1(n_0),
.B2(n_1),
.C(n_2),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_396),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_0),
.Y(n_415)
);

NAND4xp25_ASAP7_75t_SL g414 ( 
.A(n_400),
.B(n_12),
.C(n_11),
.D(n_37),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_420),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_403),
.A2(n_36),
.B(n_1),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_416),
.A2(n_418),
.B(n_4),
.Y(n_426)
);

OAI21x1_ASAP7_75t_SL g424 ( 
.A1(n_417),
.A2(n_4),
.B(n_5),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_404),
.B(n_1),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_419),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_36),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_SL g422 ( 
.A(n_421),
.B(n_3),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_426),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_428),
.A2(n_420),
.B1(n_37),
.B2(n_5),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_412),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_431),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_432),
.B(n_427),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_430),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_433),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_SL g437 ( 
.A1(n_436),
.A2(n_423),
.B(n_429),
.C(n_37),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_4),
.Y(n_438)
);


endmodule