module fake_jpeg_1670_n_500 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_500);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_500;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_9),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_54),
.Y(n_108)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_15),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_66),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_89),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_24),
.Y(n_114)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_40),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_40),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_90),
.B(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_40),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_96),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_99),
.Y(n_115)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_109),
.B(n_124),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_114),
.B(n_28),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_51),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_32),
.C(n_20),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_149),
.Y(n_196)
);

BUFx16f_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

CKINVDCx6p67_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_22),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_133),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_38),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_38),
.B1(n_23),
.B2(n_48),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_134),
.A2(n_145),
.B1(n_19),
.B2(n_47),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_81),
.A2(n_41),
.B1(n_24),
.B2(n_34),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_65),
.A2(n_23),
.B1(n_32),
.B2(n_20),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_56),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_79),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_71),
.B(n_48),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_158),
.Y(n_187)
);

BUFx16f_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_91),
.B(n_48),
.Y(n_158)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_160),
.Y(n_242)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_103),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_163),
.B(n_183),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_165),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_101),
.A2(n_75),
.B1(n_78),
.B2(n_77),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_166),
.A2(n_167),
.B1(n_175),
.B2(n_179),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_41),
.B1(n_37),
.B2(n_45),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_112),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_194),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_117),
.A2(n_41),
.B1(n_24),
.B2(n_18),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_108),
.B(n_32),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_181),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_25),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_126),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_30),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_197),
.Y(n_227)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_131),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_190),
.B(n_204),
.Y(n_251)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_201),
.Y(n_231)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_130),
.B(n_60),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_209),
.B(n_47),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx12_ASAP7_75t_R g202 ( 
.A(n_106),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_203),
.Y(n_233)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_205),
.B(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_207),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_211),
.Y(n_255)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_138),
.B(n_59),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_19),
.B1(n_100),
.B2(n_140),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_114),
.B(n_30),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_213),
.Y(n_262)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_122),
.B(n_30),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_110),
.B(n_28),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_47),
.B1(n_19),
.B2(n_73),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_76),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_218),
.B(n_239),
.C(n_247),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_46),
.B1(n_28),
.B2(n_157),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_222),
.A2(n_246),
.B1(n_252),
.B2(n_143),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_145),
.B(n_98),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_226),
.A2(n_172),
.B(n_170),
.Y(n_279)
);

BUFx2_ASAP7_75t_SL g266 ( 
.A(n_235),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_168),
.B(n_171),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_200),
.B1(n_195),
.B2(n_193),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_142),
.Y(n_239)
);

AO22x1_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_94),
.B1(n_95),
.B2(n_140),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_143),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_207),
.B1(n_203),
.B2(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_175),
.B(n_185),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_82),
.C(n_86),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_256),
.C(n_257),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_198),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_173),
.B(n_68),
.C(n_84),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_169),
.B(n_87),
.C(n_151),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_177),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_209),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_218),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_271),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_168),
.B(n_166),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_270),
.B1(n_285),
.B2(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_281),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_245),
.A2(n_177),
.B1(n_174),
.B2(n_178),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_274),
.Y(n_334)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_278),
.Y(n_330)
);

OR2x2_ASAP7_75t_SL g339 ( 
.A(n_276),
.B(n_164),
.Y(n_339)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_279),
.A2(n_296),
.B(n_233),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_248),
.B(n_168),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_280),
.B(n_282),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_238),
.B(n_182),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_220),
.B(n_182),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_286),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_160),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_221),
.B(n_227),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_294),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_238),
.B(n_120),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_291),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_231),
.B(n_120),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_121),
.B1(n_119),
.B2(n_157),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_253),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_295),
.Y(n_326)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_236),
.A2(n_164),
.B(n_165),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_142),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_219),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_302),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_228),
.B(n_15),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_251),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_301),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_17),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_262),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_230),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_263),
.A2(n_234),
.B1(n_226),
.B2(n_240),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_325),
.B1(n_119),
.B2(n_116),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_259),
.C(n_258),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_316),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_313),
.A2(n_339),
.B(n_281),
.Y(n_347)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_250),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_314),
.B(n_304),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_256),
.C(n_257),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_291),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_328),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_263),
.A2(n_240),
.B1(n_252),
.B2(n_254),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_327),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_224),
.C(n_253),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_320),
.B(n_324),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_264),
.A2(n_242),
.B1(n_260),
.B2(n_232),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_332),
.B1(n_230),
.B2(n_303),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_224),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_268),
.A2(n_242),
.B1(n_249),
.B2(n_116),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_264),
.A2(n_268),
.B1(n_292),
.B2(n_289),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_249),
.C(n_225),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_331),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_268),
.A2(n_225),
.B1(n_121),
.B2(n_151),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_281),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_268),
.Y(n_356)
);

BUFx8_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVx13_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

NOR4xp25_ASAP7_75t_SL g340 ( 
.A(n_338),
.B(n_339),
.C(n_306),
.D(n_313),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_306),
.A2(n_298),
.A3(n_295),
.B1(n_265),
.B2(n_293),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_366),
.Y(n_377)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_338),
.A2(n_279),
.B(n_302),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_343),
.A2(n_346),
.B(n_347),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_307),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_329),
.A2(n_271),
.B(n_300),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_266),
.B(n_293),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_317),
.Y(n_353)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_326),
.A2(n_272),
.B(n_274),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_356),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_270),
.Y(n_357)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_308),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_369),
.Y(n_394)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_360),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_305),
.B(n_275),
.Y(n_364)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_330),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_326),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_368),
.B1(n_319),
.B2(n_332),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_309),
.A2(n_278),
.B1(n_294),
.B2(n_277),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_315),
.B(n_282),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_370),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_371),
.A2(n_322),
.B1(n_321),
.B2(n_335),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_372),
.A2(n_355),
.B1(n_368),
.B2(n_363),
.Y(n_407)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_315),
.B1(n_335),
.B2(n_310),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_376),
.A2(n_363),
.B1(n_367),
.B2(n_365),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_320),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_395),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_328),
.C(n_316),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_391),
.C(n_399),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_312),
.C(n_324),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_346),
.Y(n_393)
);

NOR3xp33_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_34),
.C(n_164),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_314),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_336),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_398),
.C(n_370),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_333),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_331),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_357),
.C(n_366),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_406),
.C(n_410),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_388),
.A2(n_355),
.B1(n_361),
.B2(n_377),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_407),
.B1(n_413),
.B2(n_418),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_343),
.B(n_350),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_405),
.A2(n_421),
.B(n_387),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_357),
.C(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_394),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_347),
.C(n_364),
.Y(n_410)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

XOR2x2_ASAP7_75t_SL g412 ( 
.A(n_377),
.B(n_340),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_389),
.Y(n_437)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_414),
.A2(n_404),
.B1(n_388),
.B2(n_405),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_362),
.C(n_342),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_400),
.C(n_396),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_353),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_422),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_369),
.B1(n_334),
.B2(n_359),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_380),
.B(n_359),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_384),
.Y(n_432)
);

INVx13_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_420),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_376),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_360),
.B1(n_34),
.B2(n_85),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_423),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_425),
.A2(n_433),
.B1(n_437),
.B2(n_441),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_432),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_396),
.C(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_417),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_414),
.A2(n_384),
.B1(n_390),
.B2(n_392),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_389),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_437),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_387),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_31),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_374),
.Y(n_441)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_441),
.Y(n_448)
);

OAI321xp33_ASAP7_75t_L g450 ( 
.A1(n_442),
.A2(n_419),
.A3(n_420),
.B1(n_373),
.B2(n_165),
.C(n_13),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_440),
.Y(n_443)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_417),
.C(n_415),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_446),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_438),
.A2(n_421),
.B1(n_412),
.B2(n_403),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_374),
.B1(n_406),
.B2(n_375),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_452),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_426),
.B(n_432),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_26),
.C(n_31),
.Y(n_452)
);

BUFx12_ASAP7_75t_L g453 ( 
.A(n_439),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_455),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_456),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_26),
.C(n_31),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_26),
.C(n_31),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_425),
.C(n_433),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_442),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_464),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_460),
.A2(n_453),
.B(n_452),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_465),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_445),
.B(n_431),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_429),
.C(n_427),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_429),
.C(n_435),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_468),
.C(n_14),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_439),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_448),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_476),
.Y(n_481)
);

NAND2x1_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_13),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_463),
.A2(n_453),
.B1(n_457),
.B2(n_8),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_473),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_31),
.C(n_17),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_17),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_478),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_14),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_479),
.B(n_480),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_9),
.Y(n_480)
);

AOI21xp33_ASAP7_75t_L g483 ( 
.A1(n_474),
.A2(n_469),
.B(n_463),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_484),
.B(n_485),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_461),
.C(n_470),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_487),
.B(n_0),
.C(n_1),
.Y(n_491)
);

AOI322xp5_ASAP7_75t_L g488 ( 
.A1(n_481),
.A2(n_473),
.A3(n_485),
.B1(n_486),
.B2(n_484),
.C1(n_476),
.C2(n_482),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_489),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_482),
.A2(n_480),
.B(n_1),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_4),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_492),
.B(n_4),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_494),
.B(n_495),
.C(n_490),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_493),
.Y(n_495)
);

AOI322xp5_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_487),
.C1(n_493),
.C2(n_453),
.Y(n_497)
);

MAJx2_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_5),
.C(n_6),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_5),
.B(n_6),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_7),
.Y(n_500)
);


endmodule