module fake_netlist_5_1610_n_8442 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_737, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_733, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_726, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_713, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_256, n_305, n_533, n_52, n_278, n_110, n_8442);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_733;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_713;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_8442;

wire n_924;
wire n_6643;
wire n_6122;
wire n_977;
wire n_2417;
wire n_2253;
wire n_2756;
wire n_7981;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_6579;
wire n_7164;
wire n_5287;
wire n_6546;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_8174;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_6786;
wire n_7206;
wire n_7303;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_8363;
wire n_2021;
wire n_7710;
wire n_8383;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_8328;
wire n_2059;
wire n_7461;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_6649;
wire n_8060;
wire n_7154;
wire n_3202;
wire n_8002;
wire n_4977;
wire n_3813;
wire n_6810;
wire n_7660;
wire n_6276;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_7686;
wire n_4211;
wire n_7024;
wire n_3448;
wire n_7205;
wire n_6742;
wire n_3019;
wire n_2096;
wire n_8319;
wire n_6694;
wire n_877;
wire n_3776;
wire n_7616;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_1696;
wire n_7486;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_8244;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_1107;
wire n_6090;
wire n_6580;
wire n_7010;
wire n_5480;
wire n_6549;
wire n_8105;
wire n_6913;
wire n_7867;
wire n_2147;
wire n_3010;
wire n_7315;
wire n_7004;
wire n_2770;
wire n_4131;
wire n_7772;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_7641;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_1242;
wire n_7468;
wire n_5469;
wire n_2323;
wire n_6431;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_7861;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_8413;
wire n_5202;
wire n_5648;
wire n_7667;
wire n_1314;
wire n_1512;
wire n_6931;
wire n_8114;
wire n_1490;
wire n_6618;
wire n_6408;
wire n_3214;
wire n_7523;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_8158;
wire n_1449;
wire n_6698;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_8104;
wire n_5848;
wire n_5406;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_7421;
wire n_7306;
wire n_6214;
wire n_7493;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_7804;
wire n_8089;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_6939;
wire n_882;
wire n_2384;
wire n_7528;
wire n_3156;
wire n_8262;
wire n_8290;
wire n_3376;
wire n_7562;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_6586;
wire n_2202;
wire n_2648;
wire n_8147;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_8310;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_6707;
wire n_2276;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_8380;
wire n_845;
wire n_7402;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_901;
wire n_4484;
wire n_7592;
wire n_3668;
wire n_7152;
wire n_6512;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_8126;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_7801;
wire n_7992;
wire n_1151;
wire n_1405;
wire n_7463;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_8305;
wire n_6725;
wire n_7613;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_6464;
wire n_2863;
wire n_2072;
wire n_8317;
wire n_2738;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_2968;
wire n_7316;
wire n_1585;
wire n_6820;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_6098;
wire n_7019;
wire n_6686;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_7956;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_7323;
wire n_2248;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_3007;
wire n_1000;
wire n_6769;
wire n_7683;
wire n_6592;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_6062;
wire n_6191;
wire n_7903;
wire n_2258;
wire n_748;
wire n_1667;
wire n_1058;
wire n_838;
wire n_8440;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_8416;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_8064;
wire n_5909;
wire n_1385;
wire n_7575;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_6043;
wire n_2987;
wire n_1527;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_7701;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_8214;
wire n_5055;
wire n_2175;
wire n_6793;
wire n_7873;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_7127;
wire n_5397;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_7568;
wire n_3208;
wire n_6021;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_5695;
wire n_7814;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_6926;
wire n_3649;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_7965;
wire n_2514;
wire n_6304;
wire n_5862;
wire n_8228;
wire n_8210;
wire n_5189;
wire n_6956;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_1027;
wire n_4160;
wire n_6782;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_7002;
wire n_8387;
wire n_1412;
wire n_3981;
wire n_8410;
wire n_7141;
wire n_5936;
wire n_6126;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_6027;
wire n_6598;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_870;
wire n_1711;
wire n_6638;
wire n_1891;
wire n_7308;
wire n_5254;
wire n_3526;
wire n_6900;
wire n_2546;
wire n_965;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_7457;
wire n_4613;
wire n_7718;
wire n_4649;
wire n_7617;
wire n_1888;
wire n_6269;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_7768;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_7974;
wire n_6013;
wire n_7357;
wire n_2449;
wire n_5083;
wire n_8247;
wire n_6927;
wire n_7975;
wire n_1194;
wire n_6503;
wire n_5888;
wire n_8172;
wire n_2297;
wire n_4186;
wire n_7310;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_7593;
wire n_6256;
wire n_7716;
wire n_2876;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_5870;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_7076;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_6982;
wire n_1680;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_7848;
wire n_6727;
wire n_3317;
wire n_8218;
wire n_7539;
wire n_1121;
wire n_7229;
wire n_4391;
wire n_949;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_8368;
wire n_4681;
wire n_8334;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_8159;
wire n_3455;
wire n_6097;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_1195;
wire n_7797;
wire n_4707;
wire n_2577;
wire n_8216;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_2796;
wire n_757;
wire n_7869;
wire n_6466;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_8337;
wire n_8257;
wire n_7983;
wire n_2805;
wire n_7781;
wire n_8125;
wire n_1145;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_1153;
wire n_741;
wire n_7624;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_1163;
wire n_8063;
wire n_6805;
wire n_6185;
wire n_5010;
wire n_1207;
wire n_7762;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_6568;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_8295;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_940;
wire n_6351;
wire n_7552;
wire n_8059;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_8146;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_6901;
wire n_8082;
wire n_2947;
wire n_978;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_6411;
wire n_3515;
wire n_8339;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_7746;
wire n_5435;
wire n_1431;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_8032;
wire n_7139;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4232;
wire n_4125;
wire n_8351;
wire n_4949;
wire n_2941;
wire n_8196;
wire n_6594;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_7857;
wire n_962;
wire n_2536;
wire n_6387;
wire n_1336;
wire n_7223;
wire n_1758;
wire n_7890;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_7964;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_6019;
wire n_6222;
wire n_7165;
wire n_8110;
wire n_3505;
wire n_6223;
wire n_4610;
wire n_6435;
wire n_3730;
wire n_4489;
wire n_7235;
wire n_974;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_5657;
wire n_957;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_6844;
wire n_3001;
wire n_7795;
wire n_7404;
wire n_3945;
wire n_4542;
wire n_2729;
wire n_2261;
wire n_6295;
wire n_3597;
wire n_8087;
wire n_8119;
wire n_1612;
wire n_7885;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_5857;
wire n_8173;
wire n_4534;
wire n_4500;
wire n_7437;
wire n_5014;
wire n_6241;
wire n_8420;
wire n_3185;
wire n_1300;
wire n_6087;
wire n_1127;
wire n_8019;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_6041;
wire n_7822;
wire n_2017;
wire n_2604;
wire n_6994;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_7329;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_6790;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_7194;
wire n_6273;
wire n_3474;
wire n_3984;
wire n_6807;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_8221;
wire n_1913;
wire n_7708;
wire n_1823;
wire n_7696;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_7115;
wire n_4189;
wire n_5670;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_7958;
wire n_8128;
wire n_4687;
wire n_948;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_6218;
wire n_7281;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_8106;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_6824;
wire n_1552;
wire n_6189;
wire n_3618;
wire n_2593;
wire n_8299;
wire n_5262;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_8287;
wire n_815;
wire n_4594;
wire n_6153;
wire n_7989;
wire n_3424;
wire n_5970;
wire n_1381;
wire n_6418;
wire n_1037;
wire n_6564;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_8197;
wire n_2786;
wire n_8081;
wire n_7192;
wire n_3171;
wire n_6671;
wire n_1437;
wire n_6591;
wire n_6266;
wire n_7161;
wire n_7580;
wire n_7153;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_6517;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_7350;
wire n_5690;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_6967;
wire n_5885;
wire n_2254;
wire n_6433;
wire n_1382;
wire n_3546;
wire n_925;
wire n_7535;
wire n_6893;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_4575;
wire n_3012;
wire n_7632;
wire n_8140;
wire n_3244;
wire n_6501;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_8137;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_6798;
wire n_5702;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_7844;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_4572;
wire n_3073;
wire n_1157;
wire n_8423;
wire n_5527;
wire n_6986;
wire n_802;
wire n_8090;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_6745;
wire n_8260;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_6209;
wire n_2263;
wire n_6875;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_7905;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_5551;
wire n_7594;
wire n_7766;
wire n_3715;
wire n_7803;
wire n_7340;
wire n_6699;
wire n_7747;
wire n_6073;
wire n_972;
wire n_8205;
wire n_5767;
wire n_8401;
wire n_6324;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_2499;
wire n_1200;
wire n_8284;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_6138;
wire n_7603;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_7726;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_8024;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_6477;
wire n_3734;
wire n_8133;
wire n_8373;
wire n_4778;
wire n_2429;
wire n_883;
wire n_6159;
wire n_6283;
wire n_7396;
wire n_5322;
wire n_856;
wire n_7116;
wire n_1793;
wire n_4352;
wire n_7519;
wire n_4441;
wire n_6943;
wire n_918;
wire n_4761;
wire n_6827;
wire n_6173;
wire n_8318;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_6312;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_7770;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1096;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_7664;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_6300;
wire n_7815;
wire n_2043;
wire n_2751;
wire n_8163;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_6537;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_7023;
wire n_1807;
wire n_2618;
wire n_7428;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_6783;
wire n_4748;
wire n_7465;
wire n_3931;
wire n_2295;
wire n_4010;
wire n_1219;
wire n_8293;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_7961;
wire n_1722;
wire n_7847;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_7149;
wire n_2795;
wire n_8252;
wire n_6459;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_7700;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_8367;
wire n_3538;
wire n_6869;
wire n_8078;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_7914;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_7967;
wire n_4728;
wire n_7117;
wire n_789;
wire n_4247;
wire n_4933;
wire n_6977;
wire n_4018;
wire n_3900;
wire n_7984;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_8361;
wire n_6313;
wire n_3872;
wire n_4336;
wire n_6569;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_6555;
wire n_3877;
wire n_6639;
wire n_7516;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3977;
wire n_3547;
wire n_1102;
wire n_7596;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_6490;
wire n_8301;
wire n_2633;
wire n_6961;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_5460;
wire n_7628;
wire n_4304;
wire n_6761;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_6294;
wire n_6767;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_4805;
wire n_4885;
wire n_7838;
wire n_8364;
wire n_7786;
wire n_5983;
wire n_1661;
wire n_5804;
wire n_7979;
wire n_6376;
wire n_3565;
wire n_6167;
wire n_7926;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_861;
wire n_6582;
wire n_1658;
wire n_7752;
wire n_1904;
wire n_6996;
wire n_1345;
wire n_1899;
wire n_6974;
wire n_7731;
wire n_6765;
wire n_7577;
wire n_8388;
wire n_8321;
wire n_1003;
wire n_6921;
wire n_2067;
wire n_8044;
wire n_8091;
wire n_2219;
wire n_7845;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_7709;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_6898;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_8261;
wire n_1657;
wire n_5886;
wire n_768;
wire n_7080;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_7744;
wire n_1491;
wire n_754;
wire n_8034;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_6960;
wire n_8201;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_1915;
wire n_5610;
wire n_1109;
wire n_5239;
wire n_6836;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_6972;
wire n_2924;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_5785;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_6093;
wire n_4538;
wire n_5994;
wire n_8093;
wire n_766;
wire n_6010;
wire n_7247;
wire n_8061;
wire n_1117;
wire n_6833;
wire n_2754;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_7481;
wire n_5204;
wire n_7292;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_7687;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_6265;
wire n_1650;
wire n_1137;
wire n_6821;
wire n_3934;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_5788;
wire n_8191;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_6676;
wire n_2372;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_8136;
wire n_2430;
wire n_7742;
wire n_2433;
wire n_3293;
wire n_7955;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_7758;
wire n_7547;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_6648;
wire n_7880;
wire n_4601;
wire n_8075;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_909;
wire n_5630;
wire n_1497;
wire n_8071;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_7513;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_1981;
wire n_7540;
wire n_1663;
wire n_1718;
wire n_4858;
wire n_4509;
wire n_3700;
wire n_5504;
wire n_7622;
wire n_7005;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_7353;
wire n_6219;
wire n_1889;
wire n_8315;
wire n_6965;
wire n_5025;
wire n_1489;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_8314;
wire n_6720;
wire n_1569;
wire n_8149;
wire n_2188;
wire n_6032;
wire n_7174;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_756;
wire n_1429;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_7607;
wire n_8209;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_7816;
wire n_3170;
wire n_7591;
wire n_5775;
wire n_8141;
wire n_2748;
wire n_3311;
wire n_7830;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_8302;
wire n_2898;
wire n_2717;
wire n_7151;
wire n_6229;
wire n_1861;
wire n_760;
wire n_5731;
wire n_5581;
wire n_3628;
wire n_3691;
wire n_6668;
wire n_7446;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_7053;
wire n_5831;
wire n_2573;
wire n_7473;
wire n_4435;
wire n_2939;
wire n_8070;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_886;
wire n_5653;
wire n_8248;
wire n_7966;
wire n_6258;
wire n_7070;
wire n_1221;
wire n_5394;
wire n_6755;
wire n_2774;
wire n_7276;
wire n_7351;
wire n_1707;
wire n_7942;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_6084;
wire n_4827;
wire n_8411;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_2488;
wire n_7666;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_7211;
wire n_4399;
wire n_6531;
wire n_2781;
wire n_5309;
wire n_7901;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_7368;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_6771;
wire n_2526;
wire n_6389;
wire n_2703;
wire n_8004;
wire n_2167;
wire n_8375;
wire n_5764;
wire n_5428;
wire n_6910;
wire n_6442;
wire n_3391;
wire n_6102;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_6441;
wire n_5543;
wire n_816;
wire n_5678;
wire n_5935;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_7677;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_871;
wire n_7929;
wire n_3738;
wire n_8399;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_4526;
wire n_2018;
wire n_3464;
wire n_6331;
wire n_1555;
wire n_6006;
wire n_8421;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_6278;
wire n_6787;
wire n_6872;
wire n_4899;
wire n_796;
wire n_6208;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_6632;
wire n_1012;
wire n_5411;
wire n_7754;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_8001;
wire n_5671;
wire n_3076;
wire n_8322;
wire n_6990;
wire n_8403;
wire n_3535;
wire n_2182;
wire n_6349;
wire n_3251;
wire n_1061;
wire n_2931;
wire n_7631;
wire n_6830;
wire n_5185;
wire n_7939;
wire n_7898;
wire n_1193;
wire n_6359;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_8313;
wire n_2146;
wire n_7763;
wire n_1487;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_781;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_6301;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_7945;
wire n_5945;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_6744;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_7381;
wire n_5565;
wire n_4081;
wire n_1103;
wire n_7948;
wire n_3132;
wire n_4407;
wire n_8102;
wire n_7291;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_7430;
wire n_3267;
wire n_4995;
wire n_7870;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_4446;
wire n_3373;
wire n_2279;
wire n_6104;
wire n_3884;
wire n_6475;
wire n_6465;
wire n_3726;
wire n_6496;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_8238;
wire n_6998;
wire n_6145;
wire n_3577;
wire n_2820;
wire n_7305;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_7980;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_7075;
wire n_7545;
wire n_7846;
wire n_1448;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_8438;
wire n_6194;
wire n_7695;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_8095;
wire n_7537;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_7489;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_8112;
wire n_1186;
wire n_5883;
wire n_6985;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_7451;
wire n_6238;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_6548;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_6366;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_7236;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_7269;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_3256;
wire n_7560;
wire n_7326;
wire n_7060;
wire n_2386;
wire n_1501;
wire n_7572;
wire n_3086;
wire n_1007;
wire n_6885;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_6529;
wire n_8169;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_8017;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_6423;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_7140;
wire n_7233;
wire n_819;
wire n_5088;
wire n_2302;
wire n_6558;
wire n_5457;
wire n_7352;
wire n_951;
wire n_7986;
wire n_7134;
wire n_5532;
wire n_1494;
wire n_2069;
wire n_6950;
wire n_7246;
wire n_6525;
wire n_7650;
wire n_3434;
wire n_1806;
wire n_933;
wire n_6631;
wire n_6892;
wire n_8203;
wire n_1563;
wire n_7663;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_2482;
wire n_2677;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_7729;
wire n_3987;
wire n_7339;
wire n_902;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_8138;
wire n_6658;
wire n_6264;
wire n_6925;
wire n_5919;
wire n_1698;
wire n_2329;
wire n_8206;
wire n_1098;
wire n_2142;
wire n_7767;
wire n_8190;
wire n_6176;
wire n_5410;
wire n_3332;
wire n_7146;
wire n_1135;
wire n_8092;
wire n_3048;
wire n_3937;
wire n_6124;
wire n_7672;
wire n_2203;
wire n_8242;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_7482;
wire n_6864;
wire n_7893;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_8331;
wire n_7090;
wire n_3786;
wire n_7158;
wire n_2888;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_6494;
wire n_5503;
wire n_8323;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_6199;
wire n_8296;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_3022;
wire n_7839;
wire n_4264;
wire n_7504;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_7360;
wire n_7681;
wire n_8076;
wire n_7301;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_8277;
wire n_3060;
wire n_4276;
wire n_7794;
wire n_7366;
wire n_8184;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_7025;
wire n_8304;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_6947;
wire n_1723;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_7309;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_6863;
wire n_6637;
wire n_798;
wire n_6100;
wire n_7860;
wire n_6735;
wire n_2659;
wire n_1414;
wire n_8212;
wire n_4975;
wire n_6358;
wire n_7911;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_7876;
wire n_6050;
wire n_2470;
wire n_7244;
wire n_7960;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_7610;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_5903;
wire n_6371;
wire n_813;
wire n_1284;
wire n_7043;
wire n_3440;
wire n_6171;
wire n_7751;
wire n_6510;
wire n_1748;
wire n_4569;
wire n_6468;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_7788;
wire n_1064;
wire n_5842;
wire n_858;
wire n_6352;
wire n_8300;
wire n_2985;
wire n_5722;
wire n_7534;
wire n_5636;
wire n_7719;
wire n_5065;
wire n_2753;
wire n_7287;
wire n_1582;
wire n_7032;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_6850;
wire n_8435;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_7119;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_2700;
wire n_7851;
wire n_1211;
wire n_6332;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_5877;
wire n_907;
wire n_3096;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_6434;
wire n_2356;
wire n_6751;
wire n_7068;
wire n_892;
wire n_4556;
wire n_6322;
wire n_8353;
wire n_5454;
wire n_7704;
wire n_2620;
wire n_7773;
wire n_6667;
wire n_7526;
wire n_1581;
wire n_6530;
wire n_4089;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_5621;
wire n_2919;
wire n_8213;
wire n_4327;
wire n_7973;
wire n_953;
wire n_4218;
wire n_6429;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_7239;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_5573;
wire n_6405;
wire n_6613;
wire n_4353;
wire n_8043;
wire n_2042;
wire n_7969;
wire n_6248;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_7821;
wire n_1854;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_6894;
wire n_1856;
wire n_7267;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_6204;
wire n_2462;
wire n_1532;
wire n_7915;
wire n_3625;
wire n_8121;
wire n_1156;
wire n_794;
wire n_7387;
wire n_7431;
wire n_7654;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_847;
wire n_4844;
wire n_6296;
wire n_2979;
wire n_5257;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_8276;
wire n_8182;
wire n_2548;
wire n_822;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_6140;
wire n_1779;
wire n_8359;
wire n_7441;
wire n_4738;
wire n_6211;
wire n_1369;
wire n_3909;
wire n_8211;
wire n_8430;
wire n_6307;
wire n_8007;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_7394;
wire n_8311;
wire n_809;
wire n_8441;
wire n_4434;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_1942;
wire n_6860;
wire n_2510;
wire n_4219;
wire n_3659;
wire n_2804;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_8198;
wire n_5697;
wire n_7188;
wire n_1810;
wire n_7573;
wire n_2813;
wire n_7879;
wire n_4438;
wire n_2009;
wire n_7087;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_7985;
wire n_6515;
wire n_6011;
wire n_8278;
wire n_7722;
wire n_7935;
wire n_6645;
wire n_8226;
wire n_3150;
wire n_747;
wire n_6984;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_7193;
wire n_3775;
wire n_4133;
wire n_6897;
wire n_7256;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_2181;
wire n_1829;
wire n_6183;
wire n_7522;
wire n_5882;
wire n_4030;
wire n_7881;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_4397;
wire n_1710;
wire n_7502;
wire n_1128;
wire n_2928;
wire n_7335;
wire n_7103;
wire n_1734;
wire n_4820;
wire n_6246;
wire n_3770;
wire n_8025;
wire n_1308;
wire n_5094;
wire n_6383;
wire n_4938;
wire n_7020;
wire n_8434;
wire n_4179;
wire n_3469;
wire n_8175;
wire n_5336;
wire n_2723;
wire n_5672;
wire n_4641;
wire n_3220;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_8046;
wire n_6904;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_8239;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_7825;
wire n_8183;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_7533;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_6611;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_906;
wire n_6116;
wire n_919;
wire n_7186;
wire n_4356;
wire n_8230;
wire n_6819;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_7936;
wire n_1740;
wire n_6473;
wire n_4291;
wire n_1586;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_8391;
wire n_6310;
wire n_7840;
wire n_1692;
wire n_2982;
wire n_8202;
wire n_2481;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_7906;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7462;
wire n_7658;
wire n_7828;
wire n_8340;
wire n_4935;
wire n_6365;
wire n_4785;
wire n_3426;
wire n_3820;
wire n_3454;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_7401;
wire n_6828;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_6355;
wire n_5596;
wire n_7887;
wire n_8058;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_6777;
wire n_5728;
wire n_2346;
wire n_8394;
wire n_4493;
wire n_3990;
wire n_7835;
wire n_3475;
wire n_1215;
wire n_8181;
wire n_1592;
wire n_6420;
wire n_6945;
wire n_2882;
wire n_1721;
wire n_7356;
wire n_2338;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_7124;
wire n_3672;
wire n_7294;
wire n_5290;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_2721;
wire n_7321;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_6754;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_7691;
wire n_5928;
wire n_3845;
wire n_7108;
wire n_6882;
wire n_2081;
wire n_7585;
wire n_4570;
wire n_7386;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7417;
wire n_7888;
wire n_2418;
wire n_7187;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_1416;
wire n_2521;
wire n_1724;
wire n_8224;
wire n_7544;
wire n_3458;
wire n_5712;
wire n_1420;
wire n_3330;
wire n_1132;
wire n_4606;
wire n_6166;
wire n_4774;
wire n_2477;
wire n_6966;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_7255;
wire n_4093;
wire n_1486;
wire n_8037;
wire n_8084;
wire n_7120;
wire n_7218;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_4174;
wire n_8289;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_8045;
wire n_5633;
wire n_2896;
wire n_8077;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_1927;
wire n_5583;
wire n_1349;
wire n_4460;
wire n_8026;
wire n_1031;
wire n_3645;
wire n_7889;
wire n_3223;
wire n_3929;
wire n_6110;
wire n_6064;
wire n_6237;
wire n_834;
wire n_7196;
wire n_2255;
wire n_2272;
wire n_893;
wire n_6341;
wire n_1965;
wire n_1902;
wire n_6590;
wire n_1941;
wire n_5501;
wire n_7923;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_6697;
wire n_874;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_7559;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_7081;
wire n_3189;
wire n_2066;
wire n_6449;
wire n_993;
wire n_7832;
wire n_7968;
wire n_3154;
wire n_1551;
wire n_6141;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_7584;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_6983;
wire n_970;
wire n_7843;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_7222;
wire n_3242;
wire n_6071;
wire n_3525;
wire n_8161;
wire n_3486;
wire n_6808;
wire n_8271;
wire n_2405;
wire n_6724;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_6571;
wire n_921;
wire n_5100;
wire n_7470;
wire n_1795;
wire n_5849;
wire n_6251;
wire n_7400;
wire n_2578;
wire n_3483;
wire n_6635;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_8056;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_7623;
wire n_3524;
wire n_5616;
wire n_7597;
wire n_5034;
wire n_6733;
wire n_1708;
wire n_7071;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_7859;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_6522;
wire n_7109;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_1776;
wire n_4807;
wire n_6562;
wire n_6150;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_8157;
wire n_1757;
wire n_890;
wire n_8346;
wire n_1919;
wire n_960;
wire n_4230;
wire n_7882;
wire n_3419;
wire n_1290;
wire n_8309;
wire n_8344;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_1252;
wire n_5754;
wire n_6016;
wire n_8096;
wire n_8100;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_7212;
wire n_1553;
wire n_3678;
wire n_7908;
wire n_2664;
wire n_8222;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_6726;
wire n_8406;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_967;
wire n_6689;
wire n_2731;
wire n_6143;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_7777;
wire n_2998;
wire n_6277;
wire n_4684;
wire n_7395;
wire n_5981;
wire n_6095;
wire n_7671;
wire n_8020;
wire n_6247;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_6880;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_1283;
wire n_762;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_6499;
wire n_6837;
wire n_4423;
wire n_4096;
wire n_7393;
wire n_2881;
wire n_8400;
wire n_6616;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_7871;
wire n_6946;
wire n_4996;
wire n_2475;
wire n_8055;
wire n_8333;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_7484;
wire n_5173;
wire n_6305;
wire n_1228;
wire n_6317;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_7649;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_945;
wire n_6693;
wire n_3743;
wire n_6734;
wire n_7135;
wire n_7014;
wire n_8263;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_984;
wire n_6382;
wire n_7328;
wire n_1983;
wire n_7635;
wire n_6404;
wire n_5975;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_6379;
wire n_7703;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_1977;
wire n_1147;
wire n_2153;
wire n_6235;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_7265;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_6789;
wire n_7184;
wire n_6440;
wire n_6417;
wire n_1470;
wire n_2318;
wire n_1735;
wire n_833;
wire n_8177;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_7728;
wire n_3442;
wire n_1201;
wire n_7690;
wire n_1114;
wire n_7219;
wire n_7479;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_7270;
wire n_1176;
wire n_5940;
wire n_8170;
wire n_1149;
wire n_7390;
wire n_1020;
wire n_7805;
wire n_7807;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_8320;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_6272;
wire n_8153;
wire n_7699;
wire n_6484;
wire n_7674;
wire n_6236;
wire n_5576;
wire n_4668;
wire n_8298;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_849;
wire n_6871;
wire n_8235;
wire n_1786;
wire n_5284;
wire n_8370;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_6768;
wire n_4759;
wire n_7951;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_7506;
wire n_2340;
wire n_3552;
wire n_875;
wire n_6717;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_5578;
wire n_2361;
wire n_8395;
wire n_1173;
wire n_1603;
wire n_969;
wire n_1401;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_8097;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_7330;
wire n_3206;
wire n_7928;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_6992;
wire n_4183;
wire n_778;
wire n_4068;
wire n_1122;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_2649;
wire n_6655;
wire n_7892;
wire n_7304;
wire n_5792;
wire n_1187;
wire n_6657;
wire n_7756;
wire n_8129;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_7990;
wire n_4625;
wire n_3914;
wire n_1174;
wire n_3324;
wire n_8122;
wire n_2558;
wire n_8259;
wire n_2063;
wire n_3803;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_2252;
wire n_7612;
wire n_6113;
wire n_7789;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_8094;
wire n_6242;
wire n_7902;
wire n_7088;
wire n_6519;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_8120;
wire n_6842;
wire n_7588;
wire n_3390;
wire n_1573;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_6801;
wire n_8099;
wire n_774;
wire n_2493;
wire n_4930;
wire n_7680;
wire n_5276;
wire n_6308;
wire n_1059;
wire n_7398;
wire n_1133;
wire n_6906;
wire n_5078;
wire n_4537;
wire n_7230;
wire n_2885;
wire n_6629;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_6968;
wire n_4282;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_6398;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_6415;
wire n_2994;
wire n_6857;
wire n_3135;
wire n_2401;
wire n_5476;
wire n_7842;
wire n_2003;
wire n_5856;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_6413;
wire n_7679;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_6361;
wire n_3438;
wire n_6231;
wire n_7783;
wire n_4098;
wire n_872;
wire n_5684;
wire n_5861;
wire n_8108;
wire n_1297;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_7862;
wire n_2806;
wire n_5312;
wire n_1184;
wire n_2184;
wire n_985;
wire n_5850;
wire n_3425;
wire n_3217;
wire n_3404;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_7820;
wire n_7167;
wire n_7833;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_7643;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_6712;
wire n_1602;
wire n_1178;
wire n_5687;
wire n_4779;
wire n_8062;
wire n_2286;
wire n_4966;
wire n_8000;
wire n_2065;
wire n_4017;
wire n_8233;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_6953;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1318;
wire n_780;
wire n_2977;
wire n_6303;
wire n_6474;
wire n_6182;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_5674;
wire n_3600;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_1388;
wire n_8352;
wire n_7993;
wire n_7930;
wire n_2836;
wire n_5682;
wire n_8385;
wire n_6392;
wire n_8166;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_7999;
wire n_5612;
wire n_6125;
wire n_6599;
wire n_7963;
wire n_6685;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_8389;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_6560;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_8439;
wire n_8369;
wire n_5301;
wire n_7800;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_7615;
wire n_5898;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1024;
wire n_7298;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_7581;
wire n_4049;
wire n_6641;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_5563;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_6673;
wire n_7172;
wire n_7074;
wire n_5497;
wire n_8234;
wire n_4724;
wire n_5832;
wire n_1238;
wire n_7190;
wire n_7112;
wire n_7678;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_5526;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_6195;
wire n_862;
wire n_3584;
wire n_6356;
wire n_3756;
wire n_2889;
wire n_7001;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_2772;
wire n_7369;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_7829;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_6559;
wire n_7359;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_7144;
wire n_4833;
wire n_6841;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_6653;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_786;
wire n_1142;
wire n_8042;
wire n_2579;
wire n_6825;
wire n_6923;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_8021;
wire n_1756;
wire n_1716;
wire n_6112;
wire n_2788;
wire n_6547;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_6399;
wire n_1873;
wire n_3201;
wire n_6275;
wire n_1087;
wire n_5666;
wire n_6575;
wire n_3472;
wire n_7924;
wire n_7732;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7191;
wire n_1247;
wire n_7459;
wire n_7096;
wire n_3050;
wire n_1478;
wire n_8280;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_6826;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_8372;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_7551;
wire n_4045;
wire n_6678;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_8282;
wire n_7750;
wire n_5015;
wire n_2702;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_6748;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_8336;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_6752;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_2209;
wire n_7652;
wire n_7808;
wire n_6500;
wire n_4270;
wire n_8135;
wire n_2797;
wire n_1255;
wire n_7051;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_6628;
wire n_844;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_6975;
wire n_1601;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_7536;
wire n_5688;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_6293;
wire n_8417;
wire n_7952;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2505;
wire n_2427;
wire n_7991;
wire n_7676;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_7553;
wire n_6905;
wire n_7425;
wire n_2594;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_8355;
wire n_4767;
wire n_7998;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_6581;
wire n_1379;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_7064;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_6577;
wire n_6899;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_8237;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_8171;
wire n_4591;
wire n_6370;
wire n_3266;
wire n_7210;
wire n_4646;
wire n_7899;
wire n_5769;
wire n_6065;
wire n_1130;
wire n_7039;
wire n_6987;
wire n_4725;
wire n_4563;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_6190;
wire n_6859;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_6309;
wire n_6623;
wire n_7723;
wire n_2426;
wire n_6527;
wire n_7443;
wire n_7811;
wire n_5341;
wire n_4320;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_6929;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_8279;
wire n_5622;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_7348;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_2689;
wire n_3259;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_7155;
wire n_8227;
wire n_3688;
wire n_6865;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_6535;
wire n_904;
wire n_3338;
wire n_7213;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_8270;
wire n_4209;
wire n_1271;
wire n_5966;
wire n_1542;
wire n_7456;
wire n_8335;
wire n_5041;
wire n_7420;
wire n_8054;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_3261;
wire n_2200;
wire n_6482;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_8150;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_7715;
wire n_1780;
wire n_3732;
wire n_6605;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_7007;
wire n_8358;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_7909;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_8281;
wire n_5908;
wire n_6018;
wire n_4202;
wire n_7168;
wire n_5212;
wire n_7736;
wire n_5000;
wire n_8396;
wire n_2853;
wire n_1323;
wire n_5939;
wire n_7177;
wire n_3766;
wire n_1353;
wire n_800;
wire n_7780;
wire n_2880;
wire n_7379;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_8223;
wire n_5931;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_7813;
wire n_864;
wire n_7030;
wire n_5420;
wire n_1264;
wire n_6311;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_6424;
wire n_6654;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_1607;
wire n_8379;
wire n_6879;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_5679;
wire n_947;
wire n_5938;
wire n_3710;
wire n_6702;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_1230;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_6452;
wire n_929;
wire n_3379;
wire n_4374;
wire n_6791;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_7280;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_6915;
wire n_7110;
wire n_1104;
wire n_1294;
wire n_7511;
wire n_1257;
wire n_6856;
wire n_1182;
wire n_7941;
wire n_7791;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_7232;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_6364;
wire n_6451;
wire n_6552;
wire n_1845;
wire n_2193;
wire n_8325;
wire n_2478;
wire n_5140;
wire n_6328;
wire n_4816;
wire n_8382;
wire n_7827;
wire n_1483;
wire n_6363;
wire n_2983;
wire n_7159;
wire n_8127;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_6406;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_6978;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_8232;
wire n_2651;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_7363;
wire n_6612;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_955;
wire n_5511;
wire n_7863;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_1146;
wire n_7295;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_897;
wire n_5280;
wire n_6375;
wire n_6479;
wire n_1428;
wire n_6866;
wire n_7831;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_6170;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_7466;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_6130;
wire n_1513;
wire n_2970;
wire n_7651;
wire n_2235;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_8179;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_6935;
wire n_1590;
wire n_7530;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_8308;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_8378;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_6907;
wire n_6158;
wire n_7661;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_8412;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_7145;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_6338;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_8425;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_8241;
wire n_7823;
wire n_7467;
wire n_5097;
wire n_7932;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_7541;
wire n_2784;
wire n_3718;
wire n_3470;
wire n_4862;
wire n_3092;
wire n_7241;
wire n_7717;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_4850;
wire n_6625;
wire n_3781;
wire n_4912;
wire n_4813;
wire n_7464;
wire n_2590;
wire n_6302;
wire n_8274;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_8152;
wire n_3328;
wire n_6706;
wire n_944;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_8264;
wire n_7434;
wire n_7636;
wire n_6999;
wire n_7054;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_6228;
wire n_857;
wire n_5650;
wire n_2636;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_4702;
wire n_6888;
wire n_8266;
wire n_4252;
wire n_4457;
wire n_6063;
wire n_971;
wire n_6800;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_6922;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_7503;
wire n_2808;
wire n_6070;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7273;
wire n_6647;
wire n_7296;
wire n_2930;
wire n_5733;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_7543;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_6184;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_7507;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_7555;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_914;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_7578;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_759;
wire n_8195;
wire n_5585;
wire n_6397;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_7033;
wire n_6121;
wire n_1571;
wire n_3119;
wire n_7531;
wire n_4142;
wire n_4082;
wire n_1189;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_8377;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_6954;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_5875;
wire n_8428;
wire n_8103;
wire n_4262;
wire n_2671;
wire n_6646;
wire n_8414;
wire n_8362;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_7131;
wire n_7769;
wire n_6903;
wire n_1647;
wire n_4685;
wire n_6101;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_6941;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_8324;
wire n_6106;
wire n_6604;
wire n_4014;
wire n_7418;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_7688;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_8348;
wire n_5607;
wire n_1615;
wire n_4175;
wire n_8288;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_8269;
wire n_5006;
wire n_7806;
wire n_6566;
wire n_1443;
wire n_946;
wire n_1539;
wire n_5734;
wire n_6081;
wire n_4892;
wire n_7204;
wire n_3823;
wire n_8180;
wire n_1866;
wire n_4173;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_8306;
wire n_6047;
wire n_2960;
wire n_8167;
wire n_1090;
wire n_5438;
wire n_4627;
wire n_758;
wire n_7354;
wire n_7448;
wire n_6244;
wire n_2290;
wire n_6861;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_7852;
wire n_1049;
wire n_2145;
wire n_5725;
wire n_1639;
wire n_7925;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_5163;
wire n_2039;
wire n_7748;
wire n_5768;
wire n_4961;
wire n_7556;
wire n_3753;
wire n_7640;
wire n_8187;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_7422;
wire n_7920;
wire n_8433;
wire n_2509;
wire n_4317;
wire n_3236;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_6588;
wire n_3396;
wire n_1445;
wire n_7900;
wire n_7050;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_7136;
wire n_8316;
wire n_7318;
wire n_6055;
wire n_5138;
wire n_1017;
wire n_8397;
wire n_5374;
wire n_6108;
wire n_8115;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_6165;
wire n_1828;
wire n_6621;
wire n_2320;
wire n_1045;
wire n_7175;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_7810;
wire n_4640;
wire n_2583;
wire n_6323;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_2087;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_6597;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_7817;
wire n_8294;
wire n_2523;
wire n_6933;
wire n_4387;
wire n_7878;
wire n_8338;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_1578;
wire n_7289;
wire n_5805;
wire n_7665;
wire n_8131;
wire n_3719;
wire n_7855;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_7764;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_8027;
wire n_6216;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_8162;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_2725;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_7263;
wire n_743;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_6911;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_6327;
wire n_2595;
wire n_761;
wire n_6607;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_7850;
wire n_7509;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_7240;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_7725;
wire n_8398;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_4614;
wire n_1265;
wire n_8307;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_8010;
wire n_1015;
wire n_7278;
wire n_1651;
wire n_8347;
wire n_7630;
wire n_2775;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_1101;
wire n_8354;
wire n_4326;
wire n_1106;
wire n_6695;
wire n_3557;
wire n_8204;
wire n_2230;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_7565;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_7883;
wire n_1455;
wire n_6600;
wire n_767;
wire n_2490;
wire n_1407;
wire n_7410;
wire n_4213;
wire n_2849;
wire n_7097;
wire n_3692;
wire n_2204;
wire n_6421;
wire n_5747;
wire n_7414;
wire n_7495;
wire n_5969;
wire n_8312;
wire n_4929;
wire n_8040;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_6458;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_6746;
wire n_8132;
wire n_2508;
wire n_4031;
wire n_7586;
wire n_7720;
wire n_6719;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_2461;
wire n_6506;
wire n_2243;
wire n_4583;
wire n_6287;
wire n_6662;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_6851;
wire n_8116;
wire n_6687;
wire n_2890;
wire n_6884;
wire n_2554;
wire n_8356;
wire n_8013;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_1082;
wire n_3961;
wire n_1630;
wire n_6780;
wire n_6513;
wire n_4891;
wire n_7841;
wire n_6619;
wire n_8193;
wire n_1023;
wire n_5603;
wire n_6804;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_6516;
wire n_5208;
wire n_7490;
wire n_1056;
wire n_3588;
wire n_7792;
wire n_6924;
wire n_2308;
wire n_4590;
wire n_7492;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_8329;
wire n_5237;
wire n_7809;
wire n_4664;
wire n_3860;
wire n_8154;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_7073;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_6788;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_6393;
wire n_2333;
wire n_8086;
wire n_2916;
wire n_6249;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_6572;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_7569;
wire n_7003;
wire n_7897;
wire n_4773;
wire n_7962;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_2472;
wire n_4611;
wire n_8113;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_7419;
wire n_5827;
wire n_1560;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_7784;
wire n_1953;
wire n_4422;
wire n_6123;
wire n_6934;
wire n_2589;
wire n_7094;
wire n_7500;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_6082;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_7864;
wire n_5228;
wire n_1504;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_7790;
wire n_3572;
wire n_992;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_842;
wire n_8107;
wire n_7642;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_7045;
wire n_1643;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_7238;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_7126;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_7931;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3078;
wire n_6979;
wire n_6203;
wire n_7405;
wire n_7739;
wire n_894;
wire n_3253;
wire n_7207;
wire n_4027;
wire n_7934;
wire n_831;
wire n_2280;
wire n_7454;
wire n_4599;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_6596;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_6870;
wire n_7639;
wire n_5613;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_7251;
wire n_2303;
wire n_7776;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_7059;
wire n_8255;
wire n_7035;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_8029;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_6713;
wire n_5513;
wire n_6747;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_5132;
wire n_830;
wire n_5191;
wire n_6333;
wire n_6262;
wire n_3085;
wire n_5869;
wire n_8130;
wire n_5925;
wire n_1655;
wire n_749;
wire n_6240;
wire n_5359;
wire n_6412;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_7782;
wire n_7220;
wire n_4316;
wire n_939;
wire n_3697;
wire n_7438;
wire n_1232;
wire n_2638;
wire n_7515;
wire n_7574;
wire n_4044;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_7065;
wire n_1338;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_7894;
wire n_1522;
wire n_7868;
wire n_6973;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_7285;
wire n_8286;
wire n_5200;
wire n_1653;
wire n_5659;
wire n_1506;
wire n_5618;
wire n_6325;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_8178;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_7008;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_8432;
wire n_6111;
wire n_1834;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_8047;
wire n_6260;
wire n_7501;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_6665;
wire n_7566;
wire n_7937;
wire n_7055;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_8268;
wire n_8053;
wire n_5858;
wire n_5817;
wire n_6690;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_7113;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_7872;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_7242;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_2205;
wire n_1777;
wire n_1335;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_7954;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_7819;
wire n_6570;
wire n_1410;
wire n_8022;
wire n_8415;
wire n_6498;
wire n_3902;
wire n_4730;
wire n_7228;
wire n_6692;
wire n_937;
wire n_6074;
wire n_2779;
wire n_7561;
wire n_1584;
wire n_6380;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_8386;
wire n_8426;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_7994;
wire n_6045;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_2811;
wire n_3348;
wire n_7415;
wire n_7793;
wire n_5796;
wire n_7702;
wire n_7598;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_895;
wire n_3358;
wire n_8192;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_6772;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_6823;
wire n_6877;
wire n_6806;
wire n_7426;
wire n_5906;
wire n_8350;
wire n_4743;
wire n_1067;
wire n_3805;
wire n_7957;
wire n_3825;
wire n_8048;
wire n_6831;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_7217;
wire n_2692;
wire n_2008;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_799;
wire n_6785;
wire n_8254;
wire n_1213;
wire n_6374;
wire n_6930;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_7735;
wire n_8265;
wire n_1689;
wire n_8049;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_6838;
wire n_869;
wire n_5736;
wire n_6937;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_1352;
wire n_2197;
wire n_7558;
wire n_2199;
wire n_5069;
wire n_7442;
wire n_8272;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_6674;
wire n_2480;
wire n_6034;
wire n_7499;
wire n_2363;
wire n_4072;
wire n_916;
wire n_5579;
wire n_1115;
wire n_8381;
wire n_7085;
wire n_4781;
wire n_3606;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_2550;
wire n_6762;
wire n_7341;
wire n_7895;
wire n_4424;
wire n_823;
wire n_8366;
wire n_8101;
wire n_7611;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_8384;
wire n_5642;
wire n_3553;
wire n_7224;
wire n_5880;
wire n_6169;
wire n_4746;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_1683;
wire n_1530;
wire n_8023;
wire n_8052;
wire n_997;
wire n_7627;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_2996;
wire n_1268;
wire n_5793;
wire n_5591;
wire n_7856;
wire n_1320;
wire n_4050;
wire n_7496;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_5623;
wire n_1063;
wire n_5681;
wire n_4853;
wire n_981;
wire n_7399;
wire n_867;
wire n_2422;
wire n_6213;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_7605;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_6814;
wire n_7342;
wire n_2057;
wire n_4008;
wire n_8014;
wire n_5507;
wire n_905;
wire n_7214;
wire n_7472;
wire n_5077;
wire n_782;
wire n_8371;
wire n_5872;
wire n_3858;
wire n_7408;
wire n_8231;
wire n_1901;
wire n_6115;
wire n_4502;
wire n_6858;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_1330;
wire n_8164;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_7837;
wire n_8357;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_8143;
wire n_6430;
wire n_6193;
wire n_934;
wire n_5314;
wire n_6462;
wire n_1618;
wire n_8422;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_6518;
wire n_6797;
wire n_2799;
wire n_4454;
wire n_7938;
wire n_8253;
wire n_4229;
wire n_1083;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_787;
wire n_6916;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_7812;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_6152;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_8243;
wire n_1577;
wire n_8236;
wire n_8292;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_5777;
wire n_2764;
wire n_7949;
wire n_1498;
wire n_7046;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_8011;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_6589;
wire n_7579;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_8139;
wire n_8123;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_7917;
wire n_5951;
wire n_7092;
wire n_2442;
wire n_6197;
wire n_6971;
wire n_928;
wire n_8424;
wire n_1943;
wire n_7460;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_8156;
wire n_3351;
wire n_3527;
wire n_7698;
wire n_7886;
wire n_6154;
wire n_7344;
wire n_1396;
wire n_1348;
wire n_6020;
wire n_2883;
wire n_1752;
wire n_7904;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_7079;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_7774;
wire n_5797;
wire n_7922;
wire n_8189;
wire n_6696;
wire n_4839;
wire n_5222;
wire n_8285;
wire n_5743;
wire n_1028;
wire n_4016;
wire n_6210;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_6964;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_8117;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_7670;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_6681;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_6661;
wire n_8018;
wire n_3303;
wire n_1654;
wire n_6640;
wire n_3916;
wire n_7940;
wire n_2569;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_6455;
wire n_2196;
wire n_3591;
wire n_7721;
wire n_4273;
wire n_3024;
wire n_7606;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_6832;
wire n_7836;
wire n_1595;
wire n_2161;
wire n_6160;
wire n_7564;
wire n_2404;
wire n_2083;
wire n_7884;
wire n_6718;
wire n_2503;
wire n_6542;
wire n_1540;
wire n_1936;
wire n_6031;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_2500;
wire n_7653;
wire n_1918;
wire n_5656;
wire n_863;
wire n_6763;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_2414;
wire n_6438;
wire n_1402;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_6758;
wire n_2004;
wire n_7976;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_6874;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_8341;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_6030;
wire n_8199;
wire n_6077;
wire n_8005;
wire n_4119;
wire n_3799;
wire n_7743;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_4474;
wire n_1089;
wire n_6386;
wire n_5217;
wire n_1004;
wire n_8016;
wire n_5957;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_8283;
wire n_3585;
wire n_2975;
wire n_7655;
wire n_5490;
wire n_5029;
wire n_8291;
wire n_2704;
wire n_4214;
wire n_8176;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7737;
wire n_7433;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_7347;
wire n_8145;
wire n_4580;
wire n_6792;
wire n_7633;
wire n_1263;
wire n_6177;
wire n_5912;
wire n_1126;
wire n_7798;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_1859;
wire n_1677;
wire n_5557;
wire n_7397;
wire n_7389;
wire n_5472;
wire n_7602;
wire n_2955;
wire n_4112;
wire n_8069;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_5396;
wire n_7693;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_6557;
wire n_7300;
wire n_956;
wire n_2134;
wire n_5960;
wire n_8041;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_7532;
wire n_5143;
wire n_7724;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_1545;
wire n_2374;
wire n_5859;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_854;
wire n_4734;
wire n_8374;
wire n_1939;
wire n_2486;
wire n_6163;
wire n_4635;
wire n_3501;
wire n_1152;
wire n_7118;
wire n_1869;
wire n_8006;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_6285;
wire n_6778;
wire n_7946;
wire n_6025;
wire n_7257;
wire n_4242;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_7933;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_8409;
wire n_7669;
wire n_5268;
wire n_6318;
wire n_8215;
wire n_8220;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_7927;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_7910;
wire n_1261;
wire n_6315;
wire n_938;
wire n_3186;
wire n_7970;
wire n_4955;
wire n_1154;
wire n_8407;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_6343;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_920;
wire n_2515;
wire n_7865;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_6886;
wire n_1949;
wire n_976;
wire n_1946;
wire n_2936;
wire n_6912;
wire n_8326;
wire n_5914;
wire n_775;
wire n_8250;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_8408;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_7252;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_7133;
wire n_1850;
wire n_6883;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_8155;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_7518;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_6378;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_8275;
wire n_1218;
wire n_2632;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_1547;
wire n_777;
wire n_6407;
wire n_1755;
wire n_8297;
wire n_6749;
wire n_6839;
wire n_7711;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_7705;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_4942;
wire n_6217;
wire n_6680;
wire n_5844;
wire n_2432;
wire n_7972;
wire n_1521;
wire n_6532;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_8072;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_7854;
wire n_2337;
wire n_7707;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_8050;
wire n_6736;
wire n_5344;
wire n_923;
wire n_6526;
wire n_8142;
wire n_4629;
wire n_6339;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_8151;
wire n_6350;
wire n_7013;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_4376;
wire n_3986;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_7656;
wire n_3885;
wire n_6845;
wire n_7105;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_5574;
wire n_5126;
wire n_1039;
wire n_6508;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_7570;
wire n_8246;
wire n_7771;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_2688;
wire n_5368;
wire n_1202;
wire n_8057;
wire n_8349;
wire n_5626;
wire n_6603;
wire n_6114;
wire n_1463;
wire n_6576;
wire n_3651;
wire n_7943;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_7208;
wire n_6245;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_7714;
wire n_4815;
wire n_7202;
wire n_4246;
wire n_3580;
wire n_7011;
wire n_2139;
wire n_4609;
wire n_7621;
wire n_5291;
wire n_8068;
wire n_5876;
wire n_6970;
wire n_5114;
wire n_2674;
wire n_6409;
wire n_6704;
wire n_1565;
wire n_4088;
wire n_6876;
wire n_7778;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_7028;
wire n_4472;
wire n_4462;
wire n_3433;
wire n_7313;
wire n_6255;
wire n_7320;
wire n_7343;
wire n_1072;
wire n_5288;
wire n_5540;
wire n_2305;
wire n_5699;
wire n_7525;
wire n_2450;
wire n_7875;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_6938;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_8327;
wire n_2625;
wire n_2271;
wire n_7337;
wire n_6989;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_3989;
wire n_4475;
wire n_7753;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_8168;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_8392;
wire n_7038;
wire n_4683;
wire n_5366;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_6360;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_887;
wire n_6270;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_8419;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_1997;
wire n_6691;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_7392;
wire n_2215;
wire n_5053;
wire n_7912;
wire n_8245;
wire n_1259;
wire n_6239;
wire n_4553;
wire n_746;
wire n_6803;
wire n_7919;
wire n_784;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_4809;
wire n_8109;
wire n_5226;
wire n_1244;
wire n_7657;
wire n_1925;
wire n_3660;
wire n_7995;
wire n_1815;
wire n_5867;
wire n_6048;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_913;
wire n_6773;
wire n_3833;
wire n_5632;
wire n_865;
wire n_8390;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_6336;
wire n_3814;
wire n_7041;
wire n_1415;
wire n_2592;
wire n_7802;
wire n_2838;
wire n_4911;
wire n_4842;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_1191;
wire n_7557;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_6776;
wire n_3128;
wire n_5426;
wire n_6463;
wire n_744;
wire n_2631;
wire n_7896;
wire n_2178;
wire n_1767;
wire n_6372;
wire n_7176;
wire n_1529;
wire n_2469;
wire n_5625;
wire n_5778;
wire n_6396;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_6669;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_7826;
wire n_3000;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_7590;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_8208;
wire n_1933;
wire n_6995;
wire n_7185;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_6254;
wire n_6161;
wire n_3457;
wire n_1678;
wire n_7987;
wire n_8134;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_908;
wire n_6128;
wire n_4086;
wire n_7037;
wire n_2412;
wire n_4814;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_8427;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_959;
wire n_3031;
wire n_7258;
wire n_7432;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_6334;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_6848;
wire n_8345;
wire n_2171;
wire n_4708;
wire n_6321;
wire n_7765;
wire n_2768;
wire n_2314;
wire n_6794;
wire n_4826;
wire n_3343;
wire n_2420;
wire n_1079;
wire n_7761;
wire n_7197;
wire n_5489;
wire n_1593;
wire n_6400;
wire n_3767;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_2299;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_6705;
wire n_7775;
wire n_2162;
wire n_7619;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_750;
wire n_742;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_8083;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_6495;
wire n_5013;
wire n_2312;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5569;
wire n_8038;
wire n_5439;
wire n_8229;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_6481;
wire n_3607;
wire n_4925;
wire n_7548;
wire n_1921;
wire n_1309;
wire n_6534;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_6181;
wire n_3276;
wire n_1177;
wire n_6728;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_8085;
wire n_6133;
wire n_6528;
wire n_7604;
wire n_7407;
wire n_1119;
wire n_1240;
wire n_8185;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_6670;
wire n_6774;
wire n_8365;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_6038;
wire n_4818;
wire n_7727;
wire n_4514;
wire n_4800;
wire n_1366;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_6282;
wire n_1568;
wire n_2110;
wire n_8035;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_6700;
wire n_7334;
wire n_7684;
wire n_1591;
wire n_2033;
wire n_7755;
wire n_8098;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_5932;
wire n_6178;
wire n_1111;
wire n_2132;
wire n_6234;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_7787;
wire n_4140;
wire n_8067;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_7849;
wire n_5186;
wire n_7367;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_6715;
wire n_5828;
wire n_2831;
wire n_7200;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_6337;
wire n_4868;
wire n_1885;
wire n_8332;
wire n_2452;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_7877;
wire n_1849;
wire n_1131;
wire n_7799;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_5631;
wire n_8028;
wire n_2467;
wire n_6539;
wire n_1094;
wire n_7243;
wire n_7179;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_1209;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_5326;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_8404;
wire n_4669;
wire n_4339;
wire n_6595;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_7738;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_8073;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_7785;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_7373;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_6257;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_6852;
wire n_2789;
wire n_6346;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_764;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_7587;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_7874;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_2328;
wire n_7760;
wire n_4248;
wire n_5915;
wire n_6818;
wire n_5452;
wire n_7226;
wire n_4754;
wire n_7057;
wire n_7685;
wire n_8031;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6753;
wire n_6815;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_7730;
wire n_8405;
wire n_1699;
wire n_3334;
wire n_7913;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_6764;
wire n_5535;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_7706;
wire n_7891;
wire n_6391;
wire n_4003;
wire n_8088;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_1050;
wire n_841;
wire n_4586;
wire n_4048;
wire n_1954;
wire n_6471;
wire n_1844;
wire n_3777;
wire n_6627;
wire n_5761;
wire n_4784;
wire n_7203;
wire n_8429;
wire n_2999;
wire n_7512;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_7215;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_7388;
wire n_7694;
wire n_1179;
wire n_6243;
wire n_753;
wire n_6488;
wire n_4286;
wire n_1048;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_6457;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_7982;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_8225;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_6867;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_1688;
wire n_6633;
wire n_8080;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_6574;
wire n_1992;
wire n_6395;
wire n_4402;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_7996;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3382;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_7198;
wire n_1557;
wire n_4201;
wire n_6784;
wire n_6168;
wire n_896;
wire n_8431;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_2192;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_7950;
wire n_7249;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_814;
wire n_2707;
wire n_6799;
wire n_8015;
wire n_5920;
wire n_6672;
wire n_2471;
wire n_1472;
wire n_6149;
wire n_1671;
wire n_8256;
wire n_7142;
wire n_3230;
wire n_5808;
wire n_3342;
wire n_1062;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_7916;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_6450;
wire n_3729;
wire n_8074;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_783;
wire n_1928;
wire n_8039;
wire n_5244;
wire n_6523;
wire n_5382;
wire n_8065;
wire n_1188;
wire n_6107;
wire n_3957;
wire n_6775;
wire n_5274;
wire n_3848;
wire n_8194;
wire n_4284;
wire n_2600;
wire n_8207;
wire n_3919;
wire n_6232;
wire n_6445;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_3608;
wire n_6056;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_7759;
wire n_2352;
wire n_7818;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_8217;
wire n_1110;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_1088;
wire n_8437;
wire n_5249;
wire n_3393;
wire n_7447;
wire n_866;
wire n_7944;
wire n_5198;
wire n_5360;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_6252;
wire n_5866;
wire n_6493;
wire n_7947;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_5899;
wire n_7629;
wire n_8051;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_7601;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_7757;
wire n_8030;
wire n_5865;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_7138;
wire n_7290;
wire n_8249;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_6679;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_5924;
wire n_2206;
wire n_3182;
wire n_7625;
wire n_5822;
wire n_2564;
wire n_6259;
wire n_4947;
wire n_876;
wire n_7284;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_3450;
wire n_966;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_7971;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_6630;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_6279;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_1168;
wire n_6813;
wire n_5564;
wire n_8273;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_7106;
wire n_6042;
wire n_7644;
wire n_1853;
wire n_1356;
wire n_6057;
wire n_1787;
wire n_4137;
wire n_7529;
wire n_6675;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_6476;
wire n_8200;
wire n_3972;
wire n_7907;
wire n_8188;
wire n_6207;
wire n_5539;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_3308;
wire n_6524;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_8267;
wire n_1720;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_7199;
wire n_5273;
wire n_8360;
wire n_4677;
wire n_3901;
wire n_8036;
wire n_1480;
wire n_5261;
wire n_6520;
wire n_7853;
wire n_7648;
wire n_3757;
wire n_8393;
wire n_8160;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_7866;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_1170;
wire n_6425;
wire n_2213;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_7638;
wire n_5703;
wire n_8240;
wire n_4634;
wire n_3337;
wire n_7988;
wire n_2527;
wire n_855;
wire n_5534;
wire n_6432;
wire n_1461;
wire n_3204;
wire n_8258;
wire n_7259;
wire n_2136;
wire n_6540;
wire n_6955;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_7237;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_4506;
wire n_2375;
wire n_6388;
wire n_5904;
wire n_4880;
wire n_6760;
wire n_1907;
wire n_2686;
wire n_8009;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_1417;
wire n_5061;
wire n_1295;
wire n_5572;
wire n_5750;
wire n_7063;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_8012;
wire n_7576;
wire n_1762;
wire n_1013;
wire n_8008;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_8079;
wire n_6664;
wire n_5815;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_6487;
wire n_4737;
wire n_7734;
wire n_6729;
wire n_3647;
wire n_5755;
wire n_825;
wire n_2819;
wire n_5949;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_7858;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_7385;
wire n_3720;
wire n_4535;
wire n_7668;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_5955;
wire n_7476;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_792;
wire n_8436;
wire n_8124;
wire n_8148;
wire n_8033;
wire n_6843;
wire n_3140;
wire n_7953;
wire n_8343;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_8118;
wire n_2104;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_4196;
wire n_6969;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_6485;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5783;
wire n_5183;
wire n_6075;
wire n_7082;
wire n_3084;
wire n_6120;
wire n_1727;
wire n_6659;
wire n_2735;
wire n_6750;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_1046;
wire n_8376;
wire n_3761;
wire n_7689;
wire n_4889;
wire n_7132;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_7824;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_7796;
wire n_6478;
wire n_2172;
wire n_6066;
wire n_7034;
wire n_6086;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_1129;
wire n_8303;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_7084;
wire n_5845;
wire n_7293;
wire n_1225;
wire n_8251;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_7253;
wire n_2423;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_994;
wire n_8003;
wire n_6410;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_6059;
wire n_5130;
wire n_1567;
wire n_7520;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_6267;
wire n_8165;
wire n_1797;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_1250;
wire n_8330;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_6610;
wire n_7918;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7514;
wire n_7163;
wire n_7620;
wire n_2570;
wire n_1086;
wire n_1858;
wire n_1619;
wire n_5473;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_5946;
wire n_2744;
wire n_6711;
wire n_4287;
wire n_2397;
wire n_7445;
wire n_2208;
wire n_6847;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_7123;
wire n_6384;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_7959;
wire n_1676;
wire n_1113;
wire n_7563;
wire n_6298;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_7361;
wire n_852;
wire n_4602;
wire n_5172;
wire n_8186;
wire n_4449;
wire n_1864;
wire n_7322;
wire n_8219;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_5070;
wire n_6377;
wire n_1337;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_1627;
wire n_4870;
wire n_1245;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_6348;
wire n_7713;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_6834;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_2823;
wire n_1076;
wire n_1408;
wire n_1761;
wire n_8066;
wire n_5874;
wire n_7977;
wire n_8342;
wire n_7508;
wire n_7021;
wire n_5270;
wire n_5956;
wire n_7834;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_6078;
wire n_7000;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_7921;
wire n_2655;
wire n_4185;
wire n_8402;
wire n_4797;
wire n_2366;
wire n_7130;
wire n_1526;
wire n_5823;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_7538;
wire n_7517;
wire n_1583;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_7077;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_6642;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_7333;
wire n_4364;
wire n_4245;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_6942;
wire n_8418;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_6511;
wire n_3721;
wire n_1254;
wire n_6507;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_1032;
wire n_7319;
wire n_7997;
wire n_2991;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_6606;
wire n_4560;
wire n_3473;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_8144;
wire n_3699;
wire n_5067;
wire n_7107;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_7469;
wire n_2728;
wire n_3857;
wire n_8111;

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_353),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_525),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_136),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_658),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_20),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_549),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_150),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_491),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_196),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_385),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_731),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_102),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_236),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_427),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_210),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_130),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_658),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_394),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_495),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_605),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_603),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_419),
.Y(n_760)
);

BUFx10_ASAP7_75t_L g761 ( 
.A(n_16),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_389),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_283),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_513),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_86),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_661),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_603),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_202),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_383),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_691),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_476),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_184),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_148),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_49),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_360),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_287),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_195),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_233),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_136),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_66),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_213),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_246),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_582),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_445),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_498),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_295),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_623),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_228),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_621),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_556),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_246),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_506),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_131),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_459),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_403),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_3),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_284),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_175),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_539),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_722),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_637),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_542),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_165),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_249),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_3),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_451),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_103),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_516),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_192),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_628),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_596),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_443),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_103),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_724),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_224),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_461),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_243),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_173),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_513),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_202),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_702),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_114),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_99),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_703),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_87),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_308),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_427),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_510),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_632),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_696),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_122),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_1),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_109),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_567),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_557),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_121),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_492),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_416),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_31),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_360),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_133),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_28),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_425),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_487),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_247),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_135),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_375),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_505),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_355),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_539),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_439),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_298),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_176),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_260),
.Y(n_854)
);

CKINVDCx16_ASAP7_75t_R g855 ( 
.A(n_440),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_83),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_305),
.Y(n_857)
);

CKINVDCx14_ASAP7_75t_R g858 ( 
.A(n_38),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_387),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_505),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_712),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_74),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_290),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_264),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_358),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_357),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_479),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_183),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_215),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_297),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_694),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_119),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_384),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_449),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_323),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_586),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_234),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_396),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_415),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_643),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_104),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_481),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_461),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_243),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_675),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_480),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_546),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_340),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_33),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_683),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_363),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_328),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_259),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_592),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_174),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_225),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_719),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_241),
.Y(n_898)
);

CKINVDCx14_ASAP7_75t_R g899 ( 
.A(n_218),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_654),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_286),
.Y(n_901)
);

BUFx10_ASAP7_75t_L g902 ( 
.A(n_677),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_24),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_451),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_717),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_295),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_479),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_416),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_411),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_478),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_212),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_421),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_102),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_36),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_483),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_297),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_349),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_235),
.Y(n_918)
);

CKINVDCx14_ASAP7_75t_R g919 ( 
.A(n_331),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_106),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_69),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_366),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_620),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_604),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_325),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_733),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_498),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_292),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_609),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_643),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_158),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_566),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_478),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_689),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_726),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_618),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_81),
.Y(n_937)
);

BUFx5_ASAP7_75t_L g938 ( 
.A(n_358),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_454),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_76),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_29),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_181),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_618),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_420),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_463),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_527),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_392),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_493),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_39),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_722),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_160),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_135),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_443),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_83),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_464),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_650),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_387),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_364),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_362),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_577),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_115),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_325),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_411),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_268),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_58),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_244),
.Y(n_966)
);

CKINVDCx14_ASAP7_75t_R g967 ( 
.A(n_568),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_523),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_69),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_66),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_575),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_33),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_384),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_687),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_184),
.Y(n_975)
);

BUFx10_ASAP7_75t_L g976 ( 
.A(n_698),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_442),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_711),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_349),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_493),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_264),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_169),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_656),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_487),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_286),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_244),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_446),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_171),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_21),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_283),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_467),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_31),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_401),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_521),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_398),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_81),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_664),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_552),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_421),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_375),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_694),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_524),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_590),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_506),
.Y(n_1004)
);

CKINVDCx14_ASAP7_75t_R g1005 ( 
.A(n_622),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_168),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_444),
.Y(n_1007)
);

BUFx8_ASAP7_75t_SL g1008 ( 
.A(n_459),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_122),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_104),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_734),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_125),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_452),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_685),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_233),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_158),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_307),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_336),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_280),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_24),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_640),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_367),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_198),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_692),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_692),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_168),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_484),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_404),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_321),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_248),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_702),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_361),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_270),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_159),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_163),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_638),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_525),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_381),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_2),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_57),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_355),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_583),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_97),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_473),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_610),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_203),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_489),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_304),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_301),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_563),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_728),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_257),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_322),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_631),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_364),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_92),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_262),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_288),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_589),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_323),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_637),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_27),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_414),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_704),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_330),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_35),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_137),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_259),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_544),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_106),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_9),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_569),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_596),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_187),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_79),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_510),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_153),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_584),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_390),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_569),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_431),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_185),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_471),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_701),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_220),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_684),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_276),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_418),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_111),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_509),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_436),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_567),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_337),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_663),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_203),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_216),
.Y(n_1096)
);

INVx4_ASAP7_75t_R g1097 ( 
.A(n_121),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_296),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_407),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_336),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_576),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_561),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_684),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_127),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_598),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_68),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_672),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_256),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_215),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_256),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_241),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_36),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_90),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_281),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_725),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_19),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_61),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_312),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_634),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_610),
.Y(n_1120)
);

CKINVDCx14_ASAP7_75t_R g1121 ( 
.A(n_685),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_645),
.Y(n_1122)
);

BUFx5_ASAP7_75t_L g1123 ( 
.A(n_621),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_258),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_483),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_234),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_337),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_32),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_709),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_291),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_174),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_620),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_273),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_428),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_471),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_45),
.Y(n_1136)
);

CKINVDCx16_ASAP7_75t_R g1137 ( 
.A(n_564),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_491),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_450),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_632),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_363),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_371),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_662),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_11),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_405),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_545),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_342),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_393),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_515),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_204),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_150),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_263),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_661),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_368),
.Y(n_1154)
);

CKINVDCx14_ASAP7_75t_R g1155 ( 
.A(n_133),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_199),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_499),
.Y(n_1157)
);

BUFx10_ASAP7_75t_L g1158 ( 
.A(n_22),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_669),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_294),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_86),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_408),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_11),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_732),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_55),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_181),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_251),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_324),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_177),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_204),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_437),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_96),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_677),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_187),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_383),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_581),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_156),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_94),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_79),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_149),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_27),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_507),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_172),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_463),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_308),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_226),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_315),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_500),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_115),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_535),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_597),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_721),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_9),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_345),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_572),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_12),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_663),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_650),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_80),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_198),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_302),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_172),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_43),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_142),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_408),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_143),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_622),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_595),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_226),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_626),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_467),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_324),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_108),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_563),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_263),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_59),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_365),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_673),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_630),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_652),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_475),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_17),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_42),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_191),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_111),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_85),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_385),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_688),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_609),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_217),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_455),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_124),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_496),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_472),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_401),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_84),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_690),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_676),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_209),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_432),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_16),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_189),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_298),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_18),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_575),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_377),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_240),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_351),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_484),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_649),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_379),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_98),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_208),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_14),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_735),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_91),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_113),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_161),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_192),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_604),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_730),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_294),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_213),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_180),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_593),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_289),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_394),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_693),
.Y(n_1269)
);

BUFx10_ASAP7_75t_L g1270 ( 
.A(n_92),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_80),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_535),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_521),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_320),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_469),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_290),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_229),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_37),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_5),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_151),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_141),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_23),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_207),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_359),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_74),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_186),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_139),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_577),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_690),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_634),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_409),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_376),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_727),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_112),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_682),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_585),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_193),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_502),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_141),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_55),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_546),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_281),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1115),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1115),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_938),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1008),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_938),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_938),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_749),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_967),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1005),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_938),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_938),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_938),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_858),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_938),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_858),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_899),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_899),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_793),
.Y(n_1320)
);

BUFx10_ASAP7_75t_L g1321 ( 
.A(n_753),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_938),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_919),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_938),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_919),
.Y(n_1325)
);

CKINVDCx16_ASAP7_75t_R g1326 ( 
.A(n_1299),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_938),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1121),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1123),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_753),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1121),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_799),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1155),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1123),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_806),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1123),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1123),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1123),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1123),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1123),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1155),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1123),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_793),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1123),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1299),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_855),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1123),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_814),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_844),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_844),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_855),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_844),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_844),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_799),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1068),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_799),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1068),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1137),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_865),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_865),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1137),
.Y(n_1361)
);

XOR2xp5_ASAP7_75t_L g1362 ( 
.A(n_1226),
.B(n_719),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_865),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1226),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1283),
.Y(n_1365)
);

INVxp67_ASAP7_75t_SL g1366 ( 
.A(n_793),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_876),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_876),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_876),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1283),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_882),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_882),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_739),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_745),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_746),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_882),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_747),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_909),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_909),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_909),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_760),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1164),
.B(n_721),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_748),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_750),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_977),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_806),
.B(n_0),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_926),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_977),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_751),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_977),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_752),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_760),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1001),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_756),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_758),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_759),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_862),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_764),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_765),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_935),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1011),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1001),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1051),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1255),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1001),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1232),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1262),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1232),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1232),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1293),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1257),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1302),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1257),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1257),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_793),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_793),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_766),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_767),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_769),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_793),
.Y(n_1420)
);

CKINVDCx14_ASAP7_75t_R g1421 ( 
.A(n_786),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_862),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_786),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_869),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_869),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_869),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_869),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_869),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_770),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_763),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_771),
.Y(n_1431)
);

CKINVDCx16_ASAP7_75t_R g1432 ( 
.A(n_761),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_869),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_927),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_927),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_761),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_795),
.Y(n_1437)
);

CKINVDCx14_ASAP7_75t_R g1438 ( 
.A(n_1125),
.Y(n_1438)
);

CKINVDCx16_ASAP7_75t_R g1439 ( 
.A(n_761),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_772),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_890),
.B(n_0),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_927),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_773),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_927),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_774),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_927),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_775),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_776),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_780),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_781),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_927),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_784),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_785),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_965),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_965),
.Y(n_1455)
);

CKINVDCx16_ASAP7_75t_R g1456 ( 
.A(n_761),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_789),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_965),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_808),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_791),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_818),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_843),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_965),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1164),
.B(n_4),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_965),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_965),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1004),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1004),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_792),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_880),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_794),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_800),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1004),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_802),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1004),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_790),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_804),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1004),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_953),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_805),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1004),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_809),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1079),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_810),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_813),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1079),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1079),
.Y(n_1487)
);

CKINVDCx14_ASAP7_75t_R g1488 ( 
.A(n_1125),
.Y(n_1488)
);

BUFx10_ASAP7_75t_L g1489 ( 
.A(n_890),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_815),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_817),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_986),
.B(n_2),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_986),
.B(n_4),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_819),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1079),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_820),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1036),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1079),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_823),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_824),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1079),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_825),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1050),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1074),
.Y(n_1504)
);

CKINVDCx12_ASAP7_75t_R g1505 ( 
.A(n_742),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_829),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1117),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_830),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1117),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1117),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1117),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1117),
.Y(n_1512)
);

NOR2xp67_ASAP7_75t_L g1513 ( 
.A(n_1074),
.B(n_5),
.Y(n_1513)
);

INVxp33_ASAP7_75t_L g1514 ( 
.A(n_1256),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_831),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1117),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_832),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1184),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1184),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1054),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1184),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1184),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_833),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_834),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_835),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1056),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1184),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1184),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1201),
.Y(n_1529)
);

BUFx10_ASAP7_75t_L g1530 ( 
.A(n_1256),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1201),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_836),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1201),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_839),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1201),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_841),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_842),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_846),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1201),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_847),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1201),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1250),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1250),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_851),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1066),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1250),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1250),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_852),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1250),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1250),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_740),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_740),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1279),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_742),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_856),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_859),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_860),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_861),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_863),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_864),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_741),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_741),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_790),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_866),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_754),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_870),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_754),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_872),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_755),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_873),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_874),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_877),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_755),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_757),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_878),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_879),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_1279),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_742),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_881),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_883),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_884),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_744),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_757),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_887),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_888),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_744),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_892),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_893),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_894),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_768),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_895),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_768),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_896),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_897),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_900),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1072),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_901),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_903),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_904),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_905),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_790),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1081),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_777),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1099),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_777),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_906),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_910),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_778),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_778),
.B(n_6),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_911),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_912),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_913),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_779),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1119),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_914),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1136),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_915),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_779),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_921),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_790),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_931),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_782),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_932),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_744),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_762),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_762),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_933),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_782),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_787),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_787),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_788),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_788),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_934),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_796),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1162),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_796),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_798),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_762),
.Y(n_1638)
);

CKINVDCx16_ASAP7_75t_R g1639 ( 
.A(n_797),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_798),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_940),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1186),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_803),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_803),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_941),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_807),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_942),
.Y(n_1647)
);

NOR2xp67_ASAP7_75t_L g1648 ( 
.A(n_1020),
.B(n_6),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_946),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_947),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_807),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_948),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_950),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_811),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_951),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_811),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_783),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_956),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1210),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_958),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_816),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1211),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_816),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1214),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_959),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_783),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_821),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_821),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_822),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_822),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_826),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_826),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_961),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_963),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_964),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_797),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_968),
.Y(n_1677)
);

BUFx5_ASAP7_75t_L g1678 ( 
.A(n_827),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_969),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_970),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_827),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_828),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_971),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_972),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_974),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1231),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_975),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_980),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_983),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_987),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_828),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_988),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_838),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_838),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_840),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_993),
.Y(n_1696)
);

NOR2xp67_ASAP7_75t_L g1697 ( 
.A(n_1020),
.B(n_7),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_840),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_845),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_845),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_853),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_995),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1238),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_996),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_853),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_857),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_997),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_797),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_999),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1000),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1003),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_857),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1006),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_783),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_868),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_868),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_871),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_1243),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_871),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1007),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_875),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1009),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1013),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1015),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1016),
.Y(n_1725)
);

BUFx10_ASAP7_75t_L g1726 ( 
.A(n_743),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_875),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1281),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1017),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_812),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_886),
.Y(n_1731)
);

CKINVDCx14_ASAP7_75t_R g1732 ( 
.A(n_797),
.Y(n_1732)
);

CKINVDCx14_ASAP7_75t_R g1733 ( 
.A(n_801),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1019),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1021),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_886),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1023),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1291),
.Y(n_1738)
);

CKINVDCx20_ASAP7_75t_R g1739 ( 
.A(n_1298),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_891),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1025),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1026),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1027),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_891),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1028),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1301),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_898),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1029),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1030),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_812),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_898),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_907),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_801),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_801),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_907),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_908),
.Y(n_1756)
);

CKINVDCx14_ASAP7_75t_R g1757 ( 
.A(n_801),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_812),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_908),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1031),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1037),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_917),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_917),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_918),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_918),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1040),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_920),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1042),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_920),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1043),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_922),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1045),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_837),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1046),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1052),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1726),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_1430),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1366),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1349),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1349),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1563),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1400),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1345),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1401),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1350),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1352),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_1437),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1459),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1353),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1467),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1467),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1563),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1403),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1416),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1415),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1404),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1420),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1425),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1426),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1427),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1407),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1710),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1345),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1433),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1435),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1442),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1444),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1446),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1451),
.Y(n_1809)
);

INVxp33_ASAP7_75t_L g1810 ( 
.A(n_1743),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1454),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1416),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1348),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1387),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1455),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1473),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1410),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1461),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1309),
.Y(n_1819)
);

CKINVDCx16_ASAP7_75t_R g1820 ( 
.A(n_1311),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1658),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1458),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1463),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1465),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1466),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1468),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1475),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_1462),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1478),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1601),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1481),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1483),
.Y(n_1832)
);

INVxp33_ASAP7_75t_SL g1833 ( 
.A(n_1310),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1486),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1601),
.Y(n_1835)
);

INVxp67_ASAP7_75t_SL g1836 ( 
.A(n_1620),
.Y(n_1836)
);

CKINVDCx16_ASAP7_75t_R g1837 ( 
.A(n_1326),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1487),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1501),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1310),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1470),
.Y(n_1841)
);

CKINVDCx20_ASAP7_75t_R g1842 ( 
.A(n_1479),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1507),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1509),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1770),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1510),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1511),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1512),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1516),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1775),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1519),
.Y(n_1851)
);

INVxp33_ASAP7_75t_SL g1852 ( 
.A(n_1315),
.Y(n_1852)
);

INVxp67_ASAP7_75t_SL g1853 ( 
.A(n_1620),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1521),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1412),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1522),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1417),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1418),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1473),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1527),
.Y(n_1860)
);

CKINVDCx20_ASAP7_75t_R g1861 ( 
.A(n_1503),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1528),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1529),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1531),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1520),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1533),
.Y(n_1866)
);

INVxp67_ASAP7_75t_SL g1867 ( 
.A(n_1753),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1419),
.Y(n_1868)
);

CKINVDCx16_ASAP7_75t_R g1869 ( 
.A(n_1732),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1429),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1539),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1541),
.Y(n_1872)
);

CKINVDCx16_ASAP7_75t_R g1873 ( 
.A(n_1733),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1542),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1431),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1495),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1545),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1440),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1443),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1346),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1596),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1445),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1447),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1448),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1543),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1449),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1547),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1450),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1550),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1753),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1354),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1356),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1359),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1360),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1363),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1367),
.Y(n_1896)
);

INVxp33_ASAP7_75t_L g1897 ( 
.A(n_1330),
.Y(n_1897)
);

CKINVDCx20_ASAP7_75t_R g1898 ( 
.A(n_1602),
.Y(n_1898)
);

CKINVDCx16_ASAP7_75t_R g1899 ( 
.A(n_1757),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1368),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1452),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1369),
.Y(n_1902)
);

CKINVDCx20_ASAP7_75t_R g1903 ( 
.A(n_1604),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1614),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1371),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1754),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1372),
.Y(n_1907)
);

INVxp33_ASAP7_75t_SL g1908 ( 
.A(n_1315),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1453),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1457),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1460),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1376),
.Y(n_1912)
);

CKINVDCx16_ASAP7_75t_R g1913 ( 
.A(n_1432),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_SL g1914 ( 
.A(n_1321),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1378),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1379),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1495),
.Y(n_1917)
);

INVxp33_ASAP7_75t_SL g1918 ( 
.A(n_1317),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1380),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1385),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1616),
.Y(n_1921)
);

CKINVDCx20_ASAP7_75t_R g1922 ( 
.A(n_1635),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1659),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1388),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_1662),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1754),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1390),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1346),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1393),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1436),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1402),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1351),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1469),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1351),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1703),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1405),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1471),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1406),
.Y(n_1938)
);

INVxp33_ASAP7_75t_SL g1939 ( 
.A(n_1317),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1436),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1355),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1408),
.Y(n_1942)
);

CKINVDCx16_ASAP7_75t_R g1943 ( 
.A(n_1439),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1472),
.Y(n_1944)
);

CKINVDCx20_ASAP7_75t_R g1945 ( 
.A(n_1718),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1411),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1474),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1355),
.Y(n_1948)
);

CKINVDCx20_ASAP7_75t_R g1949 ( 
.A(n_1728),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1476),
.Y(n_1950)
);

INVxp67_ASAP7_75t_SL g1951 ( 
.A(n_1332),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1477),
.Y(n_1952)
);

CKINVDCx16_ASAP7_75t_R g1953 ( 
.A(n_1456),
.Y(n_1953)
);

CKINVDCx20_ASAP7_75t_R g1954 ( 
.A(n_1738),
.Y(n_1954)
);

INVxp67_ASAP7_75t_SL g1955 ( 
.A(n_1332),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1498),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1413),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1414),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1549),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_1739),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1549),
.Y(n_1961)
);

BUFx3_ASAP7_75t_L g1962 ( 
.A(n_1409),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1357),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1480),
.Y(n_1964)
);

INVxp67_ASAP7_75t_SL g1965 ( 
.A(n_1409),
.Y(n_1965)
);

INVxp67_ASAP7_75t_SL g1966 ( 
.A(n_1434),
.Y(n_1966)
);

CKINVDCx20_ASAP7_75t_R g1967 ( 
.A(n_1746),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1303),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1482),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1304),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1484),
.Y(n_1971)
);

CKINVDCx16_ASAP7_75t_R g1972 ( 
.A(n_1639),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1304),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1304),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1304),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1434),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1434),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1304),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_1421),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1485),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1305),
.Y(n_1981)
);

CKINVDCx16_ASAP7_75t_R g1982 ( 
.A(n_1438),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1307),
.Y(n_1983)
);

CKINVDCx16_ASAP7_75t_R g1984 ( 
.A(n_1488),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1308),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1320),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1314),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1496),
.Y(n_1988)
);

INVxp67_ASAP7_75t_SL g1989 ( 
.A(n_1320),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1316),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1322),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1324),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1329),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1357),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_1358),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1476),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1334),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1499),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1336),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1337),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1338),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1339),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1320),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1340),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1342),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1344),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1358),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1320),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1500),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1502),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1361),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1506),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1347),
.Y(n_2013)
);

INVxp67_ASAP7_75t_SL g2014 ( 
.A(n_1320),
.Y(n_2014)
);

BUFx10_ASAP7_75t_L g2015 ( 
.A(n_1306),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1498),
.Y(n_2016)
);

BUFx10_ASAP7_75t_L g2017 ( 
.A(n_1306),
.Y(n_2017)
);

CKINVDCx20_ASAP7_75t_R g2018 ( 
.A(n_1361),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1343),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1535),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_1364),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1676),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1535),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1546),
.Y(n_2024)
);

CKINVDCx16_ASAP7_75t_R g2025 ( 
.A(n_1497),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1546),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1551),
.Y(n_2027)
);

INVxp67_ASAP7_75t_L g2028 ( 
.A(n_1676),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1552),
.Y(n_2029)
);

CKINVDCx16_ASAP7_75t_R g2030 ( 
.A(n_1526),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1364),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1365),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1561),
.Y(n_2033)
);

HB1xp67_ASAP7_75t_L g2034 ( 
.A(n_1365),
.Y(n_2034)
);

CKINVDCx20_ASAP7_75t_R g2035 ( 
.A(n_1370),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1508),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1562),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1565),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1567),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1515),
.Y(n_2040)
);

CKINVDCx20_ASAP7_75t_R g2041 ( 
.A(n_1370),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1642),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1517),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1343),
.Y(n_2044)
);

INVxp67_ASAP7_75t_SL g2045 ( 
.A(n_1343),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1569),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1573),
.Y(n_2047)
);

INVxp33_ASAP7_75t_SL g2048 ( 
.A(n_1318),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1574),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1583),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1523),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1664),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1524),
.Y(n_2053)
);

CKINVDCx14_ASAP7_75t_R g2054 ( 
.A(n_1318),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1590),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1592),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1525),
.Y(n_2057)
);

INVxp67_ASAP7_75t_SL g2058 ( 
.A(n_1343),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1603),
.Y(n_2059)
);

INVxp33_ASAP7_75t_L g2060 ( 
.A(n_1397),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1532),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1534),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1536),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1343),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1537),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1605),
.Y(n_2066)
);

INVxp67_ASAP7_75t_L g2067 ( 
.A(n_1708),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1608),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1613),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1618),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1622),
.Y(n_2071)
);

INVxp33_ASAP7_75t_L g2072 ( 
.A(n_1514),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1538),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1540),
.Y(n_2074)
);

INVxp67_ASAP7_75t_SL g2075 ( 
.A(n_1424),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1628),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1629),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1630),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1544),
.Y(n_2079)
);

INVxp67_ASAP7_75t_SL g2080 ( 
.A(n_1424),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1631),
.Y(n_2081)
);

INVxp67_ASAP7_75t_SL g2082 ( 
.A(n_1424),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1632),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1548),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1686),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1634),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1636),
.Y(n_2087)
);

CKINVDCx20_ASAP7_75t_R g2088 ( 
.A(n_1319),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_1319),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1555),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1424),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1637),
.Y(n_2092)
);

CKINVDCx20_ASAP7_75t_R g2093 ( 
.A(n_1323),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1640),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_1323),
.Y(n_2095)
);

CKINVDCx20_ASAP7_75t_R g2096 ( 
.A(n_1325),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1424),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1643),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1644),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1556),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1428),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1646),
.Y(n_2102)
);

CKINVDCx16_ASAP7_75t_R g2103 ( 
.A(n_1321),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1428),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1651),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1654),
.Y(n_2106)
);

CKINVDCx20_ASAP7_75t_R g2107 ( 
.A(n_1325),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1557),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1428),
.Y(n_2109)
);

INVxp67_ASAP7_75t_SL g2110 ( 
.A(n_1428),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1656),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1428),
.Y(n_2112)
);

CKINVDCx20_ASAP7_75t_R g2113 ( 
.A(n_1328),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1661),
.Y(n_2114)
);

INVxp33_ASAP7_75t_SL g2115 ( 
.A(n_1328),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1663),
.Y(n_2116)
);

INVxp67_ASAP7_75t_SL g2117 ( 
.A(n_1518),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1667),
.Y(n_2118)
);

CKINVDCx16_ASAP7_75t_R g2119 ( 
.A(n_1321),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1558),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1668),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_1559),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1669),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1670),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1671),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1672),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1518),
.Y(n_2127)
);

CKINVDCx20_ASAP7_75t_R g2128 ( 
.A(n_1331),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_1560),
.Y(n_2129)
);

INVxp67_ASAP7_75t_L g2130 ( 
.A(n_1708),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1681),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1564),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1682),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1566),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1691),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1518),
.Y(n_2136)
);

INVxp67_ASAP7_75t_SL g2137 ( 
.A(n_1518),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1568),
.Y(n_2138)
);

INVxp67_ASAP7_75t_SL g2139 ( 
.A(n_1518),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1693),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1694),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1570),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1695),
.Y(n_2143)
);

INVxp67_ASAP7_75t_L g2144 ( 
.A(n_1381),
.Y(n_2144)
);

CKINVDCx20_ASAP7_75t_R g2145 ( 
.A(n_1331),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1698),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1582),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1699),
.Y(n_2148)
);

CKINVDCx20_ASAP7_75t_R g2149 ( 
.A(n_1333),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1700),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1571),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1701),
.Y(n_2152)
);

CKINVDCx14_ASAP7_75t_R g2153 ( 
.A(n_1333),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1705),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1706),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1712),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1715),
.Y(n_2157)
);

INVxp67_ASAP7_75t_L g2158 ( 
.A(n_1392),
.Y(n_2158)
);

INVxp67_ASAP7_75t_SL g2159 ( 
.A(n_1422),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1572),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1582),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1575),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1716),
.Y(n_2163)
);

INVxp67_ASAP7_75t_SL g2164 ( 
.A(n_1504),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1794),
.Y(n_2165)
);

AND2x6_ASAP7_75t_L g2166 ( 
.A(n_1981),
.B(n_837),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1790),
.Y(n_2167)
);

BUFx6f_ASAP7_75t_L g2168 ( 
.A(n_2064),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_1790),
.B(n_1791),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1951),
.B(n_1576),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1794),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1812),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1776),
.B(n_1579),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1791),
.B(n_1554),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_2064),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_2064),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_1959),
.A2(n_1313),
.B(n_1312),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_2158),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1955),
.B(n_1580),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1977),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1802),
.A2(n_1581),
.B1(n_1585),
.B2(n_1584),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_1961),
.B(n_1554),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1812),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1891),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_1977),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_1962),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_2003),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1892),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_2147),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1965),
.B(n_1966),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1976),
.B(n_1587),
.Y(n_2191)
);

BUFx12f_ASAP7_75t_L g2192 ( 
.A(n_2015),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1813),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1814),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_1962),
.B(n_1578),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_2161),
.A2(n_1313),
.B(n_1312),
.Y(n_2196)
);

BUFx12f_ASAP7_75t_L g2197 ( 
.A(n_2015),
.Y(n_2197)
);

BUFx3_ASAP7_75t_L g2198 ( 
.A(n_2147),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1816),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_2003),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1816),
.Y(n_2201)
);

CKINVDCx16_ASAP7_75t_R g2202 ( 
.A(n_1982),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_R g2203 ( 
.A1(n_1845),
.A2(n_1362),
.B1(n_1057),
.B2(n_1058),
.Y(n_2203)
);

OAI21x1_ASAP7_75t_L g2204 ( 
.A1(n_2161),
.A2(n_1327),
.B(n_1773),
.Y(n_2204)
);

INVx5_ASAP7_75t_L g2205 ( 
.A(n_2003),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2101),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1859),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1785),
.B(n_1578),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1859),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1893),
.B(n_1624),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_2072),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1778),
.B(n_1588),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_2101),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1983),
.B(n_1985),
.Y(n_2214)
);

CKINVDCx6p67_ASAP7_75t_R g2215 ( 
.A(n_1869),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1876),
.Y(n_2216)
);

INVx6_ASAP7_75t_L g2217 ( 
.A(n_1873),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_SL g2218 ( 
.A1(n_2042),
.A2(n_1423),
.B1(n_1049),
.B2(n_1274),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1817),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1876),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1917),
.Y(n_2221)
);

INVx5_ASAP7_75t_L g2222 ( 
.A(n_2101),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1894),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1895),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1917),
.Y(n_2225)
);

CKINVDCx6p67_ASAP7_75t_R g2226 ( 
.A(n_1899),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1786),
.B(n_1624),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1956),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1817),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1821),
.A2(n_1589),
.B1(n_1593),
.B2(n_1591),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1956),
.Y(n_2231)
);

INVx4_ASAP7_75t_L g2232 ( 
.A(n_2044),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1896),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2044),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_2091),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1900),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1789),
.B(n_1625),
.Y(n_2237)
);

CKINVDCx6p67_ASAP7_75t_R g2238 ( 
.A(n_1984),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2016),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1902),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_2091),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_2025),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2159),
.A2(n_1382),
.B1(n_1464),
.B2(n_1492),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2020),
.Y(n_2244)
);

OA21x2_ASAP7_75t_L g2245 ( 
.A1(n_1987),
.A2(n_1327),
.B(n_1625),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_1905),
.B(n_1657),
.Y(n_2246)
);

AND2x6_ASAP7_75t_L g2247 ( 
.A(n_1990),
.B(n_837),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2164),
.A2(n_1594),
.B1(n_1597),
.B2(n_1595),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1907),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_2030),
.Y(n_2250)
);

BUFx6f_ASAP7_75t_L g2251 ( 
.A(n_2097),
.Y(n_2251)
);

CKINVDCx8_ASAP7_75t_R g2252 ( 
.A(n_1837),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_1912),
.B(n_1657),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2072),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1915),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1991),
.B(n_1598),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1992),
.B(n_1599),
.Y(n_2257)
);

INVx4_ASAP7_75t_L g2258 ( 
.A(n_2097),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2023),
.Y(n_2259)
);

BUFx8_ASAP7_75t_L g2260 ( 
.A(n_1914),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_2104),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_1782),
.A2(n_1600),
.B1(n_1607),
.B2(n_1606),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2024),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_1845),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2026),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_1916),
.B(n_1666),
.Y(n_2266)
);

OA21x2_ASAP7_75t_L g2267 ( 
.A1(n_1993),
.A2(n_1714),
.B(n_1666),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_1997),
.Y(n_2268)
);

OAI22xp5_ASAP7_75t_SL g2269 ( 
.A1(n_2042),
.A2(n_849),
.B1(n_928),
.B2(n_867),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1795),
.Y(n_2270)
);

INVx5_ASAP7_75t_L g2271 ( 
.A(n_2109),
.Y(n_2271)
);

AND2x2_ASAP7_75t_SL g2272 ( 
.A(n_2051),
.B(n_1609),
.Y(n_2272)
);

OAI21x1_ASAP7_75t_L g2273 ( 
.A1(n_2109),
.A2(n_1773),
.B(n_1730),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1919),
.Y(n_2274)
);

INVx5_ASAP7_75t_L g2275 ( 
.A(n_2112),
.Y(n_2275)
);

INVx6_ASAP7_75t_L g2276 ( 
.A(n_1986),
.Y(n_2276)
);

BUFx6f_ASAP7_75t_L g2277 ( 
.A(n_2127),
.Y(n_2277)
);

AND2x6_ASAP7_75t_L g2278 ( 
.A(n_1999),
.B(n_848),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_2127),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2136),
.A2(n_1730),
.B(n_1714),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2000),
.B(n_1610),
.Y(n_2281)
);

BUFx12f_ASAP7_75t_L g2282 ( 
.A(n_2015),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_1783),
.Y(n_2283)
);

BUFx12f_ASAP7_75t_L g2284 ( 
.A(n_2017),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1920),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_2052),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1924),
.Y(n_2287)
);

BUFx8_ASAP7_75t_L g2288 ( 
.A(n_1914),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1797),
.Y(n_2289)
);

CKINVDCx6p67_ASAP7_75t_R g2290 ( 
.A(n_1979),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1927),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1798),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2052),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2001),
.B(n_1611),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1799),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1850),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_1776),
.Y(n_2297)
);

OAI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_1930),
.A2(n_1341),
.B1(n_1441),
.B2(n_1386),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_1970),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1973),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_1784),
.A2(n_1612),
.B1(n_1341),
.B2(n_1374),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_2085),
.Y(n_2302)
);

AND2x2_ASAP7_75t_SL g2303 ( 
.A(n_2057),
.B(n_848),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2002),
.B(n_1373),
.Y(n_2304)
);

BUFx6f_ASAP7_75t_L g2305 ( 
.A(n_1974),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_1929),
.B(n_1750),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2144),
.B(n_1553),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_1931),
.B(n_1750),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1850),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1800),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1936),
.Y(n_2311)
);

INVx5_ASAP7_75t_L g2312 ( 
.A(n_1989),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1968),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_1938),
.B(n_1942),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2085),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1946),
.B(n_1717),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1804),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1957),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_1975),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1805),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_1958),
.B(n_1719),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2004),
.B(n_1373),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_1940),
.A2(n_1513),
.B1(n_1493),
.B2(n_1375),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_2005),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_1793),
.A2(n_1375),
.B1(n_1377),
.B2(n_1374),
.Y(n_2325)
);

AND2x6_ASAP7_75t_L g2326 ( 
.A(n_2006),
.B(n_848),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_1950),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_1978),
.Y(n_2328)
);

INVx2_ASAP7_75t_SL g2329 ( 
.A(n_1803),
.Y(n_2329)
);

BUFx3_ASAP7_75t_L g2330 ( 
.A(n_2013),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_1796),
.A2(n_1383),
.B1(n_1384),
.B2(n_1377),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_1806),
.Y(n_2332)
);

OAI22x1_ASAP7_75t_R g2333 ( 
.A1(n_1777),
.A2(n_1774),
.B1(n_1384),
.B2(n_1389),
.Y(n_2333)
);

BUFx3_ASAP7_75t_L g2334 ( 
.A(n_2027),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2029),
.Y(n_2335)
);

INVx4_ASAP7_75t_L g2336 ( 
.A(n_1807),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1808),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1809),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1811),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2033),
.B(n_1721),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2037),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_1815),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_1822),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1823),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_1824),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2038),
.Y(n_2346)
);

BUFx8_ASAP7_75t_L g2347 ( 
.A(n_1914),
.Y(n_2347)
);

CKINVDCx11_ASAP7_75t_R g2348 ( 
.A(n_2017),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2039),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2046),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_1996),
.B(n_1383),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2047),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1825),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1826),
.Y(n_2354)
);

BUFx8_ASAP7_75t_SL g2355 ( 
.A(n_1777),
.Y(n_2355)
);

CKINVDCx11_ASAP7_75t_R g2356 ( 
.A(n_2017),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_1827),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_1829),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2022),
.B(n_1389),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2049),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1831),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1832),
.Y(n_2362)
);

BUFx12f_ASAP7_75t_L g2363 ( 
.A(n_1840),
.Y(n_2363)
);

CKINVDCx6p67_ASAP7_75t_R g2364 ( 
.A(n_1979),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2008),
.B(n_1391),
.Y(n_2365)
);

BUFx6f_ASAP7_75t_L g2366 ( 
.A(n_1834),
.Y(n_2366)
);

OA21x2_ASAP7_75t_L g2367 ( 
.A1(n_1838),
.A2(n_1763),
.B(n_1762),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1839),
.Y(n_2368)
);

OA21x2_ASAP7_75t_L g2369 ( 
.A1(n_1843),
.A2(n_1765),
.B(n_1764),
.Y(n_2369)
);

OAI22x1_ASAP7_75t_R g2370 ( 
.A1(n_1787),
.A2(n_1761),
.B1(n_1766),
.B2(n_1760),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_1844),
.Y(n_2371)
);

INVx6_ASAP7_75t_L g2372 ( 
.A(n_2014),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1846),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2050),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1847),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2055),
.B(n_1727),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2056),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2059),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2019),
.B(n_1391),
.Y(n_2379)
);

AND2x6_ASAP7_75t_L g2380 ( 
.A(n_2095),
.B(n_885),
.Y(n_2380)
);

INVxp33_ASAP7_75t_SL g2381 ( 
.A(n_1840),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_2028),
.B(n_1394),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_1848),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1849),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2067),
.B(n_1394),
.Y(n_2385)
);

OA21x2_ASAP7_75t_L g2386 ( 
.A1(n_1851),
.A2(n_1769),
.B(n_1767),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_1854),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2066),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_SL g2389 ( 
.A1(n_1994),
.A2(n_849),
.B1(n_928),
.B2(n_867),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_1856),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2068),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_1860),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_1862),
.Y(n_2393)
);

HB1xp67_ASAP7_75t_L g2394 ( 
.A(n_2130),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_1819),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1810),
.B(n_1395),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2069),
.B(n_1731),
.Y(n_2397)
);

INVx2_ASAP7_75t_SL g2398 ( 
.A(n_1880),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2070),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2071),
.B(n_1726),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1863),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2076),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_1830),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2077),
.Y(n_2404)
);

OA21x2_ASAP7_75t_L g2405 ( 
.A1(n_1864),
.A2(n_1740),
.B(n_1736),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2078),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2081),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_1866),
.Y(n_2408)
);

BUFx3_ASAP7_75t_L g2409 ( 
.A(n_2083),
.Y(n_2409)
);

BUFx2_ASAP7_75t_L g2410 ( 
.A(n_1994),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_1871),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_1872),
.Y(n_2412)
);

BUFx6f_ASAP7_75t_L g2413 ( 
.A(n_1874),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1885),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_1887),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_1835),
.Y(n_2416)
);

XOR2xp5_ASAP7_75t_L g2417 ( 
.A(n_1787),
.B(n_1395),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2086),
.B(n_1744),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_1810),
.B(n_1396),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1889),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2087),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2092),
.B(n_2094),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_1779),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_2098),
.Y(n_2424)
);

INVx3_ASAP7_75t_L g2425 ( 
.A(n_1780),
.Y(n_2425)
);

AND2x6_ASAP7_75t_L g2426 ( 
.A(n_2099),
.B(n_885),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2102),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_1890),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_2105),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2106),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_1995),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2111),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2114),
.Y(n_2433)
);

AOI22x1_ASAP7_75t_SL g2434 ( 
.A1(n_1819),
.A2(n_990),
.B1(n_998),
.B2(n_930),
.Y(n_2434)
);

CKINVDCx16_ASAP7_75t_R g2435 ( 
.A(n_1913),
.Y(n_2435)
);

OAI21x1_ASAP7_75t_L g2436 ( 
.A1(n_2045),
.A2(n_889),
.B(n_885),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2116),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2118),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_SL g2439 ( 
.A1(n_1995),
.A2(n_990),
.B1(n_998),
.B2(n_930),
.Y(n_2439)
);

OAI22xp5_ASAP7_75t_SL g2440 ( 
.A1(n_2011),
.A2(n_1049),
.B1(n_1085),
.B2(n_1035),
.Y(n_2440)
);

BUFx8_ASAP7_75t_L g2441 ( 
.A(n_2163),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2121),
.B(n_1747),
.Y(n_2442)
);

INVx4_ASAP7_75t_L g2443 ( 
.A(n_1801),
.Y(n_2443)
);

HB1xp67_ASAP7_75t_L g2444 ( 
.A(n_1906),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2123),
.Y(n_2445)
);

BUFx2_ASAP7_75t_L g2446 ( 
.A(n_2011),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2124),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_2125),
.Y(n_2448)
);

BUFx6f_ASAP7_75t_L g2449 ( 
.A(n_2126),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_2018),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2131),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_2133),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2135),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2140),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2141),
.Y(n_2455)
);

AOI22xp5_ASAP7_75t_L g2456 ( 
.A1(n_2162),
.A2(n_1398),
.B1(n_1399),
.B2(n_1396),
.Y(n_2456)
);

INVx5_ASAP7_75t_L g2457 ( 
.A(n_2058),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2075),
.B(n_1398),
.Y(n_2458)
);

BUFx12f_ASAP7_75t_L g2459 ( 
.A(n_1901),
.Y(n_2459)
);

BUFx3_ASAP7_75t_L g2460 ( 
.A(n_2143),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_1781),
.B(n_1399),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2146),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2148),
.Y(n_2463)
);

NOR2x1_ASAP7_75t_L g2464 ( 
.A(n_2150),
.B(n_1648),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2152),
.B(n_1726),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_2154),
.Y(n_2466)
);

OA21x2_ASAP7_75t_L g2467 ( 
.A1(n_2080),
.A2(n_1752),
.B(n_1751),
.Y(n_2467)
);

OAI22xp5_ASAP7_75t_R g2468 ( 
.A1(n_1901),
.A2(n_1059),
.B1(n_1060),
.B2(n_1053),
.Y(n_2468)
);

CKINVDCx6p67_ASAP7_75t_R g2469 ( 
.A(n_1943),
.Y(n_2469)
);

AND2x4_ASAP7_75t_L g2470 ( 
.A(n_2155),
.B(n_1755),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2156),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2157),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_1792),
.B(n_1756),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2082),
.Y(n_2474)
);

BUFx8_ASAP7_75t_SL g2475 ( 
.A(n_1788),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2110),
.Y(n_2476)
);

OA21x2_ASAP7_75t_L g2477 ( 
.A1(n_2117),
.A2(n_1771),
.B(n_1759),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2137),
.B(n_1490),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2139),
.Y(n_2479)
);

OA21x2_ASAP7_75t_L g2480 ( 
.A1(n_1836),
.A2(n_916),
.B(n_889),
.Y(n_2480)
);

CKINVDCx11_ASAP7_75t_R g2481 ( 
.A(n_1788),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_2054),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_1853),
.B(n_889),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1867),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_1926),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1855),
.B(n_1490),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_1857),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_1858),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_1928),
.B(n_916),
.Y(n_2489)
);

INVx3_ASAP7_75t_L g2490 ( 
.A(n_1868),
.Y(n_2490)
);

INVx5_ASAP7_75t_L g2491 ( 
.A(n_1953),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1870),
.B(n_1491),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_1875),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1932),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_1878),
.Y(n_2495)
);

BUFx12f_ASAP7_75t_L g2496 ( 
.A(n_1980),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_1879),
.B(n_1491),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_1882),
.B(n_1494),
.Y(n_2498)
);

OAI21x1_ASAP7_75t_L g2499 ( 
.A1(n_1934),
.A2(n_952),
.B(n_916),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1941),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_1883),
.Y(n_2501)
);

CKINVDCx8_ASAP7_75t_R g2502 ( 
.A(n_1972),
.Y(n_2502)
);

AOI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_1852),
.A2(n_1615),
.B1(n_1617),
.B2(n_1494),
.Y(n_2503)
);

BUFx8_ASAP7_75t_SL g2504 ( 
.A(n_1818),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_1897),
.B(n_1678),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_1948),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_1884),
.Y(n_2507)
);

INVxp67_ASAP7_75t_L g2508 ( 
.A(n_1963),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_1886),
.B(n_1615),
.Y(n_2509)
);

BUFx12f_ASAP7_75t_L g2510 ( 
.A(n_1980),
.Y(n_2510)
);

BUFx6f_ASAP7_75t_L g2511 ( 
.A(n_1888),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2007),
.B(n_952),
.Y(n_2512)
);

INVx4_ASAP7_75t_L g2513 ( 
.A(n_1909),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_1910),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2032),
.Y(n_2515)
);

AND2x2_ASAP7_75t_SL g2516 ( 
.A(n_2034),
.B(n_952),
.Y(n_2516)
);

INVxp67_ASAP7_75t_L g2517 ( 
.A(n_1988),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_1911),
.Y(n_2518)
);

OAI22x1_ASAP7_75t_R g2519 ( 
.A1(n_1818),
.A2(n_1774),
.B1(n_1619),
.B2(n_1621),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_1933),
.Y(n_2520)
);

BUFx2_ASAP7_75t_L g2521 ( 
.A(n_2018),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_1937),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_1944),
.Y(n_2523)
);

OA21x2_ASAP7_75t_L g2524 ( 
.A1(n_1947),
.A2(n_982),
.B(n_979),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_1952),
.B(n_979),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1964),
.Y(n_2526)
);

OA21x2_ASAP7_75t_L g2527 ( 
.A1(n_1969),
.A2(n_982),
.B(n_979),
.Y(n_2527)
);

INVxp67_ASAP7_75t_L g2528 ( 
.A(n_1988),
.Y(n_2528)
);

AND2x4_ASAP7_75t_L g2529 ( 
.A(n_1971),
.B(n_982),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2073),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2160),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2074),
.B(n_1617),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2079),
.Y(n_2533)
);

HB1xp67_ASAP7_75t_L g2534 ( 
.A(n_1897),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2084),
.Y(n_2535)
);

AND2x4_ASAP7_75t_L g2536 ( 
.A(n_2090),
.B(n_994),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2100),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2060),
.B(n_1678),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2108),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2120),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2122),
.Y(n_2541)
);

BUFx3_ASAP7_75t_L g2542 ( 
.A(n_2129),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2132),
.B(n_994),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2134),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2138),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2142),
.Y(n_2546)
);

OAI22xp5_ASAP7_75t_SL g2547 ( 
.A1(n_2021),
.A2(n_1085),
.B1(n_1102),
.B2(n_1035),
.Y(n_2547)
);

BUFx2_ASAP7_75t_L g2548 ( 
.A(n_2021),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_1852),
.A2(n_1619),
.B1(n_1623),
.B2(n_1621),
.Y(n_2549)
);

BUFx6f_ASAP7_75t_L g2550 ( 
.A(n_2151),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_1998),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_1998),
.Y(n_2552)
);

OAI21x1_ASAP7_75t_L g2553 ( 
.A1(n_2153),
.A2(n_1034),
.B(n_994),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_2009),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2009),
.Y(n_2555)
);

INVx6_ASAP7_75t_L g2556 ( 
.A(n_1820),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2010),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2060),
.Y(n_2558)
);

OA21x2_ASAP7_75t_L g2559 ( 
.A1(n_2010),
.A2(n_1039),
.B(n_1034),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2012),
.B(n_1623),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2031),
.Y(n_2561)
);

CKINVDCx16_ASAP7_75t_R g2562 ( 
.A(n_2103),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2012),
.B(n_1678),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_1908),
.A2(n_1627),
.B1(n_1641),
.B2(n_1633),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_L g2565 ( 
.A(n_2036),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_1908),
.A2(n_1627),
.B1(n_1641),
.B2(n_1633),
.Y(n_2566)
);

INVxp67_ASAP7_75t_L g2567 ( 
.A(n_2036),
.Y(n_2567)
);

INVx4_ASAP7_75t_L g2568 ( 
.A(n_2040),
.Y(n_2568)
);

INVx5_ASAP7_75t_L g2569 ( 
.A(n_2119),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2040),
.Y(n_2570)
);

OAI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_1918),
.A2(n_1647),
.B1(n_1649),
.B2(n_1645),
.Y(n_2571)
);

OA21x2_ASAP7_75t_L g2572 ( 
.A1(n_2043),
.A2(n_1039),
.B(n_1034),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_1918),
.B(n_1645),
.Y(n_2573)
);

HB1xp67_ASAP7_75t_L g2574 ( 
.A(n_2043),
.Y(n_2574)
);

OA21x2_ASAP7_75t_L g2575 ( 
.A1(n_2053),
.A2(n_1067),
.B(n_1039),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2053),
.B(n_1647),
.Y(n_2576)
);

HB1xp67_ASAP7_75t_L g2577 ( 
.A(n_2061),
.Y(n_2577)
);

INVx4_ASAP7_75t_L g2578 ( 
.A(n_2061),
.Y(n_2578)
);

BUFx2_ASAP7_75t_L g2579 ( 
.A(n_2031),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2062),
.B(n_1067),
.Y(n_2580)
);

INVx2_ASAP7_75t_SL g2581 ( 
.A(n_2062),
.Y(n_2581)
);

INVx3_ASAP7_75t_L g2582 ( 
.A(n_2063),
.Y(n_2582)
);

AND2x2_ASAP7_75t_SL g2583 ( 
.A(n_1939),
.B(n_1067),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2063),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2065),
.Y(n_2585)
);

OAI21x1_ASAP7_75t_L g2586 ( 
.A1(n_1939),
.A2(n_1098),
.B(n_1073),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2048),
.A2(n_1649),
.B1(n_1652),
.B2(n_1650),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2065),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2048),
.B(n_1650),
.Y(n_2589)
);

INVx5_ASAP7_75t_L g2590 ( 
.A(n_2115),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_1828),
.Y(n_2591)
);

BUFx6f_ASAP7_75t_L g2592 ( 
.A(n_2115),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_1833),
.B(n_1652),
.Y(n_2593)
);

BUFx6f_ASAP7_75t_L g2594 ( 
.A(n_1833),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2088),
.B(n_1653),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2088),
.B(n_1653),
.Y(n_2596)
);

OAI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2089),
.A2(n_1660),
.B1(n_1665),
.B2(n_1655),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2089),
.B(n_1073),
.Y(n_2598)
);

BUFx6f_ASAP7_75t_L g2599 ( 
.A(n_2149),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2093),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2093),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_2096),
.B(n_1655),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2096),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2107),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2107),
.B(n_1660),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_2113),
.Y(n_2606)
);

INVx6_ASAP7_75t_L g2607 ( 
.A(n_2113),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2128),
.B(n_1678),
.Y(n_2608)
);

CKINVDCx11_ASAP7_75t_R g2609 ( 
.A(n_1828),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2128),
.Y(n_2610)
);

INVx6_ASAP7_75t_L g2611 ( 
.A(n_2145),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2174),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2355),
.Y(n_2613)
);

NOR2xp33_ASAP7_75t_R g2614 ( 
.A(n_2193),
.B(n_1841),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2355),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2174),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2178),
.B(n_1665),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_2180),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2267),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_2193),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2174),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2267),
.Y(n_2622)
);

INVx3_ASAP7_75t_L g2623 ( 
.A(n_2177),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2194),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2505),
.B(n_1673),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_2194),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_2475),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2180),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2212),
.B(n_1673),
.Y(n_2629)
);

CKINVDCx16_ASAP7_75t_R g2630 ( 
.A(n_2435),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2422),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2475),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2504),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2211),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2267),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2422),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2182),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2245),
.Y(n_2638)
);

INVx3_ASAP7_75t_L g2639 ( 
.A(n_2177),
.Y(n_2639)
);

CKINVDCx20_ASAP7_75t_R g2640 ( 
.A(n_2242),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2254),
.Y(n_2641)
);

AND2x4_ASAP7_75t_L g2642 ( 
.A(n_2169),
.B(n_1073),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_2504),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2245),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2245),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2273),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2182),
.Y(n_2647)
);

NAND2xp33_ASAP7_75t_L g2648 ( 
.A(n_2166),
.B(n_1678),
.Y(n_2648)
);

NOR2xp67_ASAP7_75t_L g2649 ( 
.A(n_2491),
.B(n_1674),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_2481),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2481),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2273),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2609),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2505),
.B(n_1674),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2538),
.B(n_1675),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2396),
.B(n_2419),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2280),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2182),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2538),
.B(n_1675),
.Y(n_2659)
);

CKINVDCx20_ASAP7_75t_R g2660 ( 
.A(n_2242),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2609),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2427),
.Y(n_2662)
);

CKINVDCx5p33_ASAP7_75t_R g2663 ( 
.A(n_2250),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2427),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2534),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2430),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2280),
.Y(n_2667)
);

INVxp67_ASAP7_75t_L g2668 ( 
.A(n_2307),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2430),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2250),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2432),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_2459),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2563),
.B(n_1677),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2204),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2204),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2563),
.B(n_1677),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2432),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2433),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2459),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2496),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2196),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2433),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2438),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2438),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_2496),
.Y(n_2685)
);

OAI21x1_ASAP7_75t_L g2686 ( 
.A1(n_2436),
.A2(n_1108),
.B(n_1098),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2453),
.Y(n_2687)
);

BUFx8_ASAP7_75t_L g2688 ( 
.A(n_2286),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2315),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2510),
.Y(n_2690)
);

BUFx8_ASAP7_75t_L g2691 ( 
.A(n_2410),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2196),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2165),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_2510),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2453),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2462),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2293),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2462),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2471),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2471),
.Y(n_2700)
);

INVx1_ASAP7_75t_SL g2701 ( 
.A(n_2302),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2165),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2608),
.B(n_1679),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2472),
.Y(n_2704)
);

CKINVDCx5p33_ASAP7_75t_R g2705 ( 
.A(n_2348),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2171),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2348),
.Y(n_2707)
);

CKINVDCx5p33_ASAP7_75t_R g2708 ( 
.A(n_2356),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2171),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2472),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2195),
.Y(n_2711)
);

CKINVDCx20_ASAP7_75t_R g2712 ( 
.A(n_2591),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2195),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2356),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2195),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2341),
.Y(n_2716)
);

OR2x6_ASAP7_75t_L g2717 ( 
.A(n_2488),
.B(n_743),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2346),
.Y(n_2718)
);

CKINVDCx20_ASAP7_75t_R g2719 ( 
.A(n_2591),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2349),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_2180),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2350),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2180),
.Y(n_2723)
);

OA21x2_ASAP7_75t_L g2724 ( 
.A1(n_2436),
.A2(n_1680),
.B(n_1679),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_2395),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2352),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2360),
.Y(n_2727)
);

HB1xp67_ASAP7_75t_L g2728 ( 
.A(n_2558),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2374),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2377),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2378),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_L g2732 ( 
.A(n_2191),
.B(n_1680),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2180),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2395),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2186),
.B(n_1683),
.Y(n_2735)
);

CKINVDCx20_ASAP7_75t_R g2736 ( 
.A(n_2202),
.Y(n_2736)
);

OA21x2_ASAP7_75t_L g2737 ( 
.A1(n_2586),
.A2(n_1684),
.B(n_1683),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2172),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2388),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2391),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_2219),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2399),
.Y(n_2742)
);

BUFx2_ASAP7_75t_L g2743 ( 
.A(n_2608),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2525),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_2185),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2172),
.Y(n_2746)
);

CKINVDCx20_ASAP7_75t_R g2747 ( 
.A(n_2562),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2400),
.B(n_1684),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2219),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2183),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2402),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2404),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2229),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2307),
.Y(n_2754)
);

INVxp67_ASAP7_75t_L g2755 ( 
.A(n_2359),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2380),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2229),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2264),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2406),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2264),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2407),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_SL g2762 ( 
.A(n_2303),
.B(n_1685),
.Y(n_2762)
);

BUFx6f_ASAP7_75t_L g2763 ( 
.A(n_2185),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2421),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2525),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2437),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2296),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2400),
.B(n_2465),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2451),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2232),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2296),
.Y(n_2771)
);

AND2x6_ASAP7_75t_L g2772 ( 
.A(n_2484),
.B(n_2485),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2465),
.B(n_1685),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2184),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2188),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2232),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2223),
.Y(n_2777)
);

OA21x2_ASAP7_75t_L g2778 ( 
.A1(n_2586),
.A2(n_1688),
.B(n_1687),
.Y(n_2778)
);

CKINVDCx20_ASAP7_75t_R g2779 ( 
.A(n_2469),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2224),
.Y(n_2780)
);

CKINVDCx20_ASAP7_75t_R g2781 ( 
.A(n_2469),
.Y(n_2781)
);

CKINVDCx20_ASAP7_75t_R g2782 ( 
.A(n_2238),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_2238),
.Y(n_2783)
);

BUFx6f_ASAP7_75t_L g2784 ( 
.A(n_2185),
.Y(n_2784)
);

BUFx8_ASAP7_75t_L g2785 ( 
.A(n_2431),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2233),
.Y(n_2786)
);

CKINVDCx20_ASAP7_75t_R g2787 ( 
.A(n_2252),
.Y(n_2787)
);

INVx1_ASAP7_75t_SL g2788 ( 
.A(n_2446),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_2482),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2236),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2256),
.B(n_1687),
.Y(n_2791)
);

CKINVDCx5p33_ASAP7_75t_R g2792 ( 
.A(n_2482),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2183),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2186),
.B(n_1688),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2327),
.B(n_2394),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2240),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2199),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2249),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2255),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2274),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2285),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2199),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2525),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2185),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2287),
.Y(n_2805)
);

HB1xp67_ASAP7_75t_L g2806 ( 
.A(n_2529),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_2192),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2529),
.Y(n_2808)
);

CKINVDCx20_ASAP7_75t_R g2809 ( 
.A(n_2252),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2190),
.B(n_1689),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2201),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_2192),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2303),
.B(n_1689),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2169),
.B(n_1098),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2185),
.Y(n_2815)
);

CKINVDCx5p33_ASAP7_75t_R g2816 ( 
.A(n_2197),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2291),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2311),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2318),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2208),
.Y(n_2820)
);

BUFx6f_ASAP7_75t_L g2821 ( 
.A(n_2198),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_2197),
.Y(n_2822)
);

AND2x4_ASAP7_75t_L g2823 ( 
.A(n_2169),
.B(n_1108),
.Y(n_2823)
);

AND2x6_ASAP7_75t_L g2824 ( 
.A(n_2483),
.B(n_1108),
.Y(n_2824)
);

CKINVDCx16_ASAP7_75t_R g2825 ( 
.A(n_2333),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2282),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2208),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2227),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_2282),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2201),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2297),
.B(n_2329),
.Y(n_2831)
);

INVx1_ASAP7_75t_SL g2832 ( 
.A(n_2450),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2207),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2227),
.Y(n_2834)
);

OA21x2_ASAP7_75t_L g2835 ( 
.A1(n_2499),
.A2(n_1692),
.B(n_1690),
.Y(n_2835)
);

BUFx6f_ASAP7_75t_L g2836 ( 
.A(n_2198),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_2284),
.Y(n_2837)
);

CKINVDCx20_ASAP7_75t_R g2838 ( 
.A(n_2417),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2447),
.B(n_2476),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_R g2840 ( 
.A(n_2309),
.B(n_1841),
.Y(n_2840)
);

INVx3_ASAP7_75t_L g2841 ( 
.A(n_2232),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2284),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2529),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2207),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2516),
.B(n_2297),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_SL g2846 ( 
.A(n_2516),
.B(n_1690),
.Y(n_2846)
);

NOR2xp33_ASAP7_75t_R g2847 ( 
.A(n_2309),
.B(n_1842),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_2363),
.Y(n_2848)
);

AND2x6_ASAP7_75t_L g2849 ( 
.A(n_2483),
.B(n_1161),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2237),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2258),
.Y(n_2851)
);

CKINVDCx20_ASAP7_75t_R g2852 ( 
.A(n_2521),
.Y(n_2852)
);

CKINVDCx20_ASAP7_75t_R g2853 ( 
.A(n_2548),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2237),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2447),
.B(n_1692),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2209),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2447),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_2363),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2314),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2209),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2329),
.B(n_1696),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2314),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2314),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_2215),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2215),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2334),
.Y(n_2866)
);

CKINVDCx20_ASAP7_75t_R g2867 ( 
.A(n_2561),
.Y(n_2867)
);

OR2x2_ASAP7_75t_L g2868 ( 
.A(n_2580),
.B(n_1696),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2189),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2216),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2216),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2220),
.Y(n_2872)
);

CKINVDCx20_ASAP7_75t_R g2873 ( 
.A(n_2579),
.Y(n_2873)
);

NAND2x1p5_ASAP7_75t_L g2874 ( 
.A(n_2559),
.B(n_1582),
.Y(n_2874)
);

CKINVDCx20_ASAP7_75t_R g2875 ( 
.A(n_2290),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2334),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2536),
.B(n_1702),
.Y(n_2877)
);

CKINVDCx5p33_ASAP7_75t_R g2878 ( 
.A(n_2226),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2220),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2272),
.A2(n_1702),
.B1(n_1707),
.B2(n_1704),
.Y(n_2880)
);

BUFx2_ASAP7_75t_L g2881 ( 
.A(n_2380),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2335),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2398),
.B(n_1704),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2335),
.Y(n_2884)
);

NOR2xp67_ASAP7_75t_L g2885 ( 
.A(n_2491),
.B(n_1707),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2556),
.Y(n_2886)
);

BUFx6f_ASAP7_75t_L g2887 ( 
.A(n_2189),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2398),
.B(n_1709),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2226),
.Y(n_2889)
);

CKINVDCx5p33_ASAP7_75t_R g2890 ( 
.A(n_2290),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2409),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2409),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_2364),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2476),
.B(n_1709),
.Y(n_2894)
);

CKINVDCx5p33_ASAP7_75t_R g2895 ( 
.A(n_2487),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2479),
.B(n_1711),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2258),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2221),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2424),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2221),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2225),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2382),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2424),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2479),
.B(n_1711),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2487),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2515),
.B(n_1713),
.Y(n_2906)
);

CKINVDCx20_ASAP7_75t_R g2907 ( 
.A(n_2364),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2474),
.B(n_1713),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_2487),
.Y(n_2909)
);

CKINVDCx20_ASAP7_75t_R g2910 ( 
.A(n_2502),
.Y(n_2910)
);

INVx3_ASAP7_75t_L g2911 ( 
.A(n_2258),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2225),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2235),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2214),
.B(n_1720),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2429),
.Y(n_2915)
);

CKINVDCx5p33_ASAP7_75t_R g2916 ( 
.A(n_2487),
.Y(n_2916)
);

BUFx6f_ASAP7_75t_L g2917 ( 
.A(n_2189),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2488),
.Y(n_2918)
);

CKINVDCx5p33_ASAP7_75t_R g2919 ( 
.A(n_2488),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2429),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_2167),
.B(n_1161),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2488),
.Y(n_2922)
);

CKINVDCx20_ASAP7_75t_R g2923 ( 
.A(n_2502),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2460),
.Y(n_2924)
);

INVx3_ASAP7_75t_L g2925 ( 
.A(n_2235),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2228),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2473),
.B(n_1720),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2473),
.B(n_1722),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2473),
.B(n_1722),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2536),
.B(n_1723),
.Y(n_2930)
);

INVx3_ASAP7_75t_L g2931 ( 
.A(n_2235),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2228),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2460),
.Y(n_2933)
);

CKINVDCx20_ASAP7_75t_R g2934 ( 
.A(n_2370),
.Y(n_2934)
);

INVxp67_ASAP7_75t_SL g2935 ( 
.A(n_2168),
.Y(n_2935)
);

BUFx6f_ASAP7_75t_L g2936 ( 
.A(n_2313),
.Y(n_2936)
);

BUFx6f_ASAP7_75t_L g2937 ( 
.A(n_2313),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2235),
.Y(n_2938)
);

CKINVDCx20_ASAP7_75t_R g2939 ( 
.A(n_2519),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2515),
.B(n_2385),
.Y(n_2940)
);

BUFx6f_ASAP7_75t_L g2941 ( 
.A(n_2313),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2210),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2210),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2210),
.Y(n_2944)
);

BUFx2_ASAP7_75t_L g2945 ( 
.A(n_2380),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2246),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2231),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2246),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2246),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2253),
.Y(n_2950)
);

CKINVDCx20_ASAP7_75t_R g2951 ( 
.A(n_2607),
.Y(n_2951)
);

BUFx6f_ASAP7_75t_L g2952 ( 
.A(n_2313),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2403),
.B(n_1723),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2483),
.B(n_1724),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2253),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2253),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_R g2957 ( 
.A(n_2582),
.B(n_1842),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2266),
.Y(n_2958)
);

CKINVDCx20_ASAP7_75t_R g2959 ( 
.A(n_2607),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_2488),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_2495),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2268),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2266),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2266),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2268),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_2495),
.Y(n_2966)
);

INVx6_ASAP7_75t_L g2967 ( 
.A(n_2491),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2536),
.B(n_1724),
.Y(n_2968)
);

BUFx6f_ASAP7_75t_L g2969 ( 
.A(n_2324),
.Y(n_2969)
);

INVxp67_ASAP7_75t_L g2970 ( 
.A(n_2416),
.Y(n_2970)
);

BUFx6f_ASAP7_75t_L g2971 ( 
.A(n_2324),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2306),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2231),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2425),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2425),
.Y(n_2975)
);

CKINVDCx5p33_ASAP7_75t_R g2976 ( 
.A(n_2495),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2425),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2543),
.B(n_1725),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2239),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2239),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2244),
.Y(n_2981)
);

CKINVDCx5p33_ASAP7_75t_R g2982 ( 
.A(n_2260),
.Y(n_2982)
);

CKINVDCx5p33_ASAP7_75t_R g2983 ( 
.A(n_2260),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_2380),
.Y(n_2984)
);

HB1xp67_ASAP7_75t_L g2985 ( 
.A(n_2543),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2244),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2260),
.Y(n_2987)
);

CKINVDCx5p33_ASAP7_75t_R g2988 ( 
.A(n_2288),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_2288),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2306),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2306),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2308),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2259),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2308),
.Y(n_2994)
);

NAND2xp33_ASAP7_75t_SL g2995 ( 
.A(n_2243),
.B(n_743),
.Y(n_2995)
);

INVx4_ASAP7_75t_L g2996 ( 
.A(n_2467),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2257),
.B(n_1725),
.Y(n_2997)
);

AOI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2272),
.A2(n_2583),
.B1(n_2543),
.B2(n_2580),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2288),
.Y(n_2999)
);

AND2x4_ASAP7_75t_L g3000 ( 
.A(n_2340),
.B(n_1161),
.Y(n_3000)
);

INVxp67_ASAP7_75t_L g3001 ( 
.A(n_2428),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2330),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2330),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2308),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2316),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2259),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2316),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2316),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2263),
.Y(n_3009)
);

BUFx6f_ASAP7_75t_L g3010 ( 
.A(n_2467),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2336),
.B(n_1729),
.Y(n_3011)
);

CKINVDCx5p33_ASAP7_75t_R g3012 ( 
.A(n_2347),
.Y(n_3012)
);

INVxp67_ASAP7_75t_L g3013 ( 
.A(n_2444),
.Y(n_3013)
);

AND3x2_ASAP7_75t_L g3014 ( 
.A(n_2574),
.B(n_1239),
.C(n_1092),
.Y(n_3014)
);

INVx3_ASAP7_75t_L g3015 ( 
.A(n_2235),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2581),
.B(n_2533),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2321),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2321),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_2347),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2263),
.Y(n_3020)
);

CKINVDCx20_ASAP7_75t_R g3021 ( 
.A(n_2607),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2321),
.Y(n_3022)
);

NOR2xp67_ASAP7_75t_L g3023 ( 
.A(n_2491),
.B(n_1729),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_2347),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2336),
.B(n_1734),
.Y(n_3025)
);

HB1xp67_ASAP7_75t_L g3026 ( 
.A(n_2580),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2340),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2581),
.B(n_1734),
.Y(n_3028)
);

CKINVDCx5p33_ASAP7_75t_R g3029 ( 
.A(n_2381),
.Y(n_3029)
);

BUFx6f_ASAP7_75t_L g3030 ( 
.A(n_2467),
.Y(n_3030)
);

CKINVDCx20_ASAP7_75t_R g3031 ( 
.A(n_2607),
.Y(n_3031)
);

HB1xp67_ASAP7_75t_L g3032 ( 
.A(n_2598),
.Y(n_3032)
);

BUFx2_ASAP7_75t_L g3033 ( 
.A(n_2380),
.Y(n_3033)
);

CKINVDCx5p33_ASAP7_75t_R g3034 ( 
.A(n_2381),
.Y(n_3034)
);

CKINVDCx5p33_ASAP7_75t_R g3035 ( 
.A(n_2554),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2477),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2340),
.Y(n_3037)
);

CKINVDCx5p33_ASAP7_75t_R g3038 ( 
.A(n_2554),
.Y(n_3038)
);

HB1xp67_ASAP7_75t_L g3039 ( 
.A(n_2598),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2376),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2376),
.Y(n_3041)
);

HB1xp67_ASAP7_75t_L g3042 ( 
.A(n_2598),
.Y(n_3042)
);

CKINVDCx5p33_ASAP7_75t_R g3043 ( 
.A(n_2554),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2265),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2265),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2423),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2376),
.Y(n_3047)
);

BUFx2_ASAP7_75t_SL g3048 ( 
.A(n_2495),
.Y(n_3048)
);

HB1xp67_ASAP7_75t_L g3049 ( 
.A(n_2489),
.Y(n_3049)
);

HB1xp67_ASAP7_75t_L g3050 ( 
.A(n_2489),
.Y(n_3050)
);

BUFx6f_ASAP7_75t_L g3051 ( 
.A(n_2477),
.Y(n_3051)
);

CKINVDCx5p33_ASAP7_75t_R g3052 ( 
.A(n_2554),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2423),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_2554),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2477),
.Y(n_3055)
);

BUFx2_ASAP7_75t_L g3056 ( 
.A(n_2380),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2397),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2281),
.B(n_1735),
.Y(n_3058)
);

AND2x2_ASAP7_75t_SL g3059 ( 
.A(n_2583),
.B(n_1173),
.Y(n_3059)
);

BUFx10_ASAP7_75t_L g3060 ( 
.A(n_2497),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_2557),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_2557),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2367),
.Y(n_3063)
);

CKINVDCx20_ASAP7_75t_R g3064 ( 
.A(n_2611),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2336),
.B(n_2445),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2397),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2557),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_2557),
.Y(n_3068)
);

BUFx2_ASAP7_75t_L g3069 ( 
.A(n_2599),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2367),
.Y(n_3070)
);

CKINVDCx5p33_ASAP7_75t_R g3071 ( 
.A(n_2557),
.Y(n_3071)
);

AND2x4_ASAP7_75t_L g3072 ( 
.A(n_2397),
.B(n_1173),
.Y(n_3072)
);

INVx3_ASAP7_75t_L g3073 ( 
.A(n_2241),
.Y(n_3073)
);

CKINVDCx5p33_ASAP7_75t_R g3074 ( 
.A(n_2565),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2418),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_2565),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2367),
.Y(n_3077)
);

CKINVDCx5p33_ASAP7_75t_R g3078 ( 
.A(n_2565),
.Y(n_3078)
);

CKINVDCx5p33_ASAP7_75t_R g3079 ( 
.A(n_2565),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2418),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2418),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2442),
.Y(n_3082)
);

CKINVDCx5p33_ASAP7_75t_R g3083 ( 
.A(n_2565),
.Y(n_3083)
);

CKINVDCx5p33_ASAP7_75t_R g3084 ( 
.A(n_2588),
.Y(n_3084)
);

OA21x2_ASAP7_75t_L g3085 ( 
.A1(n_2499),
.A2(n_1737),
.B(n_1735),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2442),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2588),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2442),
.Y(n_3088)
);

CKINVDCx5p33_ASAP7_75t_R g3089 ( 
.A(n_2588),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2693),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_SL g3091 ( 
.A(n_3035),
.B(n_2588),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2693),
.Y(n_3092)
);

INVx1_ASAP7_75t_SL g3093 ( 
.A(n_2795),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2656),
.B(n_2755),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2702),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2702),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2619),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2706),
.Y(n_3098)
);

OR2x6_ASAP7_75t_L g3099 ( 
.A(n_3048),
.B(n_2495),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_3010),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2706),
.Y(n_3101)
);

INVxp33_ASAP7_75t_L g3102 ( 
.A(n_2617),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2625),
.B(n_2170),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2709),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_2614),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2709),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2738),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_3035),
.B(n_2588),
.Y(n_3108)
);

INVx3_ASAP7_75t_L g3109 ( 
.A(n_3010),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2738),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_3038),
.B(n_3043),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2746),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_3010),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2746),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2654),
.B(n_2179),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2619),
.Y(n_3116)
);

INVxp33_ASAP7_75t_L g3117 ( 
.A(n_2840),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_SL g3118 ( 
.A(n_3038),
.B(n_2501),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2831),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2750),
.Y(n_3120)
);

HB1xp67_ASAP7_75t_L g3121 ( 
.A(n_2634),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2622),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2750),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_3043),
.B(n_3052),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2793),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2793),
.Y(n_3126)
);

CKINVDCx5p33_ASAP7_75t_R g3127 ( 
.A(n_2620),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_3052),
.B(n_2501),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2622),
.Y(n_3129)
);

OR2x6_ASAP7_75t_L g3130 ( 
.A(n_2743),
.B(n_2501),
.Y(n_3130)
);

CKINVDCx5p33_ASAP7_75t_R g3131 ( 
.A(n_2624),
.Y(n_3131)
);

AO22x2_ASAP7_75t_L g3132 ( 
.A1(n_3059),
.A2(n_2551),
.B1(n_2555),
.B2(n_2552),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_SL g3133 ( 
.A(n_3054),
.B(n_2501),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_2902),
.B(n_2532),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2797),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_3010),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2797),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2802),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2802),
.Y(n_3139)
);

BUFx3_ASAP7_75t_L g3140 ( 
.A(n_2886),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_3054),
.B(n_3061),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2811),
.Y(n_3142)
);

BUFx3_ASAP7_75t_L g3143 ( 
.A(n_2886),
.Y(n_3143)
);

INVx2_ASAP7_75t_SL g3144 ( 
.A(n_2641),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2659),
.B(n_2294),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2811),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2830),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2830),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2833),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2833),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2655),
.B(n_2461),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2844),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2844),
.Y(n_3153)
);

INVx5_ASAP7_75t_L g3154 ( 
.A(n_3030),
.Y(n_3154)
);

INVx2_ASAP7_75t_SL g3155 ( 
.A(n_2665),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2856),
.Y(n_3156)
);

BUFx3_ASAP7_75t_L g3157 ( 
.A(n_2967),
.Y(n_3157)
);

INVx4_ASAP7_75t_L g3158 ( 
.A(n_2770),
.Y(n_3158)
);

OR2x2_ASAP7_75t_L g3159 ( 
.A(n_2668),
.B(n_2595),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2856),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2860),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_3030),
.Y(n_3162)
);

BUFx3_ASAP7_75t_L g3163 ( 
.A(n_2967),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2860),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_3061),
.B(n_2501),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2870),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2870),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_SL g3168 ( 
.A(n_3062),
.B(n_2511),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2871),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2871),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2872),
.Y(n_3171)
);

INVx3_ASAP7_75t_L g3172 ( 
.A(n_3030),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2635),
.Y(n_3173)
);

CKINVDCx5p33_ASAP7_75t_R g3174 ( 
.A(n_2626),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2872),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2879),
.Y(n_3176)
);

BUFx6f_ASAP7_75t_L g3177 ( 
.A(n_3030),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2635),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2638),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_SL g3180 ( 
.A(n_3062),
.B(n_2511),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2638),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2879),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2644),
.Y(n_3183)
);

BUFx4f_ASAP7_75t_L g3184 ( 
.A(n_2967),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2644),
.Y(n_3185)
);

NOR2xp33_ASAP7_75t_L g3186 ( 
.A(n_2673),
.B(n_2560),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2898),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2898),
.Y(n_3188)
);

INVx1_ASAP7_75t_SL g3189 ( 
.A(n_2701),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2900),
.Y(n_3190)
);

AND2x4_ASAP7_75t_L g3191 ( 
.A(n_2859),
.B(n_2582),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2900),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2901),
.Y(n_3193)
);

INVx8_ASAP7_75t_L g3194 ( 
.A(n_2824),
.Y(n_3194)
);

INVx1_ASAP7_75t_SL g3195 ( 
.A(n_2788),
.Y(n_3195)
);

AND3x2_ASAP7_75t_L g3196 ( 
.A(n_3069),
.B(n_2577),
.C(n_2528),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2901),
.Y(n_3197)
);

INVx2_ASAP7_75t_SL g3198 ( 
.A(n_2768),
.Y(n_3198)
);

INVx3_ASAP7_75t_L g3199 ( 
.A(n_3036),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_SL g3200 ( 
.A(n_3067),
.B(n_2511),
.Y(n_3200)
);

NAND3xp33_ASAP7_75t_L g3201 ( 
.A(n_2995),
.B(n_2527),
.C(n_2524),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2912),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2912),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2926),
.Y(n_3204)
);

NOR2xp33_ASAP7_75t_L g3205 ( 
.A(n_2676),
.B(n_2576),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2732),
.B(n_2304),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_3067),
.B(n_2511),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2926),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2932),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_SL g3210 ( 
.A(n_3068),
.B(n_2511),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2932),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_2631),
.B(n_2559),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_3068),
.B(n_2545),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_2947),
.Y(n_3214)
);

AND3x2_ASAP7_75t_L g3215 ( 
.A(n_3016),
.B(n_2567),
.C(n_2517),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_SL g3216 ( 
.A(n_3071),
.B(n_2545),
.Y(n_3216)
);

INVx5_ASAP7_75t_L g3217 ( 
.A(n_3036),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2629),
.B(n_2322),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2947),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2973),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2973),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_3071),
.B(n_2545),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2810),
.B(n_2486),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2645),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2645),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2681),
.Y(n_3226)
);

CKINVDCx6p67_ASAP7_75t_R g3227 ( 
.A(n_2630),
.Y(n_3227)
);

AND2x2_ASAP7_75t_SL g3228 ( 
.A(n_3059),
.B(n_2524),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2681),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_3036),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_3074),
.B(n_2545),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2974),
.Y(n_3232)
);

BUFx3_ASAP7_75t_L g3233 ( 
.A(n_2821),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2692),
.Y(n_3234)
);

INVxp33_ASAP7_75t_L g3235 ( 
.A(n_2847),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_3036),
.Y(n_3236)
);

AOI21x1_ASAP7_75t_L g3237 ( 
.A1(n_2839),
.A2(n_2289),
.B(n_2270),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2692),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2974),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2975),
.Y(n_3240)
);

CKINVDCx20_ASAP7_75t_R g3241 ( 
.A(n_2736),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2674),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2975),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_3074),
.B(n_3076),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2674),
.Y(n_3245)
);

INVx8_ASAP7_75t_L g3246 ( 
.A(n_2824),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2977),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2675),
.Y(n_3248)
);

INVxp33_ASAP7_75t_SL g3249 ( 
.A(n_2895),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_3076),
.B(n_2545),
.Y(n_3250)
);

INVx2_ASAP7_75t_SL g3251 ( 
.A(n_2642),
.Y(n_3251)
);

BUFx10_ASAP7_75t_L g3252 ( 
.A(n_2791),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2977),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2675),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_3078),
.B(n_2550),
.Y(n_3255)
);

INVx4_ASAP7_75t_L g3256 ( 
.A(n_2770),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2979),
.Y(n_3257)
);

BUFx6f_ASAP7_75t_SL g3258 ( 
.A(n_3060),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2646),
.Y(n_3259)
);

INVx2_ASAP7_75t_SL g3260 ( 
.A(n_2642),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2979),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_2940),
.B(n_2492),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2646),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_SL g3264 ( 
.A(n_3078),
.B(n_2550),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2652),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2652),
.Y(n_3266)
);

INVx1_ASAP7_75t_SL g3267 ( 
.A(n_2832),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_2657),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2980),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_L g3270 ( 
.A(n_2754),
.B(n_2498),
.Y(n_3270)
);

BUFx4f_ASAP7_75t_L g3271 ( 
.A(n_2772),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2657),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2980),
.Y(n_3273)
);

INVx4_ASAP7_75t_L g3274 ( 
.A(n_2770),
.Y(n_3274)
);

OR2x2_ASAP7_75t_L g3275 ( 
.A(n_2703),
.B(n_2596),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2981),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2667),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2667),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3055),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2981),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_3051),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2986),
.Y(n_3282)
);

AND3x2_ASAP7_75t_L g3283 ( 
.A(n_3032),
.B(n_2589),
.C(n_2573),
.Y(n_3283)
);

INVx4_ASAP7_75t_L g3284 ( 
.A(n_2776),
.Y(n_3284)
);

HB1xp67_ASAP7_75t_L g3285 ( 
.A(n_3039),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2986),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3055),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_SL g3288 ( 
.A(n_3079),
.B(n_2550),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_3079),
.B(n_2550),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3063),
.Y(n_3290)
);

CKINVDCx5p33_ASAP7_75t_R g3291 ( 
.A(n_2905),
.Y(n_3291)
);

INVx2_ASAP7_75t_SL g3292 ( 
.A(n_2642),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2993),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2997),
.B(n_2365),
.Y(n_3294)
);

NAND2xp33_ASAP7_75t_L g3295 ( 
.A(n_3083),
.B(n_3084),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_3063),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3070),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2993),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3070),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3006),
.Y(n_3300)
);

CKINVDCx16_ASAP7_75t_R g3301 ( 
.A(n_2957),
.Y(n_3301)
);

AND2x4_ASAP7_75t_L g3302 ( 
.A(n_2862),
.B(n_2582),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3006),
.Y(n_3303)
);

BUFx6f_ASAP7_75t_L g3304 ( 
.A(n_3051),
.Y(n_3304)
);

BUFx6f_ASAP7_75t_L g3305 ( 
.A(n_3051),
.Y(n_3305)
);

AND2x6_ASAP7_75t_L g3306 ( 
.A(n_3077),
.B(n_2550),
.Y(n_3306)
);

NOR2xp33_ASAP7_75t_L g3307 ( 
.A(n_3058),
.B(n_2509),
.Y(n_3307)
);

INVx2_ASAP7_75t_SL g3308 ( 
.A(n_2814),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3077),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3009),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3009),
.Y(n_3311)
);

INVx8_ASAP7_75t_L g3312 ( 
.A(n_2824),
.Y(n_3312)
);

INVxp67_ASAP7_75t_SL g3313 ( 
.A(n_2776),
.Y(n_3313)
);

AOI22xp5_ASAP7_75t_L g3314 ( 
.A1(n_2995),
.A2(n_2524),
.B1(n_2527),
.B2(n_2559),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3020),
.Y(n_3315)
);

CKINVDCx6p67_ASAP7_75t_R g3316 ( 
.A(n_2640),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2776),
.B(n_2379),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3020),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_3083),
.B(n_2551),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3044),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_3051),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3044),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2841),
.B(n_2458),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3045),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3045),
.Y(n_3325)
);

INVxp33_ASAP7_75t_SL g3326 ( 
.A(n_2909),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3046),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3046),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2841),
.B(n_2478),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3053),
.Y(n_3330)
);

AND3x2_ASAP7_75t_L g3331 ( 
.A(n_3042),
.B(n_1239),
.C(n_1092),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_SL g3332 ( 
.A(n_2916),
.B(n_2443),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3053),
.Y(n_3333)
);

BUFx2_ASAP7_75t_L g3334 ( 
.A(n_3084),
.Y(n_3334)
);

INVx2_ASAP7_75t_SL g3335 ( 
.A(n_2814),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2841),
.B(n_2445),
.Y(n_3336)
);

INVx2_ASAP7_75t_SL g3337 ( 
.A(n_2814),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_2851),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_2623),
.Y(n_3339)
);

INVx2_ASAP7_75t_SL g3340 ( 
.A(n_2823),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_2636),
.B(n_2572),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_3087),
.B(n_2585),
.Y(n_3342)
);

INVx4_ASAP7_75t_L g3343 ( 
.A(n_2851),
.Y(n_3343)
);

NOR2x1p5_ASAP7_75t_L g3344 ( 
.A(n_2868),
.B(n_2490),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2857),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2711),
.Y(n_3346)
);

OR2x6_ASAP7_75t_L g3347 ( 
.A(n_2756),
.B(n_2493),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3087),
.B(n_2585),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_L g3349 ( 
.A(n_2914),
.B(n_2552),
.Y(n_3349)
);

INVxp67_ASAP7_75t_L g3350 ( 
.A(n_2861),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_2623),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_2845),
.B(n_2555),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2713),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2623),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2639),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_2639),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2715),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_2639),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2851),
.B(n_2445),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2996),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_2996),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_2996),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_3089),
.B(n_2570),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_3089),
.B(n_2570),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_2998),
.A2(n_2507),
.B1(n_2514),
.B2(n_2493),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_2897),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_2897),
.Y(n_3367)
);

OR2x2_ASAP7_75t_L g3368 ( 
.A(n_2689),
.B(n_2605),
.Y(n_3368)
);

BUFx3_ASAP7_75t_L g3369 ( 
.A(n_2821),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_2897),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2612),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_2911),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2911),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2616),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2621),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_2911),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2662),
.Y(n_3377)
);

NAND2xp33_ASAP7_75t_SL g3378 ( 
.A(n_2918),
.B(n_2592),
.Y(n_3378)
);

AND3x2_ASAP7_75t_L g3379 ( 
.A(n_2744),
.B(n_1267),
.C(n_2283),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2664),
.Y(n_3380)
);

BUFx8_ASAP7_75t_SL g3381 ( 
.A(n_2787),
.Y(n_3381)
);

AO21x2_ASAP7_75t_L g3382 ( 
.A1(n_2686),
.A2(n_2553),
.B(n_2173),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_2666),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2669),
.Y(n_3384)
);

INVxp33_ASAP7_75t_SL g3385 ( 
.A(n_2919),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2671),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2820),
.B(n_2445),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2677),
.Y(n_3388)
);

INVx3_ASAP7_75t_L g3389 ( 
.A(n_2913),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_2678),
.Y(n_3390)
);

NAND2xp33_ASAP7_75t_R g3391 ( 
.A(n_2663),
.B(n_2572),
.Y(n_3391)
);

OAI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_2922),
.A2(n_2533),
.B1(n_2578),
.B2(n_2568),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_2827),
.B(n_2445),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_2682),
.Y(n_3394)
);

INVx2_ASAP7_75t_SL g3395 ( 
.A(n_2823),
.Y(n_3395)
);

NAND2xp33_ASAP7_75t_L g3396 ( 
.A(n_2960),
.B(n_2592),
.Y(n_3396)
);

BUFx10_ASAP7_75t_L g3397 ( 
.A(n_3029),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2683),
.Y(n_3398)
);

INVx3_ASAP7_75t_L g3399 ( 
.A(n_2913),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_SL g3400 ( 
.A(n_2961),
.B(n_2590),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_2684),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_2687),
.Y(n_3402)
);

OAI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_2966),
.A2(n_2578),
.B1(n_2568),
.B2(n_2490),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2695),
.Y(n_3404)
);

NAND3xp33_ASAP7_75t_L g3405 ( 
.A(n_2828),
.B(n_2527),
.C(n_2572),
.Y(n_3405)
);

BUFx6f_ASAP7_75t_L g3406 ( 
.A(n_2618),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2696),
.Y(n_3407)
);

INVx3_ASAP7_75t_L g3408 ( 
.A(n_2913),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2698),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_2699),
.Y(n_3410)
);

INVx2_ASAP7_75t_SL g3411 ( 
.A(n_2823),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2700),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_2976),
.B(n_2590),
.Y(n_3413)
);

BUFx3_ASAP7_75t_L g3414 ( 
.A(n_2821),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2704),
.Y(n_3415)
);

NAND2xp33_ASAP7_75t_L g3416 ( 
.A(n_2772),
.B(n_2824),
.Y(n_3416)
);

INVxp67_ASAP7_75t_SL g3417 ( 
.A(n_2618),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_2962),
.B(n_2590),
.Y(n_3418)
);

INVx3_ASAP7_75t_L g3419 ( 
.A(n_2925),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_2710),
.Y(n_3420)
);

INVxp33_ASAP7_75t_SL g3421 ( 
.A(n_2725),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2942),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_2943),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2944),
.Y(n_3424)
);

AND3x1_ASAP7_75t_L g3425 ( 
.A(n_2880),
.B(n_2549),
.C(n_2503),
.Y(n_3425)
);

INVx2_ASAP7_75t_SL g3426 ( 
.A(n_3026),
.Y(n_3426)
);

CKINVDCx6p67_ASAP7_75t_R g3427 ( 
.A(n_2640),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_2834),
.B(n_2448),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_2946),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_2948),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_SL g3431 ( 
.A(n_2962),
.B(n_2590),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_2962),
.B(n_2590),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_2618),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_2949),
.Y(n_3434)
);

AO21x2_ASAP7_75t_L g3435 ( 
.A1(n_2686),
.A2(n_2553),
.B(n_2173),
.Y(n_3435)
);

INVx2_ASAP7_75t_SL g3436 ( 
.A(n_3049),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2950),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2955),
.Y(n_3438)
);

BUFx3_ASAP7_75t_L g3439 ( 
.A(n_2821),
.Y(n_3439)
);

CKINVDCx6p67_ASAP7_75t_R g3440 ( 
.A(n_2660),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_2850),
.B(n_2575),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_2962),
.B(n_2490),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2956),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2854),
.B(n_2894),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_2958),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_2963),
.Y(n_3446)
);

AO21x2_ASAP7_75t_L g3447 ( 
.A1(n_3065),
.A2(n_2351),
.B(n_2289),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_2964),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_2972),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_2965),
.B(n_2540),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_2990),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2991),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_2992),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_2896),
.B(n_2448),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_2994),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_SL g3456 ( 
.A(n_2965),
.B(n_2969),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3004),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_2970),
.B(n_2568),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_2637),
.Y(n_3459)
);

CKINVDCx6p67_ASAP7_75t_R g3460 ( 
.A(n_2660),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_2647),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2904),
.B(n_2448),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2658),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_2925),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_2772),
.B(n_2448),
.Y(n_3465)
);

INVx3_ASAP7_75t_L g3466 ( 
.A(n_2925),
.Y(n_3466)
);

BUFx6f_ASAP7_75t_L g3467 ( 
.A(n_2618),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_2931),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2931),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2931),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_2772),
.B(n_2448),
.Y(n_3471)
);

CKINVDCx20_ASAP7_75t_R g3472 ( 
.A(n_2736),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_2938),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_2938),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_2938),
.Y(n_3475)
);

INVx2_ASAP7_75t_SL g3476 ( 
.A(n_3050),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3015),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3015),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3015),
.Y(n_3479)
);

BUFx2_ASAP7_75t_L g3480 ( 
.A(n_2951),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3001),
.B(n_2578),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3073),
.Y(n_3482)
);

NAND3xp33_ASAP7_75t_L g3483 ( 
.A(n_2954),
.B(n_2575),
.C(n_2480),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3073),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3073),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_2863),
.Y(n_3486)
);

INVx3_ASAP7_75t_L g3487 ( 
.A(n_2869),
.Y(n_3487)
);

INVx3_ASAP7_75t_L g3488 ( 
.A(n_2869),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_2697),
.B(n_2600),
.Y(n_3489)
);

INVx5_ASAP7_75t_L g3490 ( 
.A(n_2824),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_2874),
.Y(n_3491)
);

OAI22xp5_ASAP7_75t_L g3492 ( 
.A1(n_2881),
.A2(n_2514),
.B1(n_2518),
.B2(n_2507),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_2965),
.B(n_2540),
.Y(n_3493)
);

BUFx6f_ASAP7_75t_L g3494 ( 
.A(n_2628),
.Y(n_3494)
);

BUFx2_ASAP7_75t_L g3495 ( 
.A(n_2951),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_2874),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_2748),
.B(n_2575),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_2921),
.Y(n_3498)
);

XOR2xp5_ASAP7_75t_L g3499 ( 
.A(n_2712),
.B(n_1861),
.Y(n_3499)
);

BUFx16f_ASAP7_75t_R g3500 ( 
.A(n_2688),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_2921),
.Y(n_3501)
);

INVx3_ASAP7_75t_L g3502 ( 
.A(n_2869),
.Y(n_3502)
);

NOR2x1p5_ASAP7_75t_L g3503 ( 
.A(n_2927),
.B(n_2540),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_2936),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_2936),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_2921),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_2716),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2936),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_2772),
.B(n_2449),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_2718),
.Y(n_3510)
);

BUFx2_ASAP7_75t_L g3511 ( 
.A(n_2959),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_2773),
.B(n_3000),
.Y(n_3512)
);

BUFx8_ASAP7_75t_SL g3513 ( 
.A(n_2787),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_2720),
.Y(n_3514)
);

NOR2x1p5_ASAP7_75t_L g3515 ( 
.A(n_2928),
.B(n_2443),
.Y(n_3515)
);

BUFx4f_ASAP7_75t_L g3516 ( 
.A(n_2772),
.Y(n_3516)
);

NOR3xp33_ASAP7_75t_L g3517 ( 
.A(n_2762),
.B(n_2597),
.C(n_2602),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_2722),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3000),
.B(n_2489),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_2936),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_2855),
.B(n_2449),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_2937),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_2937),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_2726),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_2727),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_SL g3526 ( 
.A(n_2965),
.B(n_2592),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_2729),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_2937),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_2937),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_2730),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2941),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_2731),
.Y(n_3532)
);

AND2x4_ASAP7_75t_L g3533 ( 
.A(n_3005),
.B(n_2518),
.Y(n_3533)
);

BUFx10_ASAP7_75t_L g3534 ( 
.A(n_3029),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_2739),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_2740),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3000),
.B(n_2512),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_2742),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_2751),
.Y(n_3539)
);

INVx3_ASAP7_75t_L g3540 ( 
.A(n_2869),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_2752),
.B(n_2449),
.Y(n_3541)
);

NAND3xp33_ASAP7_75t_L g3542 ( 
.A(n_2759),
.B(n_2764),
.C(n_2761),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_2766),
.B(n_2449),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_2769),
.B(n_2449),
.Y(n_3544)
);

INVx2_ASAP7_75t_SL g3545 ( 
.A(n_2765),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_2774),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_2941),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_2775),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_2941),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_2777),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_2780),
.B(n_2786),
.Y(n_3551)
);

OR2x6_ASAP7_75t_L g3552 ( 
.A(n_2945),
.B(n_2522),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_2941),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_2969),
.B(n_2592),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_2969),
.B(n_2592),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_2952),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_2790),
.B(n_2452),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_2969),
.B(n_2594),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_SL g3559 ( 
.A(n_2971),
.B(n_2594),
.Y(n_3559)
);

INVx2_ASAP7_75t_SL g3560 ( 
.A(n_2803),
.Y(n_3560)
);

NAND2xp33_ASAP7_75t_L g3561 ( 
.A(n_2824),
.B(n_2594),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_2796),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_L g3563 ( 
.A(n_3013),
.B(n_2813),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_2952),
.Y(n_3564)
);

INVx3_ASAP7_75t_L g3565 ( 
.A(n_2887),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_2798),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_2799),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_2800),
.Y(n_3568)
);

INVx2_ASAP7_75t_SL g3569 ( 
.A(n_2806),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3072),
.B(n_2512),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_2952),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_2801),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_2952),
.Y(n_3573)
);

BUFx4f_ASAP7_75t_L g3574 ( 
.A(n_2849),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_2971),
.B(n_2594),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_2724),
.Y(n_3576)
);

OAI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_2984),
.A2(n_2523),
.B1(n_2526),
.B2(n_2522),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_2971),
.B(n_2594),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_2971),
.B(n_2443),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_2805),
.Y(n_3580)
);

INVx2_ASAP7_75t_SL g3581 ( 
.A(n_2808),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_2817),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_2818),
.B(n_2452),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_2846),
.B(n_2593),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_2724),
.Y(n_3585)
);

CKINVDCx5p33_ASAP7_75t_R g3586 ( 
.A(n_2734),
.Y(n_3586)
);

BUFx8_ASAP7_75t_SL g3587 ( 
.A(n_2809),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_2724),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_2819),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3007),
.Y(n_3590)
);

INVx2_ASAP7_75t_SL g3591 ( 
.A(n_2843),
.Y(n_3591)
);

INVxp33_ASAP7_75t_L g3592 ( 
.A(n_2883),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3072),
.B(n_2452),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3008),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3002),
.B(n_3003),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2835),
.Y(n_3596)
);

INVx3_ASAP7_75t_L g3597 ( 
.A(n_2887),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3072),
.B(n_2452),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_2835),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3017),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_3002),
.B(n_2513),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_2835),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3002),
.B(n_2513),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_2929),
.B(n_2325),
.Y(n_3604)
);

INVx3_ASAP7_75t_L g3605 ( 
.A(n_2887),
.Y(n_3605)
);

NAND3xp33_ASAP7_75t_L g3606 ( 
.A(n_3018),
.B(n_2480),
.C(n_2292),
.Y(n_3606)
);

INVx5_ASAP7_75t_L g3607 ( 
.A(n_2849),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3022),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3424),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3424),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_3349),
.B(n_2523),
.Y(n_3611)
);

NOR2xp33_ASAP7_75t_L g3612 ( 
.A(n_3094),
.B(n_2728),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3434),
.Y(n_3613)
);

INVx3_ASAP7_75t_L g3614 ( 
.A(n_3157),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3434),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_3134),
.B(n_2513),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3437),
.Y(n_3617)
);

INVxp33_ASAP7_75t_L g3618 ( 
.A(n_3121),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3095),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3437),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3443),
.Y(n_3621)
);

INVx2_ASAP7_75t_SL g3622 ( 
.A(n_3144),
.Y(n_3622)
);

INVx3_ASAP7_75t_L g3623 ( 
.A(n_3157),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3443),
.Y(n_3624)
);

BUFx10_ASAP7_75t_L g3625 ( 
.A(n_3127),
.Y(n_3625)
);

AOI22xp5_ASAP7_75t_L g3626 ( 
.A1(n_3307),
.A2(n_3011),
.B1(n_3025),
.B2(n_2985),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3445),
.Y(n_3627)
);

BUFx3_ASAP7_75t_L g3628 ( 
.A(n_3131),
.Y(n_3628)
);

INVx1_ASAP7_75t_SL g3629 ( 
.A(n_3189),
.Y(n_3629)
);

AND2x4_ASAP7_75t_L g3630 ( 
.A(n_3198),
.B(n_3027),
.Y(n_3630)
);

AOI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3604),
.A2(n_3028),
.B1(n_2794),
.B2(n_2735),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3445),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3186),
.B(n_2849),
.Y(n_3633)
);

INVx2_ASAP7_75t_SL g3634 ( 
.A(n_3144),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3451),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_L g3636 ( 
.A(n_3275),
.B(n_3034),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3451),
.Y(n_3637)
);

INVx1_ASAP7_75t_SL g3638 ( 
.A(n_3195),
.Y(n_3638)
);

NAND2xp33_ASAP7_75t_L g3639 ( 
.A(n_3306),
.B(n_2849),
.Y(n_3639)
);

INVx8_ASAP7_75t_L g3640 ( 
.A(n_3099),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3452),
.Y(n_3641)
);

INVx1_ASAP7_75t_SL g3642 ( 
.A(n_3267),
.Y(n_3642)
);

INVx4_ASAP7_75t_L g3643 ( 
.A(n_3099),
.Y(n_3643)
);

OR2x6_ASAP7_75t_L g3644 ( 
.A(n_3130),
.B(n_2611),
.Y(n_3644)
);

BUFx2_ASAP7_75t_L g3645 ( 
.A(n_3334),
.Y(n_3645)
);

OR2x2_ASAP7_75t_L g3646 ( 
.A(n_3093),
.B(n_2600),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3452),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3453),
.Y(n_3648)
);

INVxp67_ASAP7_75t_SL g3649 ( 
.A(n_3136),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3453),
.Y(n_3650)
);

BUFx6f_ASAP7_75t_L g3651 ( 
.A(n_3140),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_3275),
.B(n_3034),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3346),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_L g3654 ( 
.A1(n_3228),
.A2(n_2849),
.B1(n_2468),
.B2(n_3033),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3346),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_SL g3656 ( 
.A(n_3158),
.B(n_3002),
.Y(n_3656)
);

AND2x4_ASAP7_75t_L g3657 ( 
.A(n_3198),
.B(n_3037),
.Y(n_3657)
);

BUFx2_ASAP7_75t_L g3658 ( 
.A(n_3334),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3353),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3205),
.B(n_2849),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_SL g3661 ( 
.A(n_3262),
.B(n_2526),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3158),
.B(n_3003),
.Y(n_3662)
);

INVx4_ASAP7_75t_L g3663 ( 
.A(n_3099),
.Y(n_3663)
);

AO22x2_ASAP7_75t_L g3664 ( 
.A1(n_3201),
.A2(n_2610),
.B1(n_2604),
.B2(n_2434),
.Y(n_3664)
);

AO22x2_ASAP7_75t_L g3665 ( 
.A1(n_3201),
.A2(n_2610),
.B1(n_2604),
.B2(n_2602),
.Y(n_3665)
);

INVx2_ASAP7_75t_SL g3666 ( 
.A(n_3155),
.Y(n_3666)
);

NAND2x1p5_ASAP7_75t_L g3667 ( 
.A(n_3154),
.B(n_3003),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_3151),
.B(n_3060),
.Y(n_3668)
);

BUFx3_ASAP7_75t_L g3669 ( 
.A(n_3174),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3353),
.Y(n_3670)
);

BUFx2_ASAP7_75t_L g3671 ( 
.A(n_3291),
.Y(n_3671)
);

AND3x4_ASAP7_75t_L g3672 ( 
.A(n_3517),
.B(n_2584),
.C(n_2542),
.Y(n_3672)
);

NAND3xp33_ASAP7_75t_L g3673 ( 
.A(n_3223),
.B(n_2331),
.C(n_2564),
.Y(n_3673)
);

BUFx6f_ASAP7_75t_L g3674 ( 
.A(n_3140),
.Y(n_3674)
);

INVx3_ASAP7_75t_L g3675 ( 
.A(n_3157),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3357),
.Y(n_3676)
);

BUFx3_ASAP7_75t_L g3677 ( 
.A(n_3586),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_3421),
.Y(n_3678)
);

INVx3_ASAP7_75t_L g3679 ( 
.A(n_3163),
.Y(n_3679)
);

BUFx6f_ASAP7_75t_L g3680 ( 
.A(n_3140),
.Y(n_3680)
);

BUFx2_ASAP7_75t_L g3681 ( 
.A(n_3155),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3357),
.Y(n_3682)
);

AND2x2_ASAP7_75t_L g3683 ( 
.A(n_3592),
.B(n_2888),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3103),
.B(n_3040),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3480),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3371),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3218),
.B(n_3060),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3095),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3102),
.B(n_2906),
.Y(n_3689)
);

INVx4_ASAP7_75t_L g3690 ( 
.A(n_3099),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3096),
.Y(n_3691)
);

BUFx4f_ASAP7_75t_L g3692 ( 
.A(n_3227),
.Y(n_3692)
);

BUFx3_ASAP7_75t_L g3693 ( 
.A(n_3227),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3371),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3096),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3374),
.Y(n_3696)
);

AND2x6_ASAP7_75t_L g3697 ( 
.A(n_3136),
.B(n_3041),
.Y(n_3697)
);

INVx4_ASAP7_75t_L g3698 ( 
.A(n_3099),
.Y(n_3698)
);

AND2x4_ASAP7_75t_L g3699 ( 
.A(n_3512),
.B(n_3047),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_3381),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3512),
.B(n_2953),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3098),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3374),
.Y(n_3703)
);

CKINVDCx20_ASAP7_75t_R g3704 ( 
.A(n_3513),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3375),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_SL g3706 ( 
.A(n_3206),
.B(n_2535),
.Y(n_3706)
);

NOR2xp33_ASAP7_75t_L g3707 ( 
.A(n_3159),
.B(n_2508),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3375),
.Y(n_3708)
);

NAND3x1_ASAP7_75t_L g3709 ( 
.A(n_3500),
.B(n_2603),
.C(n_2601),
.Y(n_3709)
);

BUFx3_ASAP7_75t_L g3710 ( 
.A(n_3480),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3461),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3098),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3107),
.Y(n_3713)
);

AND2x6_ASAP7_75t_L g3714 ( 
.A(n_3136),
.B(n_3057),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3115),
.B(n_3066),
.Y(n_3715)
);

BUFx3_ASAP7_75t_L g3716 ( 
.A(n_3495),
.Y(n_3716)
);

AND3x2_ASAP7_75t_L g3717 ( 
.A(n_3332),
.B(n_3056),
.C(n_2539),
.Y(n_3717)
);

OAI22xp33_ASAP7_75t_L g3718 ( 
.A1(n_3294),
.A2(n_2717),
.B1(n_3080),
.B2(n_3075),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3461),
.Y(n_3719)
);

OR2x2_ASAP7_75t_L g3720 ( 
.A(n_3159),
.B(n_2741),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3270),
.B(n_2584),
.Y(n_3721)
);

OR2x2_ASAP7_75t_SL g3722 ( 
.A(n_3301),
.B(n_2825),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_SL g3723 ( 
.A(n_3271),
.B(n_2749),
.Y(n_3723)
);

AND2x6_ASAP7_75t_L g3724 ( 
.A(n_3136),
.B(n_3081),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3107),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3495),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3461),
.Y(n_3727)
);

NAND2x1p5_ASAP7_75t_L g3728 ( 
.A(n_3154),
.B(n_3003),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3135),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3145),
.B(n_3082),
.Y(n_3730)
);

INVx4_ASAP7_75t_L g3731 ( 
.A(n_3154),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3444),
.B(n_3086),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3350),
.B(n_2535),
.Y(n_3733)
);

INVx1_ASAP7_75t_SL g3734 ( 
.A(n_3489),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3119),
.B(n_2539),
.Y(n_3735)
);

NAND3xp33_ASAP7_75t_L g3736 ( 
.A(n_3584),
.B(n_2587),
.C(n_2566),
.Y(n_3736)
);

NAND3x1_ASAP7_75t_L g3737 ( 
.A(n_3458),
.B(n_2456),
.C(n_2301),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3135),
.Y(n_3738)
);

INVx2_ASAP7_75t_SL g3739 ( 
.A(n_3489),
.Y(n_3739)
);

BUFx2_ASAP7_75t_L g3740 ( 
.A(n_3511),
.Y(n_3740)
);

AO21x2_ASAP7_75t_L g3741 ( 
.A1(n_3576),
.A2(n_2908),
.B(n_2648),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3463),
.Y(n_3742)
);

NOR2xp33_ASAP7_75t_L g3743 ( 
.A(n_3385),
.B(n_2537),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3137),
.Y(n_3744)
);

OAI221xp5_ASAP7_75t_L g3745 ( 
.A1(n_3425),
.A2(n_3088),
.B1(n_1697),
.B2(n_2269),
.C(n_2439),
.Y(n_3745)
);

AND2x6_ASAP7_75t_L g3746 ( 
.A(n_3136),
.B(n_2537),
.Y(n_3746)
);

AOI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3425),
.A2(n_2930),
.B1(n_2968),
.B2(n_2877),
.Y(n_3747)
);

INVx5_ASAP7_75t_L g3748 ( 
.A(n_3162),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3137),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3511),
.Y(n_3750)
);

INVx1_ASAP7_75t_SL g3751 ( 
.A(n_3368),
.Y(n_3751)
);

AND2x4_ASAP7_75t_L g3752 ( 
.A(n_3344),
.B(n_3119),
.Y(n_3752)
);

CKINVDCx6p67_ASAP7_75t_R g3753 ( 
.A(n_3316),
.Y(n_3753)
);

AND2x6_ASAP7_75t_L g3754 ( 
.A(n_3162),
.B(n_2542),
.Y(n_3754)
);

CKINVDCx5p33_ASAP7_75t_R g3755 ( 
.A(n_3587),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3139),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3463),
.Y(n_3757)
);

AND2x4_ASAP7_75t_L g3758 ( 
.A(n_3344),
.B(n_2866),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3139),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3463),
.Y(n_3760)
);

INVx4_ASAP7_75t_L g3761 ( 
.A(n_3154),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3142),
.Y(n_3762)
);

OR2x6_ASAP7_75t_L g3763 ( 
.A(n_3130),
.B(n_2611),
.Y(n_3763)
);

INVx4_ASAP7_75t_L g3764 ( 
.A(n_3154),
.Y(n_3764)
);

INVx5_ASAP7_75t_L g3765 ( 
.A(n_3162),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3497),
.B(n_2836),
.Y(n_3766)
);

INVx5_ASAP7_75t_L g3767 ( 
.A(n_3162),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3142),
.Y(n_3768)
);

BUFx4f_ASAP7_75t_L g3769 ( 
.A(n_3316),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_SL g3770 ( 
.A(n_3252),
.B(n_3403),
.Y(n_3770)
);

NOR2xp33_ASAP7_75t_L g3771 ( 
.A(n_3249),
.B(n_2571),
.Y(n_3771)
);

INVx3_ASAP7_75t_L g3772 ( 
.A(n_3163),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3232),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3158),
.A2(n_2717),
.B1(n_3021),
.B2(n_2959),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3497),
.B(n_2836),
.Y(n_3775)
);

AND2x4_ASAP7_75t_L g3776 ( 
.A(n_3519),
.B(n_2876),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3232),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3519),
.B(n_2512),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3146),
.Y(n_3779)
);

NOR2xp33_ASAP7_75t_L g3780 ( 
.A(n_3326),
.B(n_2753),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_3158),
.B(n_2836),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3146),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3149),
.Y(n_3783)
);

BUFx8_ASAP7_75t_SL g3784 ( 
.A(n_3241),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3256),
.B(n_2836),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3279),
.B(n_2882),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3239),
.Y(n_3787)
);

INVx1_ASAP7_75t_SL g3788 ( 
.A(n_3368),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3149),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3239),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3152),
.Y(n_3791)
);

AOI22xp33_ASAP7_75t_L g3792 ( 
.A1(n_3228),
.A2(n_2468),
.B1(n_2440),
.B2(n_2389),
.Y(n_3792)
);

BUFx6f_ASAP7_75t_L g3793 ( 
.A(n_3143),
.Y(n_3793)
);

INVx4_ASAP7_75t_L g3794 ( 
.A(n_3154),
.Y(n_3794)
);

BUFx6f_ASAP7_75t_L g3795 ( 
.A(n_3143),
.Y(n_3795)
);

INVx4_ASAP7_75t_SL g3796 ( 
.A(n_3306),
.Y(n_3796)
);

INVx2_ASAP7_75t_SL g3797 ( 
.A(n_3379),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3279),
.B(n_2884),
.Y(n_3798)
);

BUFx6f_ASAP7_75t_L g3799 ( 
.A(n_3143),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3240),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_SL g3801 ( 
.A(n_3252),
.B(n_2569),
.Y(n_3801)
);

OAI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3580),
.A2(n_2717),
.B1(n_2892),
.B2(n_2891),
.Y(n_3802)
);

INVx3_ASAP7_75t_L g3803 ( 
.A(n_3163),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3240),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_SL g3805 ( 
.A(n_3252),
.B(n_2569),
.Y(n_3805)
);

CKINVDCx5p33_ASAP7_75t_R g3806 ( 
.A(n_3105),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3152),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3243),
.Y(n_3808)
);

OR2x2_ASAP7_75t_L g3809 ( 
.A(n_3285),
.B(n_2757),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3243),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3247),
.Y(n_3811)
);

INVx1_ASAP7_75t_SL g3812 ( 
.A(n_3212),
.Y(n_3812)
);

INVx2_ASAP7_75t_SL g3813 ( 
.A(n_3331),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3156),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3352),
.B(n_2758),
.Y(n_3815)
);

AND2x6_ASAP7_75t_L g3816 ( 
.A(n_3162),
.B(n_2899),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3247),
.Y(n_3817)
);

BUFx6f_ASAP7_75t_L g3818 ( 
.A(n_3233),
.Y(n_3818)
);

INVx4_ASAP7_75t_L g3819 ( 
.A(n_3217),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3253),
.Y(n_3820)
);

INVx4_ASAP7_75t_SL g3821 ( 
.A(n_3306),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_SL g3822 ( 
.A(n_3271),
.B(n_2760),
.Y(n_3822)
);

INVxp67_ASAP7_75t_L g3823 ( 
.A(n_3537),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3279),
.B(n_2903),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3253),
.Y(n_3825)
);

INVx1_ASAP7_75t_SL g3826 ( 
.A(n_3212),
.Y(n_3826)
);

NAND2xp33_ASAP7_75t_L g3827 ( 
.A(n_3306),
.B(n_2767),
.Y(n_3827)
);

AND2x4_ASAP7_75t_L g3828 ( 
.A(n_3537),
.B(n_2915),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3156),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3161),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_L g3831 ( 
.A(n_3252),
.B(n_2771),
.Y(n_3831)
);

INVx3_ASAP7_75t_L g3832 ( 
.A(n_3406),
.Y(n_3832)
);

OR2x2_ASAP7_75t_L g3833 ( 
.A(n_3545),
.B(n_2663),
.Y(n_3833)
);

OR2x2_ASAP7_75t_SL g3834 ( 
.A(n_3301),
.B(n_2611),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3257),
.Y(n_3835)
);

INVx1_ASAP7_75t_SL g3836 ( 
.A(n_3341),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3161),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3287),
.B(n_2920),
.Y(n_3838)
);

AND2x4_ASAP7_75t_L g3839 ( 
.A(n_3570),
.B(n_2924),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3257),
.Y(n_3840)
);

INVx6_ASAP7_75t_L g3841 ( 
.A(n_3397),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3570),
.B(n_2218),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3167),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3533),
.B(n_2933),
.Y(n_3844)
);

BUFx3_ASAP7_75t_L g3845 ( 
.A(n_3472),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3261),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3287),
.B(n_2480),
.Y(n_3847)
);

AND2x6_ASAP7_75t_L g3848 ( 
.A(n_3177),
.B(n_2520),
.Y(n_3848)
);

OAI21xp33_ASAP7_75t_L g3849 ( 
.A1(n_3563),
.A2(n_1741),
.B(n_1737),
.Y(n_3849)
);

CKINVDCx20_ASAP7_75t_R g3850 ( 
.A(n_3427),
.Y(n_3850)
);

OR2x2_ASAP7_75t_L g3851 ( 
.A(n_3545),
.B(n_2670),
.Y(n_3851)
);

CKINVDCx5p33_ASAP7_75t_R g3852 ( 
.A(n_3427),
.Y(n_3852)
);

NAND2x1p5_ASAP7_75t_L g3853 ( 
.A(n_3217),
.B(n_2721),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3287),
.B(n_2452),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3167),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3190),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3261),
.Y(n_3857)
);

NOR2xp33_ASAP7_75t_L g3858 ( 
.A(n_3319),
.B(n_2530),
.Y(n_3858)
);

NAND2x1p5_ASAP7_75t_L g3859 ( 
.A(n_3217),
.B(n_2733),
.Y(n_3859)
);

INVx3_ASAP7_75t_L g3860 ( 
.A(n_3406),
.Y(n_3860)
);

CKINVDCx5p33_ASAP7_75t_R g3861 ( 
.A(n_3440),
.Y(n_3861)
);

AND2x6_ASAP7_75t_L g3862 ( 
.A(n_3177),
.B(n_3230),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3269),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_SL g3864 ( 
.A(n_3256),
.B(n_2569),
.Y(n_3864)
);

AND2x6_ASAP7_75t_L g3865 ( 
.A(n_3177),
.B(n_2531),
.Y(n_3865)
);

INVx4_ASAP7_75t_L g3866 ( 
.A(n_3217),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3269),
.Y(n_3867)
);

OR2x6_ASAP7_75t_L g3868 ( 
.A(n_3130),
.B(n_2556),
.Y(n_3868)
);

NOR2xp33_ASAP7_75t_L g3869 ( 
.A(n_3342),
.B(n_2541),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3273),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3560),
.B(n_2670),
.Y(n_3871)
);

AO22x2_ASAP7_75t_L g3872 ( 
.A1(n_3405),
.A2(n_2203),
.B1(n_2978),
.B2(n_2500),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3348),
.B(n_2544),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3481),
.B(n_2494),
.Y(n_3874)
);

INVx4_ASAP7_75t_L g3875 ( 
.A(n_3217),
.Y(n_3875)
);

BUFx6f_ASAP7_75t_L g3876 ( 
.A(n_3233),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3273),
.Y(n_3877)
);

CKINVDCx16_ASAP7_75t_R g3878 ( 
.A(n_3499),
.Y(n_3878)
);

NOR2xp33_ASAP7_75t_L g3879 ( 
.A(n_3363),
.B(n_2546),
.Y(n_3879)
);

INVx4_ASAP7_75t_L g3880 ( 
.A(n_3217),
.Y(n_3880)
);

CKINVDCx5p33_ASAP7_75t_R g3881 ( 
.A(n_3440),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_3256),
.B(n_3274),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3276),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3177),
.B(n_2454),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3276),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3280),
.Y(n_3886)
);

BUFx6f_ASAP7_75t_L g3887 ( 
.A(n_3233),
.Y(n_3887)
);

NAND3xp33_ASAP7_75t_L g3888 ( 
.A(n_3365),
.B(n_2181),
.C(n_2230),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3177),
.B(n_2454),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_3460),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3436),
.B(n_2506),
.Y(n_3891)
);

CKINVDCx5p33_ASAP7_75t_R g3892 ( 
.A(n_3460),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3190),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3193),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_SL g3895 ( 
.A(n_3256),
.B(n_2569),
.Y(n_3895)
);

BUFx10_ASAP7_75t_L g3896 ( 
.A(n_3258),
.Y(n_3896)
);

BUFx10_ASAP7_75t_L g3897 ( 
.A(n_3258),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3280),
.Y(n_3898)
);

OAI22xp5_ASAP7_75t_SL g3899 ( 
.A1(n_3499),
.A2(n_2939),
.B1(n_2934),
.B2(n_1865),
.Y(n_3899)
);

AND2x2_ASAP7_75t_L g3900 ( 
.A(n_3436),
.B(n_3476),
.Y(n_3900)
);

BUFx4_ASAP7_75t_L g3901 ( 
.A(n_3258),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3406),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3282),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3282),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3193),
.Y(n_3905)
);

BUFx3_ASAP7_75t_L g3906 ( 
.A(n_3397),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3228),
.A2(n_2547),
.B1(n_2203),
.B2(n_2426),
.Y(n_3907)
);

HB1xp67_ASAP7_75t_L g3908 ( 
.A(n_3230),
.Y(n_3908)
);

NOR2xp33_ASAP7_75t_SL g3909 ( 
.A(n_3271),
.B(n_3516),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_SL g3910 ( 
.A(n_3274),
.B(n_2569),
.Y(n_3910)
);

BUFx2_ASAP7_75t_L g3911 ( 
.A(n_3130),
.Y(n_3911)
);

INVx2_ASAP7_75t_SL g3912 ( 
.A(n_3215),
.Y(n_3912)
);

INVx1_ASAP7_75t_SL g3913 ( 
.A(n_3341),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_L g3914 ( 
.A1(n_3441),
.A2(n_2426),
.B1(n_954),
.B2(n_854),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3230),
.B(n_2454),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3286),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3286),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3293),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3293),
.Y(n_3919)
);

BUFx6f_ASAP7_75t_L g3920 ( 
.A(n_3369),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3298),
.Y(n_3921)
);

BUFx6f_ASAP7_75t_L g3922 ( 
.A(n_3369),
.Y(n_3922)
);

INVx4_ASAP7_75t_L g3923 ( 
.A(n_3369),
.Y(n_3923)
);

BUFx6f_ASAP7_75t_L g3924 ( 
.A(n_3414),
.Y(n_3924)
);

BUFx3_ASAP7_75t_L g3925 ( 
.A(n_3397),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_3364),
.B(n_2262),
.Y(n_3926)
);

BUFx6f_ASAP7_75t_L g3927 ( 
.A(n_3414),
.Y(n_3927)
);

INVx4_ASAP7_75t_L g3928 ( 
.A(n_3414),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3197),
.Y(n_3929)
);

INVx4_ASAP7_75t_SL g3930 ( 
.A(n_3306),
.Y(n_3930)
);

OAI22xp5_ASAP7_75t_L g3931 ( 
.A1(n_3274),
.A2(n_2717),
.B1(n_3031),
.B2(n_3021),
.Y(n_3931)
);

BUFx6f_ASAP7_75t_L g3932 ( 
.A(n_3439),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3298),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3533),
.B(n_2491),
.Y(n_3934)
);

INVx3_ASAP7_75t_L g3935 ( 
.A(n_3406),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_SL g3936 ( 
.A(n_3274),
.B(n_2649),
.Y(n_3936)
);

INVx5_ASAP7_75t_L g3937 ( 
.A(n_3230),
.Y(n_3937)
);

NOR2xp33_ASAP7_75t_L g3938 ( 
.A(n_3111),
.B(n_2351),
.Y(n_3938)
);

CKINVDCx5p33_ASAP7_75t_R g3939 ( 
.A(n_3397),
.Y(n_3939)
);

BUFx3_ASAP7_75t_L g3940 ( 
.A(n_3534),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3230),
.B(n_2454),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3476),
.B(n_2248),
.Y(n_3942)
);

INVx3_ASAP7_75t_L g3943 ( 
.A(n_3406),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3300),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3197),
.Y(n_3945)
);

BUFx6f_ASAP7_75t_L g3946 ( 
.A(n_3439),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3281),
.B(n_2454),
.Y(n_3947)
);

AND2x6_ASAP7_75t_L g3948 ( 
.A(n_3281),
.B(n_2887),
.Y(n_3948)
);

INVx3_ASAP7_75t_L g3949 ( 
.A(n_3433),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3281),
.B(n_2455),
.Y(n_3950)
);

BUFx3_ASAP7_75t_L g3951 ( 
.A(n_3534),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3300),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3281),
.B(n_2455),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3202),
.Y(n_3954)
);

INVx4_ASAP7_75t_L g3955 ( 
.A(n_3439),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3303),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3303),
.Y(n_3957)
);

NOR2xp33_ASAP7_75t_L g3958 ( 
.A(n_3124),
.B(n_2556),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_SL g3959 ( 
.A(n_3284),
.B(n_3023),
.Y(n_3959)
);

BUFx6f_ASAP7_75t_SL g3960 ( 
.A(n_3534),
.Y(n_3960)
);

INVx3_ASAP7_75t_L g3961 ( 
.A(n_3433),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3310),
.Y(n_3962)
);

NOR2xp33_ASAP7_75t_L g3963 ( 
.A(n_3141),
.B(n_2556),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3281),
.B(n_2455),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3202),
.Y(n_3965)
);

INVx1_ASAP7_75t_SL g3966 ( 
.A(n_3441),
.Y(n_3966)
);

INVx5_ASAP7_75t_L g3967 ( 
.A(n_3304),
.Y(n_3967)
);

BUFx3_ASAP7_75t_L g3968 ( 
.A(n_3534),
.Y(n_3968)
);

BUFx6f_ASAP7_75t_L g3969 ( 
.A(n_3433),
.Y(n_3969)
);

NAND3xp33_ASAP7_75t_L g3970 ( 
.A(n_3542),
.B(n_1742),
.C(n_1741),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3304),
.B(n_2455),
.Y(n_3971)
);

NOR2xp33_ASAP7_75t_L g3972 ( 
.A(n_3244),
.B(n_2599),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3310),
.Y(n_3973)
);

NOR2xp33_ASAP7_75t_L g3974 ( 
.A(n_3117),
.B(n_2599),
.Y(n_3974)
);

BUFx6f_ASAP7_75t_L g3975 ( 
.A(n_3433),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3304),
.B(n_3305),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3203),
.Y(n_3977)
);

INVx1_ASAP7_75t_SL g3978 ( 
.A(n_3426),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3304),
.B(n_3305),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3311),
.Y(n_3980)
);

BUFx6f_ASAP7_75t_L g3981 ( 
.A(n_3433),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3311),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3203),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3204),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3560),
.B(n_2599),
.Y(n_3985)
);

INVx3_ASAP7_75t_L g3986 ( 
.A(n_3467),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3235),
.B(n_2599),
.Y(n_3987)
);

INVx3_ASAP7_75t_L g3988 ( 
.A(n_3467),
.Y(n_3988)
);

BUFx3_ASAP7_75t_L g3989 ( 
.A(n_3569),
.Y(n_3989)
);

BUFx6f_ASAP7_75t_L g3990 ( 
.A(n_3467),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3284),
.B(n_2885),
.Y(n_3991)
);

INVx1_ASAP7_75t_SL g3992 ( 
.A(n_3426),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3315),
.Y(n_3993)
);

NAND2xp33_ASAP7_75t_SL g3994 ( 
.A(n_3515),
.B(n_3031),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3315),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_SL g3996 ( 
.A(n_3284),
.B(n_2628),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3204),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3304),
.B(n_2455),
.Y(n_3998)
);

INVx2_ASAP7_75t_SL g3999 ( 
.A(n_3196),
.Y(n_3999)
);

NOR2xp33_ASAP7_75t_SL g4000 ( 
.A(n_3516),
.B(n_2672),
.Y(n_4000)
);

CKINVDCx16_ASAP7_75t_R g4001 ( 
.A(n_3391),
.Y(n_4001)
);

INVx3_ASAP7_75t_L g4002 ( 
.A(n_3467),
.Y(n_4002)
);

AND2x6_ASAP7_75t_L g4003 ( 
.A(n_3305),
.B(n_2917),
.Y(n_4003)
);

BUFx6f_ASAP7_75t_L g4004 ( 
.A(n_3467),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3320),
.Y(n_4005)
);

AOI22xp33_ASAP7_75t_L g4006 ( 
.A1(n_3132),
.A2(n_2426),
.B1(n_954),
.B2(n_854),
.Y(n_4006)
);

BUFx6f_ASAP7_75t_L g4007 ( 
.A(n_3494),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_L g4008 ( 
.A(n_3305),
.B(n_2463),
.Y(n_4008)
);

HB1xp67_ASAP7_75t_L g4009 ( 
.A(n_3305),
.Y(n_4009)
);

INVx3_ASAP7_75t_L g4010 ( 
.A(n_3494),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3320),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3321),
.B(n_2463),
.Y(n_4012)
);

HB1xp67_ASAP7_75t_L g4013 ( 
.A(n_3321),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_L g4014 ( 
.A(n_3551),
.B(n_2789),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3494),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3569),
.B(n_3581),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3325),
.Y(n_4017)
);

INVx4_ASAP7_75t_L g4018 ( 
.A(n_3184),
.Y(n_4018)
);

BUFx3_ASAP7_75t_L g4019 ( 
.A(n_3581),
.Y(n_4019)
);

INVx1_ASAP7_75t_SL g4020 ( 
.A(n_3591),
.Y(n_4020)
);

CKINVDCx5p33_ASAP7_75t_R g4021 ( 
.A(n_3130),
.Y(n_4021)
);

HB1xp67_ASAP7_75t_L g4022 ( 
.A(n_3321),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3325),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3327),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3211),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3327),
.Y(n_4026)
);

CKINVDCx20_ASAP7_75t_R g4027 ( 
.A(n_3378),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3321),
.B(n_3097),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3328),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3542),
.B(n_2789),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3321),
.B(n_3097),
.Y(n_4031)
);

INVx3_ASAP7_75t_L g4032 ( 
.A(n_3494),
.Y(n_4032)
);

OAI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_3580),
.A2(n_3589),
.B1(n_3582),
.B2(n_3510),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3328),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3097),
.B(n_2463),
.Y(n_4035)
);

BUFx2_ASAP7_75t_L g4036 ( 
.A(n_3591),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3284),
.B(n_3343),
.Y(n_4037)
);

BUFx10_ASAP7_75t_L g4038 ( 
.A(n_3283),
.Y(n_4038)
);

BUFx4f_ASAP7_75t_L g4039 ( 
.A(n_3347),
.Y(n_4039)
);

BUFx2_ASAP7_75t_L g4040 ( 
.A(n_3191),
.Y(n_4040)
);

INVx2_ASAP7_75t_SL g4041 ( 
.A(n_3503),
.Y(n_4041)
);

INVx1_ASAP7_75t_SL g4042 ( 
.A(n_3533),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3116),
.B(n_2463),
.Y(n_4043)
);

OR2x2_ASAP7_75t_L g4044 ( 
.A(n_3507),
.B(n_2606),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3116),
.B(n_2463),
.Y(n_4045)
);

INVx5_ASAP7_75t_L g4046 ( 
.A(n_3306),
.Y(n_4046)
);

INVx4_ASAP7_75t_SL g4047 ( 
.A(n_3306),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3507),
.B(n_2606),
.Y(n_4048)
);

AND2x6_ASAP7_75t_L g4049 ( 
.A(n_3100),
.B(n_2917),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_3510),
.B(n_2792),
.Y(n_4050)
);

BUFx3_ASAP7_75t_L g4051 ( 
.A(n_3533),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3330),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_L g4053 ( 
.A1(n_3132),
.A2(n_2426),
.B1(n_954),
.B2(n_854),
.Y(n_4053)
);

AND2x4_ASAP7_75t_L g4054 ( 
.A(n_3191),
.B(n_3302),
.Y(n_4054)
);

BUFx3_ASAP7_75t_L g4055 ( 
.A(n_3191),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3330),
.Y(n_4056)
);

AND2x4_ASAP7_75t_L g4057 ( 
.A(n_3191),
.B(n_3064),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3422),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3116),
.B(n_3122),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3422),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3122),
.B(n_2466),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3211),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_3494),
.Y(n_4063)
);

INVx4_ASAP7_75t_L g4064 ( 
.A(n_3184),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_3514),
.B(n_2606),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_L g4066 ( 
.A(n_3514),
.B(n_2792),
.Y(n_4066)
);

BUFx3_ASAP7_75t_L g4067 ( 
.A(n_3302),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3343),
.B(n_2606),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3423),
.Y(n_4069)
);

AND2x6_ASAP7_75t_L g4070 ( 
.A(n_3100),
.B(n_2917),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3214),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3423),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3429),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_SL g4074 ( 
.A(n_3343),
.B(n_2864),
.Y(n_4074)
);

BUFx6f_ASAP7_75t_L g4075 ( 
.A(n_3184),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3429),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3430),
.Y(n_4077)
);

AND2x4_ASAP7_75t_L g4078 ( 
.A(n_3302),
.B(n_3064),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3430),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3711),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3609),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3719),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3610),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3721),
.B(n_3518),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3730),
.B(n_3290),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3613),
.Y(n_4086)
);

CKINVDCx20_ASAP7_75t_R g4087 ( 
.A(n_3784),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3615),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3727),
.Y(n_4089)
);

INVxp67_ASAP7_75t_L g4090 ( 
.A(n_3629),
.Y(n_4090)
);

AND2x2_ASAP7_75t_L g4091 ( 
.A(n_3701),
.B(n_3518),
.Y(n_4091)
);

O2A1O1Ixp5_ASAP7_75t_L g4092 ( 
.A1(n_3616),
.A2(n_3091),
.B(n_3108),
.C(n_3118),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3730),
.B(n_3684),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3617),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3742),
.Y(n_4095)
);

NAND2xp33_ASAP7_75t_L g4096 ( 
.A(n_3746),
.B(n_3515),
.Y(n_4096)
);

OR2x2_ASAP7_75t_L g4097 ( 
.A(n_3734),
.B(n_3524),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_3612),
.B(n_3524),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3620),
.Y(n_4099)
);

AOI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_4014),
.A2(n_2910),
.B1(n_2923),
.B2(n_2809),
.Y(n_4100)
);

AOI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_4014),
.A2(n_3652),
.B1(n_3636),
.B2(n_3926),
.Y(n_4101)
);

NOR2xp33_ASAP7_75t_SL g4102 ( 
.A(n_3678),
.B(n_2672),
.Y(n_4102)
);

NOR2xp33_ASAP7_75t_L g4103 ( 
.A(n_3616),
.B(n_1861),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3621),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3684),
.B(n_3290),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_L g4106 ( 
.A(n_3687),
.B(n_1865),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_3612),
.B(n_3525),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3757),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3624),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3627),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3815),
.B(n_3392),
.Y(n_4111)
);

AND2x2_ASAP7_75t_L g4112 ( 
.A(n_3842),
.B(n_3525),
.Y(n_4112)
);

BUFx4_ASAP7_75t_L g4113 ( 
.A(n_3901),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_SL g4114 ( 
.A(n_3815),
.B(n_3302),
.Y(n_4114)
);

INVx8_ASAP7_75t_L g4115 ( 
.A(n_3640),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3715),
.B(n_3290),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3632),
.Y(n_4117)
);

NOR2xp67_ASAP7_75t_SL g4118 ( 
.A(n_3628),
.B(n_2217),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_3687),
.B(n_3516),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_3734),
.B(n_3527),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_SL g4121 ( 
.A(n_3631),
.B(n_3636),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3715),
.B(n_3296),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3732),
.B(n_3668),
.Y(n_4123)
);

AND2x4_ASAP7_75t_L g4124 ( 
.A(n_4057),
.B(n_3527),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_SL g4125 ( 
.A(n_3652),
.B(n_3530),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3760),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3732),
.B(n_3296),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3635),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3637),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3619),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3641),
.Y(n_4131)
);

OR2x2_ASAP7_75t_L g4132 ( 
.A(n_3751),
.B(n_3530),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_SL g4133 ( 
.A(n_3668),
.B(n_3532),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3812),
.B(n_3296),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_4050),
.B(n_3532),
.Y(n_4135)
);

BUFx6f_ASAP7_75t_L g4136 ( 
.A(n_3651),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3938),
.B(n_3582),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_SL g4138 ( 
.A(n_4050),
.B(n_3535),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3647),
.Y(n_4139)
);

NOR2xp33_ASAP7_75t_L g4140 ( 
.A(n_3673),
.B(n_1877),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3938),
.B(n_3589),
.Y(n_4141)
);

OR2x2_ASAP7_75t_SL g4142 ( 
.A(n_3878),
.B(n_2217),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3688),
.Y(n_4143)
);

NOR2xp67_ASAP7_75t_L g4144 ( 
.A(n_3780),
.B(n_2864),
.Y(n_4144)
);

NOR2xp33_ASAP7_75t_L g4145 ( 
.A(n_3736),
.B(n_1877),
.Y(n_4145)
);

AND2x6_ASAP7_75t_L g4146 ( 
.A(n_4042),
.B(n_3100),
.Y(n_4146)
);

BUFx3_ASAP7_75t_L g4147 ( 
.A(n_3669),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3874),
.B(n_3535),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3626),
.B(n_3536),
.Y(n_4149)
);

NOR2xp33_ASAP7_75t_L g4150 ( 
.A(n_3720),
.B(n_1881),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3629),
.Y(n_4151)
);

NOR3xp33_ASAP7_75t_L g4152 ( 
.A(n_3888),
.B(n_2323),
.C(n_2298),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3648),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3926),
.B(n_3536),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_SL g4155 ( 
.A(n_4066),
.B(n_3538),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3650),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_3691),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_3661),
.B(n_1881),
.Y(n_4158)
);

INVx2_ASAP7_75t_SL g4159 ( 
.A(n_3681),
.Y(n_4159)
);

NOR2xp33_ASAP7_75t_L g4160 ( 
.A(n_3707),
.B(n_3849),
.Y(n_4160)
);

OAI22xp5_ASAP7_75t_L g4161 ( 
.A1(n_3654),
.A2(n_3343),
.B1(n_3574),
.B2(n_3313),
.Y(n_4161)
);

AOI22xp5_ASAP7_75t_L g4162 ( 
.A1(n_4030),
.A2(n_2923),
.B1(n_2910),
.B2(n_2041),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3707),
.B(n_3538),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_3672),
.A2(n_3260),
.B1(n_3292),
.B2(n_3251),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3611),
.B(n_3539),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3653),
.Y(n_4166)
);

NOR2xp33_ASAP7_75t_L g4167 ( 
.A(n_3751),
.B(n_1898),
.Y(n_4167)
);

OAI22xp33_ASAP7_75t_L g4168 ( 
.A1(n_4001),
.A2(n_2893),
.B1(n_2890),
.B2(n_2878),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3672),
.A2(n_3260),
.B1(n_3292),
.B2(n_3251),
.Y(n_4169)
);

INVx3_ASAP7_75t_L g4170 ( 
.A(n_4075),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_SL g4171 ( 
.A(n_4066),
.B(n_3539),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3695),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3655),
.Y(n_4173)
);

AOI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_4030),
.A2(n_2041),
.B1(n_2035),
.B2(n_1903),
.Y(n_4174)
);

INVx3_ASAP7_75t_L g4175 ( 
.A(n_4075),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3659),
.Y(n_4176)
);

AOI221xp5_ASAP7_75t_L g4177 ( 
.A1(n_3745),
.A2(n_1745),
.B1(n_1749),
.B2(n_1748),
.C(n_1742),
.Y(n_4177)
);

AOI22xp33_ASAP7_75t_L g4178 ( 
.A1(n_3792),
.A2(n_3335),
.B1(n_3337),
.B2(n_3308),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3706),
.B(n_3546),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3858),
.B(n_3546),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3858),
.B(n_3548),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_3702),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_SL g4183 ( 
.A(n_3638),
.B(n_3548),
.Y(n_4183)
);

INVx2_ASAP7_75t_SL g4184 ( 
.A(n_3638),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_R g4185 ( 
.A(n_3806),
.B(n_1898),
.Y(n_4185)
);

INVxp67_ASAP7_75t_L g4186 ( 
.A(n_3642),
.Y(n_4186)
);

NOR2xp33_ASAP7_75t_L g4187 ( 
.A(n_3788),
.B(n_1903),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3812),
.B(n_3297),
.Y(n_4188)
);

INVx2_ASAP7_75t_SL g4189 ( 
.A(n_3642),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3670),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_3712),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3713),
.Y(n_4192)
);

INVxp67_ASAP7_75t_L g4193 ( 
.A(n_3809),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_3725),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3729),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_3676),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_3792),
.A2(n_3335),
.B1(n_3337),
.B2(n_3308),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_SL g4198 ( 
.A(n_3788),
.B(n_3550),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_3738),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_L g4200 ( 
.A1(n_3907),
.A2(n_3395),
.B1(n_3411),
.B2(n_3340),
.Y(n_4200)
);

A2O1A1Ixp33_ASAP7_75t_L g4201 ( 
.A1(n_3747),
.A2(n_3574),
.B(n_3561),
.C(n_3503),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_3682),
.Y(n_4202)
);

NOR2xp33_ASAP7_75t_L g4203 ( 
.A(n_3771),
.B(n_1904),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3686),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_3744),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_3749),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3869),
.B(n_3550),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_3756),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_3683),
.B(n_3689),
.Y(n_4209)
);

OAI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_3745),
.A2(n_2893),
.B1(n_2890),
.B2(n_2878),
.Y(n_4210)
);

AO221x1_ASAP7_75t_L g4211 ( 
.A1(n_3872),
.A2(n_3132),
.B1(n_3577),
.B2(n_3492),
.C(n_3487),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3826),
.B(n_3297),
.Y(n_4212)
);

AOI22xp5_ASAP7_75t_L g4213 ( 
.A1(n_3771),
.A2(n_2035),
.B1(n_1921),
.B2(n_1922),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3826),
.B(n_3297),
.Y(n_4214)
);

BUFx4_ASAP7_75t_L g4215 ( 
.A(n_3692),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_3836),
.B(n_3299),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3694),
.Y(n_4217)
);

OR2x2_ASAP7_75t_L g4218 ( 
.A(n_3646),
.B(n_3562),
.Y(n_4218)
);

OR2x2_ASAP7_75t_L g4219 ( 
.A(n_3739),
.B(n_3562),
.Y(n_4219)
);

OAI22xp33_ASAP7_75t_L g4220 ( 
.A1(n_3723),
.A2(n_2889),
.B1(n_2865),
.B2(n_2680),
.Y(n_4220)
);

A2O1A1Ixp33_ASAP7_75t_L g4221 ( 
.A1(n_3869),
.A2(n_3879),
.B(n_3873),
.C(n_3660),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3696),
.Y(n_4222)
);

AOI22xp33_ASAP7_75t_L g4223 ( 
.A1(n_3907),
.A2(n_3395),
.B1(n_3411),
.B2(n_3340),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3703),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_3618),
.B(n_1904),
.Y(n_4225)
);

INVxp67_ASAP7_75t_SL g4226 ( 
.A(n_3649),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_3759),
.Y(n_4227)
);

NOR2xp33_ASAP7_75t_L g4228 ( 
.A(n_3873),
.B(n_1921),
.Y(n_4228)
);

AOI21xp5_ASAP7_75t_L g4229 ( 
.A1(n_3882),
.A2(n_3416),
.B(n_3607),
.Y(n_4229)
);

BUFx8_ASAP7_75t_L g4230 ( 
.A(n_3960),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3879),
.B(n_3566),
.Y(n_4231)
);

AOI22xp33_ASAP7_75t_L g4232 ( 
.A1(n_3872),
.A2(n_3501),
.B1(n_3506),
.B2(n_3498),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_SL g4233 ( 
.A(n_3743),
.B(n_3566),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_3778),
.B(n_3735),
.Y(n_4234)
);

OR2x2_ASAP7_75t_L g4235 ( 
.A(n_3685),
.B(n_3567),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_3762),
.Y(n_4236)
);

AOI22xp5_ASAP7_75t_L g4237 ( 
.A1(n_3780),
.A2(n_1923),
.B1(n_1925),
.B2(n_1922),
.Y(n_4237)
);

NAND3xp33_ASAP7_75t_L g4238 ( 
.A(n_3970),
.B(n_1748),
.C(n_1745),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_SL g4239 ( 
.A(n_3743),
.B(n_3567),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_3768),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3823),
.B(n_3568),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_SL g4242 ( 
.A(n_3942),
.B(n_3568),
.Y(n_4242)
);

AOI22xp33_ASAP7_75t_L g4243 ( 
.A1(n_3872),
.A2(n_3501),
.B1(n_3506),
.B2(n_3498),
.Y(n_4243)
);

NOR2xp33_ASAP7_75t_L g4244 ( 
.A(n_3831),
.B(n_1923),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_3823),
.B(n_3572),
.Y(n_4245)
);

BUFx5_ASAP7_75t_L g4246 ( 
.A(n_3862),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3705),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_3733),
.B(n_3572),
.Y(n_4248)
);

NOR2xp33_ASAP7_75t_L g4249 ( 
.A(n_3831),
.B(n_1925),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4048),
.B(n_3295),
.Y(n_4250)
);

NOR2x1p5_ASAP7_75t_L g4251 ( 
.A(n_3753),
.B(n_2865),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3708),
.Y(n_4252)
);

NOR2xp33_ASAP7_75t_L g4253 ( 
.A(n_3833),
.B(n_1935),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_3773),
.Y(n_4254)
);

OAI22xp33_ASAP7_75t_SL g4255 ( 
.A1(n_4044),
.A2(n_3133),
.B1(n_3165),
.B2(n_3128),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_3777),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3787),
.Y(n_4257)
);

NAND2xp33_ASAP7_75t_L g4258 ( 
.A(n_3746),
.B(n_3490),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_3836),
.B(n_3299),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_SL g4260 ( 
.A(n_3851),
.B(n_2889),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_3913),
.B(n_3299),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3913),
.B(n_3309),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3966),
.B(n_3309),
.Y(n_4263)
);

OAI22xp5_ASAP7_75t_L g4264 ( 
.A1(n_3654),
.A2(n_3966),
.B1(n_4039),
.B2(n_4033),
.Y(n_4264)
);

NOR2xp33_ASAP7_75t_L g4265 ( 
.A(n_3871),
.B(n_1935),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_3891),
.B(n_3590),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3786),
.B(n_3309),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3786),
.B(n_3122),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3790),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3798),
.B(n_3129),
.Y(n_4270)
);

AND2x4_ASAP7_75t_L g4271 ( 
.A(n_4057),
.B(n_3347),
.Y(n_4271)
);

BUFx6f_ASAP7_75t_SL g4272 ( 
.A(n_3625),
.Y(n_4272)
);

INVx2_ASAP7_75t_SL g4273 ( 
.A(n_3710),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3800),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_SL g4275 ( 
.A(n_3978),
.B(n_3168),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_3798),
.B(n_3129),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_3779),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4065),
.B(n_3590),
.Y(n_4278)
);

INVxp67_ASAP7_75t_SL g4279 ( 
.A(n_3649),
.Y(n_4279)
);

AND2x4_ASAP7_75t_L g4280 ( 
.A(n_4078),
.B(n_3752),
.Y(n_4280)
);

O2A1O1Ixp5_ASAP7_75t_L g4281 ( 
.A1(n_3770),
.A2(n_3200),
.B(n_3207),
.C(n_3180),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3804),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3808),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4042),
.B(n_3594),
.Y(n_4284)
);

NAND3xp33_ASAP7_75t_L g4285 ( 
.A(n_3974),
.B(n_1760),
.C(n_1749),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4078),
.B(n_3594),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_3824),
.B(n_3129),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_SL g4288 ( 
.A(n_3978),
.B(n_3210),
.Y(n_4288)
);

O2A1O1Ixp33_ASAP7_75t_L g4289 ( 
.A1(n_3718),
.A2(n_3396),
.B(n_3213),
.C(n_3222),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_3810),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_3740),
.B(n_3600),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_SL g4292 ( 
.A(n_3992),
.B(n_3216),
.Y(n_4292)
);

NOR2xp33_ASAP7_75t_L g4293 ( 
.A(n_3992),
.B(n_1945),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_3782),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_L g4295 ( 
.A(n_4020),
.B(n_1945),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3824),
.B(n_3838),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3838),
.B(n_3173),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_3811),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3817),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4039),
.A2(n_3574),
.B1(n_3314),
.B2(n_3132),
.Y(n_4300)
);

NOR2xp33_ASAP7_75t_SL g4301 ( 
.A(n_3700),
.B(n_2679),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_3835),
.B(n_3840),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_3846),
.B(n_3173),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3820),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_3651),
.Y(n_4305)
);

INVxp67_ASAP7_75t_L g4306 ( 
.A(n_3622),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_3857),
.B(n_3173),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3825),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_3863),
.B(n_3178),
.Y(n_4309)
);

BUFx2_ASAP7_75t_L g4310 ( 
.A(n_3645),
.Y(n_4310)
);

NAND2xp33_ASAP7_75t_L g4311 ( 
.A(n_3746),
.B(n_3490),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_3867),
.B(n_3178),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3870),
.Y(n_4313)
);

INVx2_ASAP7_75t_SL g4314 ( 
.A(n_3716),
.Y(n_4314)
);

NOR3xp33_ASAP7_75t_L g4315 ( 
.A(n_3974),
.B(n_3250),
.C(n_3231),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3877),
.Y(n_4316)
);

BUFx5_ASAP7_75t_L g4317 ( 
.A(n_3862),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3883),
.Y(n_4318)
);

INVx5_ASAP7_75t_L g4319 ( 
.A(n_3862),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_SL g4320 ( 
.A(n_4020),
.B(n_3255),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3885),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_SL g4322 ( 
.A(n_3634),
.B(n_3264),
.Y(n_4322)
);

NOR2xp33_ASAP7_75t_L g4323 ( 
.A(n_3658),
.B(n_1949),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3886),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_3898),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_3666),
.B(n_3288),
.Y(n_4326)
);

INVx3_ASAP7_75t_L g4327 ( 
.A(n_4075),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_3903),
.B(n_3178),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3904),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3972),
.B(n_3600),
.Y(n_4330)
);

OR2x6_ASAP7_75t_L g4331 ( 
.A(n_3640),
.B(n_3194),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3972),
.B(n_3608),
.Y(n_4332)
);

AOI22xp33_ASAP7_75t_L g4333 ( 
.A1(n_3699),
.A2(n_3438),
.B1(n_3448),
.B2(n_3446),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_3699),
.B(n_3608),
.Y(n_4334)
);

BUFx6f_ASAP7_75t_L g4335 ( 
.A(n_3651),
.Y(n_4335)
);

OAI22xp5_ASAP7_75t_SL g4336 ( 
.A1(n_3899),
.A2(n_2939),
.B1(n_2934),
.B2(n_2719),
.Y(n_4336)
);

INVxp67_ASAP7_75t_L g4337 ( 
.A(n_3726),
.Y(n_4337)
);

NOR2xp67_ASAP7_75t_L g4338 ( 
.A(n_4041),
.B(n_2679),
.Y(n_4338)
);

INVx2_ASAP7_75t_SL g4339 ( 
.A(n_3750),
.Y(n_4339)
);

NOR2x1p5_ASAP7_75t_L g4340 ( 
.A(n_3677),
.B(n_2680),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_SL g4341 ( 
.A(n_3671),
.B(n_3723),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_3783),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_3789),
.Y(n_4343)
);

AND2x4_ASAP7_75t_L g4344 ( 
.A(n_3752),
.B(n_4054),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_4016),
.B(n_1949),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3916),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_3791),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_3776),
.A2(n_3438),
.B1(n_3448),
.B2(n_3446),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_3807),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_3917),
.Y(n_4350)
);

BUFx2_ASAP7_75t_L g4351 ( 
.A(n_3989),
.Y(n_4351)
);

BUFx5_ASAP7_75t_L g4352 ( 
.A(n_3862),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_3814),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_3844),
.B(n_3486),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_L g4355 ( 
.A(n_3987),
.B(n_1954),
.Y(n_4355)
);

INVxp67_ASAP7_75t_L g4356 ( 
.A(n_4036),
.Y(n_4356)
);

NOR2xp67_ASAP7_75t_L g4357 ( 
.A(n_3987),
.B(n_2685),
.Y(n_4357)
);

INVx1_ASAP7_75t_SL g4358 ( 
.A(n_3845),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_3829),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3918),
.Y(n_4360)
);

NOR2xp33_ASAP7_75t_L g4361 ( 
.A(n_3900),
.B(n_1954),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_3830),
.Y(n_4362)
);

NOR3xp33_ASAP7_75t_L g4363 ( 
.A(n_3958),
.B(n_3289),
.C(n_2690),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_3919),
.B(n_3179),
.Y(n_4364)
);

AND2x6_ASAP7_75t_SL g4365 ( 
.A(n_3958),
.B(n_2838),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_3921),
.B(n_3179),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_3933),
.B(n_3179),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3944),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_3952),
.B(n_3181),
.Y(n_4369)
);

INVx2_ASAP7_75t_SL g4370 ( 
.A(n_4019),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_3956),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_3837),
.Y(n_4372)
);

NAND3xp33_ASAP7_75t_L g4373 ( 
.A(n_3963),
.B(n_1766),
.C(n_1761),
.Y(n_4373)
);

NAND2xp33_ASAP7_75t_L g4374 ( 
.A(n_3746),
.B(n_3490),
.Y(n_4374)
);

INVx2_ASAP7_75t_SL g4375 ( 
.A(n_3625),
.Y(n_4375)
);

AOI22xp5_ASAP7_75t_L g4376 ( 
.A1(n_3737),
.A2(n_1967),
.B1(n_1960),
.B2(n_2852),
.Y(n_4376)
);

BUFx6f_ASAP7_75t_L g4377 ( 
.A(n_3674),
.Y(n_4377)
);

INVxp67_ASAP7_75t_R g4378 ( 
.A(n_3985),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_3957),
.B(n_3962),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_3963),
.A2(n_1967),
.B1(n_1960),
.B2(n_2852),
.Y(n_4380)
);

BUFx3_ASAP7_75t_L g4381 ( 
.A(n_3692),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_3973),
.B(n_3980),
.Y(n_4382)
);

NOR2xp33_ASAP7_75t_L g4383 ( 
.A(n_3776),
.B(n_2712),
.Y(n_4383)
);

INVxp33_ASAP7_75t_L g4384 ( 
.A(n_3828),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_3982),
.B(n_3181),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_3843),
.Y(n_4386)
);

BUFx3_ASAP7_75t_L g4387 ( 
.A(n_3693),
.Y(n_4387)
);

INVxp67_ASAP7_75t_SL g4388 ( 
.A(n_3766),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_3828),
.B(n_3486),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_SL g4390 ( 
.A(n_3822),
.B(n_2690),
.Y(n_4390)
);

INVxp33_ASAP7_75t_SL g4391 ( 
.A(n_3755),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_3993),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_3855),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_3995),
.B(n_3181),
.Y(n_4394)
);

NOR2xp33_ASAP7_75t_L g4395 ( 
.A(n_3839),
.B(n_2719),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4005),
.B(n_3183),
.Y(n_4396)
);

NOR3xp33_ASAP7_75t_L g4397 ( 
.A(n_3797),
.B(n_2694),
.C(n_2685),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_3856),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_4011),
.B(n_3183),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_3839),
.B(n_3844),
.Y(n_4400)
);

INVx2_ASAP7_75t_SL g4401 ( 
.A(n_4038),
.Y(n_4401)
);

INVx2_ASAP7_75t_L g4402 ( 
.A(n_3893),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4017),
.B(n_3183),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_SL g4404 ( 
.A(n_3822),
.B(n_4054),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_SL g4405 ( 
.A(n_4000),
.B(n_2694),
.Y(n_4405)
);

NOR2xp33_ASAP7_75t_L g4406 ( 
.A(n_3774),
.B(n_2853),
.Y(n_4406)
);

NOR2xp33_ASAP7_75t_L g4407 ( 
.A(n_3774),
.B(n_2853),
.Y(n_4407)
);

HB1xp67_ASAP7_75t_L g4408 ( 
.A(n_3674),
.Y(n_4408)
);

INVx3_ASAP7_75t_L g4409 ( 
.A(n_4018),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_SL g4410 ( 
.A(n_4000),
.B(n_2848),
.Y(n_4410)
);

BUFx4f_ASAP7_75t_L g4411 ( 
.A(n_3746),
.Y(n_4411)
);

AOI22xp33_ASAP7_75t_L g4412 ( 
.A1(n_4051),
.A2(n_3657),
.B1(n_3630),
.B2(n_3911),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_3630),
.B(n_3449),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_L g4414 ( 
.A1(n_3657),
.A2(n_3455),
.B1(n_3457),
.B2(n_3449),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4023),
.Y(n_4415)
);

INVxp33_ASAP7_75t_L g4416 ( 
.A(n_3769),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_3894),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_3931),
.B(n_2848),
.Y(n_4418)
);

NAND2xp33_ASAP7_75t_SL g4419 ( 
.A(n_4018),
.B(n_2858),
.Y(n_4419)
);

BUFx8_ASAP7_75t_L g4420 ( 
.A(n_3960),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_3905),
.Y(n_4421)
);

AOI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4040),
.A2(n_3457),
.B1(n_3459),
.B2(n_3455),
.Y(n_4422)
);

BUFx6f_ASAP7_75t_L g4423 ( 
.A(n_3674),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4024),
.Y(n_4424)
);

NAND2xp33_ASAP7_75t_L g4425 ( 
.A(n_3754),
.B(n_3490),
.Y(n_4425)
);

AND2x4_ASAP7_75t_L g4426 ( 
.A(n_4055),
.B(n_3347),
.Y(n_4426)
);

AOI22x1_ASAP7_75t_L g4427 ( 
.A1(n_3665),
.A2(n_3384),
.B1(n_3388),
.B2(n_3383),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_SL g4428 ( 
.A(n_3931),
.B(n_2858),
.Y(n_4428)
);

NOR2xp33_ASAP7_75t_L g4429 ( 
.A(n_3939),
.B(n_2867),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4033),
.B(n_3459),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_4067),
.B(n_3347),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_3766),
.B(n_3454),
.Y(n_4432)
);

INVx2_ASAP7_75t_SL g4433 ( 
.A(n_4038),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_3934),
.B(n_2441),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_3775),
.B(n_3462),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4026),
.Y(n_4436)
);

NAND2xp33_ASAP7_75t_SL g4437 ( 
.A(n_4064),
.B(n_4027),
.Y(n_4437)
);

AOI22xp33_ASAP7_75t_L g4438 ( 
.A1(n_3664),
.A2(n_3347),
.B1(n_3552),
.B2(n_3447),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4029),
.B(n_3185),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_3758),
.B(n_2867),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4034),
.B(n_3185),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4052),
.B(n_3185),
.Y(n_4442)
);

INVx1_ASAP7_75t_SL g4443 ( 
.A(n_3852),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_3664),
.B(n_3383),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_3664),
.B(n_3384),
.Y(n_4445)
);

INVxp67_ASAP7_75t_SL g4446 ( 
.A(n_3775),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4056),
.B(n_4059),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4059),
.B(n_3224),
.Y(n_4448)
);

NOR3xp33_ASAP7_75t_L g4449 ( 
.A(n_3994),
.B(n_1772),
.C(n_1768),
.Y(n_4449)
);

OR2x6_ASAP7_75t_L g4450 ( 
.A(n_3640),
.B(n_3194),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4058),
.Y(n_4451)
);

INVxp67_ASAP7_75t_L g4452 ( 
.A(n_3813),
.Y(n_4452)
);

NAND2xp33_ASAP7_75t_L g4453 ( 
.A(n_3754),
.B(n_3490),
.Y(n_4453)
);

NOR2xp33_ASAP7_75t_L g4454 ( 
.A(n_3758),
.B(n_2873),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_3929),
.Y(n_4455)
);

AOI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4037),
.A2(n_3607),
.B(n_3490),
.Y(n_4456)
);

O2A1O1Ixp33_ASAP7_75t_L g4457 ( 
.A1(n_3718),
.A2(n_3526),
.B(n_3555),
.C(n_3554),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4060),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_SL g4459 ( 
.A(n_3934),
.B(n_2441),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4069),
.B(n_3224),
.Y(n_4460)
);

INVx2_ASAP7_75t_L g4461 ( 
.A(n_3945),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_SL g4462 ( 
.A(n_4064),
.B(n_2441),
.Y(n_4462)
);

AOI21xp5_ASAP7_75t_L g4463 ( 
.A1(n_3639),
.A2(n_3607),
.B(n_3323),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4072),
.B(n_3225),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_SL g4465 ( 
.A(n_3633),
.B(n_2807),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_3954),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_SL g4467 ( 
.A(n_3633),
.B(n_2807),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4073),
.B(n_3225),
.Y(n_4468)
);

INVx2_ASAP7_75t_SL g4469 ( 
.A(n_3912),
.Y(n_4469)
);

NOR2xp33_ASAP7_75t_L g4470 ( 
.A(n_3834),
.B(n_2873),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4076),
.B(n_3109),
.Y(n_4471)
);

AND2x4_ASAP7_75t_L g4472 ( 
.A(n_3644),
.B(n_3763),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4077),
.B(n_3109),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4079),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_3965),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4028),
.B(n_3109),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_3660),
.B(n_3680),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_3977),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_SL g4479 ( 
.A(n_3680),
.B(n_2812),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_SL g4480 ( 
.A(n_3680),
.B(n_2812),
.Y(n_4480)
);

HB1xp67_ASAP7_75t_L g4481 ( 
.A(n_3793),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4028),
.B(n_3100),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_3983),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_4031),
.B(n_3109),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_R g4485 ( 
.A(n_3861),
.B(n_2747),
.Y(n_4485)
);

INVxp67_ASAP7_75t_SL g4486 ( 
.A(n_3667),
.Y(n_4486)
);

BUFx3_ASAP7_75t_L g4487 ( 
.A(n_3769),
.Y(n_4487)
);

HB1xp67_ASAP7_75t_L g4488 ( 
.A(n_4090),
.Y(n_4488)
);

AND2x4_ASAP7_75t_L g4489 ( 
.A(n_4472),
.B(n_3643),
.Y(n_4489)
);

INVxp67_ASAP7_75t_SL g4490 ( 
.A(n_4226),
.Y(n_4490)
);

INVx4_ASAP7_75t_L g4491 ( 
.A(n_4319),
.Y(n_4491)
);

OR2x2_ASAP7_75t_L g4492 ( 
.A(n_4123),
.B(n_3596),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4080),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4123),
.B(n_3665),
.Y(n_4494)
);

BUFx3_ASAP7_75t_L g4495 ( 
.A(n_4147),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4427),
.Y(n_4496)
);

AND2x2_ASAP7_75t_SL g4497 ( 
.A(n_4411),
.B(n_3909),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4082),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_4089),
.Y(n_4499)
);

OAI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_4160),
.A2(n_3521),
.B(n_3329),
.Y(n_4500)
);

INVx2_ASAP7_75t_L g4501 ( 
.A(n_4095),
.Y(n_4501)
);

OAI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_4221),
.A2(n_3317),
.B(n_3483),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_4098),
.B(n_1768),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4107),
.B(n_3665),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4154),
.B(n_3447),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_4103),
.B(n_1772),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4101),
.B(n_4163),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4084),
.B(n_4091),
.Y(n_4508)
);

BUFx6f_ASAP7_75t_L g4509 ( 
.A(n_4319),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4093),
.B(n_3447),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4302),
.Y(n_4511)
);

BUFx6f_ASAP7_75t_L g4512 ( 
.A(n_4319),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_4108),
.Y(n_4513)
);

INVx2_ASAP7_75t_SL g4514 ( 
.A(n_4136),
.Y(n_4514)
);

INVx4_ASAP7_75t_L g4515 ( 
.A(n_4319),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4093),
.B(n_3314),
.Y(n_4516)
);

AND2x2_ASAP7_75t_L g4517 ( 
.A(n_4278),
.B(n_3984),
.Y(n_4517)
);

BUFx3_ASAP7_75t_L g4518 ( 
.A(n_4351),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4137),
.B(n_3754),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4141),
.B(n_3754),
.Y(n_4520)
);

AND2x2_ASAP7_75t_L g4521 ( 
.A(n_4126),
.B(n_3997),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4303),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4081),
.Y(n_4523)
);

BUFx6f_ASAP7_75t_L g4524 ( 
.A(n_4411),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4444),
.B(n_4025),
.Y(n_4525)
);

CKINVDCx20_ASAP7_75t_R g4526 ( 
.A(n_4087),
.Y(n_4526)
);

BUFx3_ASAP7_75t_L g4527 ( 
.A(n_4310),
.Y(n_4527)
);

BUFx3_ASAP7_75t_L g4528 ( 
.A(n_4387),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4112),
.B(n_3754),
.Y(n_4529)
);

INVx1_ASAP7_75t_SL g4530 ( 
.A(n_4151),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4303),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4445),
.B(n_4062),
.Y(n_4532)
);

AND2x4_ASAP7_75t_L g4533 ( 
.A(n_4472),
.B(n_3643),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4302),
.Y(n_4534)
);

BUFx3_ASAP7_75t_L g4535 ( 
.A(n_4136),
.Y(n_4535)
);

AOI22xp5_ASAP7_75t_L g4536 ( 
.A1(n_4203),
.A2(n_2747),
.B1(n_2149),
.B2(n_2145),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4388),
.B(n_4446),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4083),
.Y(n_4538)
);

AND2x4_ASAP7_75t_L g4539 ( 
.A(n_4426),
.B(n_3663),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4180),
.B(n_4071),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4181),
.B(n_3388),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4086),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4307),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4088),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4207),
.B(n_3390),
.Y(n_4545)
);

BUFx2_ASAP7_75t_L g4546 ( 
.A(n_4279),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4231),
.B(n_3390),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4094),
.Y(n_4548)
);

NOR2xp33_ASAP7_75t_L g4549 ( 
.A(n_4228),
.B(n_2838),
.Y(n_4549)
);

NOR2xp33_ASAP7_75t_L g4550 ( 
.A(n_4106),
.B(n_2627),
.Y(n_4550)
);

OAI21xp5_ASAP7_75t_L g4551 ( 
.A1(n_4121),
.A2(n_3483),
.B(n_3405),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4148),
.B(n_4021),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4271),
.B(n_3394),
.Y(n_4553)
);

NAND2x1p5_ASAP7_75t_L g4554 ( 
.A(n_4477),
.B(n_4046),
.Y(n_4554)
);

OR2x2_ASAP7_75t_L g4555 ( 
.A(n_4330),
.B(n_3596),
.Y(n_4555)
);

INVxp67_ASAP7_75t_L g4556 ( 
.A(n_4184),
.Y(n_4556)
);

INVx2_ASAP7_75t_SL g4557 ( 
.A(n_4136),
.Y(n_4557)
);

INVx2_ASAP7_75t_SL g4558 ( 
.A(n_4305),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_4271),
.B(n_3394),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4379),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4209),
.B(n_3401),
.Y(n_4561)
);

BUFx6f_ASAP7_75t_L g4562 ( 
.A(n_4115),
.Y(n_4562)
);

BUFx3_ASAP7_75t_L g4563 ( 
.A(n_4305),
.Y(n_4563)
);

INVxp67_ASAP7_75t_SL g4564 ( 
.A(n_4097),
.Y(n_4564)
);

INVx3_ASAP7_75t_L g4565 ( 
.A(n_4331),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4307),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4309),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4332),
.B(n_3401),
.Y(n_4568)
);

INVxp67_ASAP7_75t_L g4569 ( 
.A(n_4189),
.Y(n_4569)
);

BUFx3_ASAP7_75t_L g4570 ( 
.A(n_4305),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4379),
.Y(n_4571)
);

BUFx6f_ASAP7_75t_L g4572 ( 
.A(n_4115),
.Y(n_4572)
);

INVx2_ASAP7_75t_SL g4573 ( 
.A(n_4335),
.Y(n_4573)
);

NOR2xp33_ASAP7_75t_L g4574 ( 
.A(n_4355),
.B(n_2632),
.Y(n_4574)
);

OAI21xp5_ASAP7_75t_L g4575 ( 
.A1(n_4092),
.A2(n_3543),
.B(n_3541),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4099),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4120),
.B(n_3644),
.Y(n_4577)
);

INVx2_ASAP7_75t_L g4578 ( 
.A(n_4309),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4312),
.Y(n_4579)
);

NOR2xp67_ASAP7_75t_R g4580 ( 
.A(n_4381),
.B(n_2217),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4451),
.B(n_3404),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4266),
.B(n_3644),
.Y(n_4582)
);

OAI21xp33_ASAP7_75t_L g4583 ( 
.A1(n_4140),
.A2(n_2464),
.B(n_2816),
.Y(n_4583)
);

BUFx3_ASAP7_75t_L g4584 ( 
.A(n_4335),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4382),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4234),
.B(n_3763),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4458),
.B(n_3404),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4218),
.B(n_3763),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4248),
.B(n_3410),
.Y(n_4589)
);

AND2x2_ASAP7_75t_L g4590 ( 
.A(n_4474),
.B(n_3410),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4232),
.B(n_3412),
.Y(n_4591)
);

INVx3_ASAP7_75t_L g4592 ( 
.A(n_4331),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4243),
.B(n_3412),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4312),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_SL g4595 ( 
.A(n_4158),
.B(n_3802),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4104),
.B(n_3420),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4328),
.Y(n_4597)
);

NAND2x1p5_ASAP7_75t_L g4598 ( 
.A(n_4119),
.B(n_4046),
.Y(n_4598)
);

BUFx6f_ASAP7_75t_L g4599 ( 
.A(n_4115),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4109),
.B(n_3420),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4110),
.B(n_3377),
.Y(n_4601)
);

NOR2xp33_ASAP7_75t_L g4602 ( 
.A(n_4167),
.B(n_2613),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4117),
.B(n_3377),
.Y(n_4603)
);

BUFx6f_ASAP7_75t_L g4604 ( 
.A(n_4331),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4382),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4328),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4132),
.B(n_4286),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4124),
.B(n_3014),
.Y(n_4608)
);

BUFx6f_ASAP7_75t_L g4609 ( 
.A(n_4450),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4364),
.Y(n_4610)
);

BUFx3_ASAP7_75t_L g4611 ( 
.A(n_4335),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4128),
.B(n_3380),
.Y(n_4612)
);

BUFx4f_ASAP7_75t_L g4613 ( 
.A(n_4450),
.Y(n_4613)
);

INVx2_ASAP7_75t_SL g4614 ( 
.A(n_4377),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4129),
.B(n_4131),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4124),
.B(n_3793),
.Y(n_4616)
);

BUFx2_ASAP7_75t_L g4617 ( 
.A(n_4146),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4389),
.B(n_4135),
.Y(n_4618)
);

OAI21x1_ASAP7_75t_L g4619 ( 
.A1(n_4463),
.A2(n_3237),
.B(n_3576),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4364),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4366),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4138),
.B(n_3793),
.Y(n_4622)
);

BUFx3_ASAP7_75t_L g4623 ( 
.A(n_4377),
.Y(n_4623)
);

NAND2x1p5_ASAP7_75t_L g4624 ( 
.A(n_4404),
.B(n_4046),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4155),
.B(n_3795),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4139),
.B(n_3380),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4171),
.B(n_3795),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4153),
.B(n_3386),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4366),
.Y(n_4629)
);

INVx3_ASAP7_75t_L g4630 ( 
.A(n_4450),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4156),
.B(n_3386),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4166),
.B(n_3398),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4149),
.B(n_3795),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4173),
.B(n_3398),
.Y(n_4634)
);

BUFx6f_ASAP7_75t_L g4635 ( 
.A(n_4426),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4145),
.B(n_3799),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4176),
.B(n_3402),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_SL g4638 ( 
.A(n_4244),
.B(n_3802),
.Y(n_4638)
);

INVx2_ASAP7_75t_L g4639 ( 
.A(n_4367),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4190),
.B(n_3402),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_4334),
.B(n_3799),
.Y(n_4641)
);

BUFx6f_ASAP7_75t_L g4642 ( 
.A(n_4431),
.Y(n_4642)
);

BUFx3_ASAP7_75t_L g4643 ( 
.A(n_4377),
.Y(n_4643)
);

HB1xp67_ASAP7_75t_L g4644 ( 
.A(n_4186),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_4185),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4367),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4369),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4361),
.B(n_3799),
.Y(n_4648)
);

INVx3_ASAP7_75t_L g4649 ( 
.A(n_4246),
.Y(n_4649)
);

INVx4_ASAP7_75t_L g4650 ( 
.A(n_4423),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4241),
.B(n_4074),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4196),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4202),
.B(n_3407),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4369),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4204),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4245),
.B(n_4400),
.Y(n_4656)
);

NOR2xp33_ASAP7_75t_L g4657 ( 
.A(n_4187),
.B(n_2613),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4217),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4222),
.B(n_3407),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4125),
.B(n_3409),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4224),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4413),
.B(n_3409),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_SL g4663 ( 
.A(n_4249),
.B(n_2816),
.Y(n_4663)
);

AND2x2_ASAP7_75t_SL g4664 ( 
.A(n_4258),
.B(n_3909),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4247),
.B(n_3415),
.Y(n_4665)
);

OR2x2_ASAP7_75t_SL g4666 ( 
.A(n_4373),
.B(n_3841),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4385),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4252),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4475),
.B(n_4478),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4130),
.B(n_3415),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4254),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4385),
.Y(n_4672)
);

INVx3_ASAP7_75t_L g4673 ( 
.A(n_4246),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4394),
.Y(n_4674)
);

NAND2xp5_ASAP7_75t_L g4675 ( 
.A(n_4114),
.B(n_4193),
.Y(n_4675)
);

OAI21xp5_ASAP7_75t_L g4676 ( 
.A1(n_4281),
.A2(n_3557),
.B(n_3544),
.Y(n_4676)
);

INVx3_ASAP7_75t_L g4677 ( 
.A(n_4246),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4394),
.Y(n_4678)
);

BUFx6f_ASAP7_75t_L g4679 ( 
.A(n_4431),
.Y(n_4679)
);

NOR2xp33_ASAP7_75t_L g4680 ( 
.A(n_4345),
.B(n_2615),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4256),
.Y(n_4681)
);

BUFx6f_ASAP7_75t_L g4682 ( 
.A(n_4423),
.Y(n_4682)
);

BUFx6f_ASAP7_75t_L g4683 ( 
.A(n_4423),
.Y(n_4683)
);

BUFx3_ASAP7_75t_L g4684 ( 
.A(n_4273),
.Y(n_4684)
);

HB1xp67_ASAP7_75t_L g4685 ( 
.A(n_4235),
.Y(n_4685)
);

AND2x2_ASAP7_75t_L g4686 ( 
.A(n_4143),
.B(n_4157),
.Y(n_4686)
);

AND2x4_ASAP7_75t_L g4687 ( 
.A(n_4409),
.B(n_3663),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4172),
.B(n_3552),
.Y(n_4688)
);

OR2x2_ASAP7_75t_SL g4689 ( 
.A(n_4285),
.B(n_3841),
.Y(n_4689)
);

INVx6_ASAP7_75t_L g4690 ( 
.A(n_4344),
.Y(n_4690)
);

AND2x2_ASAP7_75t_SL g4691 ( 
.A(n_4311),
.B(n_3827),
.Y(n_4691)
);

HB1xp67_ASAP7_75t_L g4692 ( 
.A(n_4291),
.Y(n_4692)
);

BUFx6f_ASAP7_75t_L g4693 ( 
.A(n_4146),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4182),
.B(n_3552),
.Y(n_4694)
);

CKINVDCx8_ASAP7_75t_R g4695 ( 
.A(n_4365),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4396),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_SL g4697 ( 
.A(n_4210),
.B(n_4357),
.Y(n_4697)
);

INVxp67_ASAP7_75t_L g4698 ( 
.A(n_4293),
.Y(n_4698)
);

INVx2_ASAP7_75t_L g4699 ( 
.A(n_4396),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_SL g4700 ( 
.A(n_4237),
.B(n_2822),
.Y(n_4700)
);

AND2x4_ASAP7_75t_L g4701 ( 
.A(n_4409),
.B(n_3690),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4354),
.B(n_4068),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4399),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4257),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4233),
.B(n_2470),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4269),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4399),
.Y(n_4707)
);

AND2x2_ASAP7_75t_SL g4708 ( 
.A(n_4374),
.B(n_3690),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4191),
.B(n_3552),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4403),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4403),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4274),
.Y(n_4712)
);

AND2x2_ASAP7_75t_SL g4713 ( 
.A(n_4425),
.B(n_3698),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4192),
.B(n_3552),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4194),
.B(n_4006),
.Y(n_4715)
);

NOR2xp33_ASAP7_75t_L g4716 ( 
.A(n_4295),
.B(n_2615),
.Y(n_4716)
);

INVx1_ASAP7_75t_SL g4717 ( 
.A(n_4358),
.Y(n_4717)
);

INVx3_ASAP7_75t_L g4718 ( 
.A(n_4246),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4439),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4439),
.Y(n_4720)
);

NOR2xp33_ASAP7_75t_L g4721 ( 
.A(n_4225),
.B(n_2633),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_4441),
.Y(n_4722)
);

AND2x2_ASAP7_75t_L g4723 ( 
.A(n_4195),
.B(n_4006),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4441),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4442),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_L g4726 ( 
.A(n_4239),
.B(n_2470),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4152),
.B(n_2470),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4159),
.Y(n_4728)
);

BUFx2_ASAP7_75t_L g4729 ( 
.A(n_4146),
.Y(n_4729)
);

INVx1_ASAP7_75t_SL g4730 ( 
.A(n_4443),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4133),
.B(n_3442),
.Y(n_4731)
);

NAND2x1p5_ASAP7_75t_L g4732 ( 
.A(n_4242),
.B(n_4046),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_SL g4733 ( 
.A(n_4174),
.B(n_2822),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4219),
.B(n_3450),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4198),
.B(n_3493),
.Y(n_4735)
);

AND2x4_ASAP7_75t_L g4736 ( 
.A(n_4280),
.B(n_3698),
.Y(n_4736)
);

INVx3_ASAP7_75t_L g4737 ( 
.A(n_4246),
.Y(n_4737)
);

INVx2_ASAP7_75t_L g4738 ( 
.A(n_4442),
.Y(n_4738)
);

AND2x2_ASAP7_75t_SL g4739 ( 
.A(n_4453),
.B(n_4053),
.Y(n_4739)
);

INVx3_ASAP7_75t_L g4740 ( 
.A(n_4246),
.Y(n_4740)
);

INVx3_ASAP7_75t_L g4741 ( 
.A(n_4317),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4199),
.B(n_4053),
.Y(n_4742)
);

BUFx2_ASAP7_75t_L g4743 ( 
.A(n_4146),
.Y(n_4743)
);

NOR2xp33_ASAP7_75t_L g4744 ( 
.A(n_4213),
.B(n_2633),
.Y(n_4744)
);

AND2x2_ASAP7_75t_SL g4745 ( 
.A(n_4438),
.B(n_3914),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4460),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4460),
.Y(n_4747)
);

INVx2_ASAP7_75t_L g4748 ( 
.A(n_4464),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4205),
.B(n_3596),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4464),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4206),
.B(n_3599),
.Y(n_4751)
);

BUFx3_ASAP7_75t_L g4752 ( 
.A(n_4314),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4208),
.B(n_3599),
.Y(n_4753)
);

BUFx6f_ASAP7_75t_L g4754 ( 
.A(n_4146),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4356),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_4468),
.Y(n_4756)
);

NOR2xp33_ASAP7_75t_R g4757 ( 
.A(n_4419),
.B(n_3704),
.Y(n_4757)
);

NOR2xp33_ASAP7_75t_L g4758 ( 
.A(n_4323),
.B(n_2643),
.Y(n_4758)
);

HB1xp67_ASAP7_75t_L g4759 ( 
.A(n_4306),
.Y(n_4759)
);

BUFx8_ASAP7_75t_L g4760 ( 
.A(n_4272),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4250),
.B(n_3717),
.Y(n_4761)
);

OAI21xp5_ASAP7_75t_L g4762 ( 
.A1(n_4238),
.A2(n_3583),
.B(n_3579),
.Y(n_4762)
);

OAI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4111),
.A2(n_3603),
.B(n_3601),
.Y(n_4763)
);

AND2x4_ASAP7_75t_L g4764 ( 
.A(n_4280),
.B(n_3868),
.Y(n_4764)
);

OR2x6_ASAP7_75t_L g4765 ( 
.A(n_4300),
.B(n_3868),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4282),
.Y(n_4766)
);

HB1xp67_ASAP7_75t_L g4767 ( 
.A(n_4408),
.Y(n_4767)
);

AND2x2_ASAP7_75t_SL g4768 ( 
.A(n_4406),
.B(n_4407),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4384),
.B(n_3717),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4283),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4227),
.B(n_3599),
.Y(n_4771)
);

OAI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4289),
.A2(n_3393),
.B(n_3387),
.Y(n_4772)
);

BUFx3_ASAP7_75t_L g4773 ( 
.A(n_4339),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4363),
.B(n_3906),
.Y(n_4774)
);

NOR2xp33_ASAP7_75t_R g4775 ( 
.A(n_4437),
.B(n_2779),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4468),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4236),
.Y(n_4777)
);

AND2x2_ASAP7_75t_L g4778 ( 
.A(n_4240),
.B(n_3602),
.Y(n_4778)
);

HB1xp67_ASAP7_75t_L g4779 ( 
.A(n_4481),
.Y(n_4779)
);

HB1xp67_ASAP7_75t_L g4780 ( 
.A(n_4337),
.Y(n_4780)
);

BUFx3_ASAP7_75t_L g4781 ( 
.A(n_4170),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_4277),
.B(n_3602),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4294),
.B(n_4342),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4343),
.B(n_3602),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4347),
.Y(n_4785)
);

AND2x2_ASAP7_75t_SL g4786 ( 
.A(n_4096),
.B(n_3914),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4290),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4183),
.B(n_4253),
.Y(n_4788)
);

NOR2xp33_ASAP7_75t_L g4789 ( 
.A(n_4265),
.B(n_2643),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4298),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_SL g4791 ( 
.A(n_4376),
.B(n_2826),
.Y(n_4791)
);

AND2x2_ASAP7_75t_L g4792 ( 
.A(n_4349),
.B(n_4353),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_SL g4793 ( 
.A(n_4144),
.B(n_2826),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4359),
.B(n_3360),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4150),
.B(n_3925),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4284),
.B(n_3940),
.Y(n_4796)
);

AND2x2_ASAP7_75t_L g4797 ( 
.A(n_4362),
.B(n_3360),
.Y(n_4797)
);

AND2x2_ASAP7_75t_L g4798 ( 
.A(n_4372),
.B(n_3360),
.Y(n_4798)
);

OAI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4177),
.A2(n_3428),
.B(n_3465),
.Y(n_4799)
);

INVx3_ASAP7_75t_L g4800 ( 
.A(n_4317),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4296),
.B(n_3951),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4296),
.B(n_3968),
.Y(n_4802)
);

INVx3_ASAP7_75t_L g4803 ( 
.A(n_4317),
.Y(n_4803)
);

AND2x2_ASAP7_75t_L g4804 ( 
.A(n_4386),
.B(n_3576),
.Y(n_4804)
);

INVxp67_ASAP7_75t_SL g4805 ( 
.A(n_4134),
.Y(n_4805)
);

HB1xp67_ASAP7_75t_L g4806 ( 
.A(n_4370),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_4344),
.B(n_3841),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4299),
.Y(n_4808)
);

INVx2_ASAP7_75t_L g4809 ( 
.A(n_4393),
.Y(n_4809)
);

INVx2_ASAP7_75t_L g4810 ( 
.A(n_4398),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4412),
.B(n_3999),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_SL g4812 ( 
.A(n_4220),
.B(n_2829),
.Y(n_4812)
);

INVx1_ASAP7_75t_SL g4813 ( 
.A(n_4485),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4402),
.B(n_3585),
.Y(n_4814)
);

INVx2_ASAP7_75t_SL g4815 ( 
.A(n_4170),
.Y(n_4815)
);

BUFx6f_ASAP7_75t_L g4816 ( 
.A(n_4175),
.Y(n_4816)
);

BUFx3_ASAP7_75t_L g4817 ( 
.A(n_4175),
.Y(n_4817)
);

INVx3_ASAP7_75t_L g4818 ( 
.A(n_4317),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4304),
.Y(n_4819)
);

AND2x2_ASAP7_75t_L g4820 ( 
.A(n_4417),
.B(n_3585),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4421),
.Y(n_4821)
);

OAI21x1_ASAP7_75t_L g4822 ( 
.A1(n_4229),
.A2(n_3237),
.B(n_3585),
.Y(n_4822)
);

BUFx6f_ASAP7_75t_L g4823 ( 
.A(n_4327),
.Y(n_4823)
);

AND2x2_ASAP7_75t_SL g4824 ( 
.A(n_4200),
.B(n_3923),
.Y(n_4824)
);

AND2x2_ASAP7_75t_L g4825 ( 
.A(n_4455),
.B(n_4461),
.Y(n_4825)
);

INVx2_ASAP7_75t_L g4826 ( 
.A(n_4466),
.Y(n_4826)
);

AND2x2_ASAP7_75t_L g4827 ( 
.A(n_4483),
.B(n_3588),
.Y(n_4827)
);

BUFx6f_ASAP7_75t_L g4828 ( 
.A(n_4327),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4308),
.Y(n_4829)
);

AND2x2_ASAP7_75t_SL g4830 ( 
.A(n_4223),
.B(n_3923),
.Y(n_4830)
);

AND2x2_ASAP7_75t_L g4831 ( 
.A(n_4313),
.B(n_3588),
.Y(n_4831)
);

AND2x2_ASAP7_75t_L g4832 ( 
.A(n_4316),
.B(n_3588),
.Y(n_4832)
);

AND2x2_ASAP7_75t_SL g4833 ( 
.A(n_4315),
.B(n_3928),
.Y(n_4833)
);

NOR2xp67_ASAP7_75t_L g4834 ( 
.A(n_4375),
.B(n_3881),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4318),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4321),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4324),
.B(n_3345),
.Y(n_4837)
);

OR2x2_ASAP7_75t_L g4838 ( 
.A(n_4432),
.B(n_3868),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4435),
.B(n_3818),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4325),
.Y(n_4840)
);

INVx2_ASAP7_75t_SL g4841 ( 
.A(n_4215),
.Y(n_4841)
);

INVx3_ASAP7_75t_L g4842 ( 
.A(n_4317),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4329),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4346),
.Y(n_4844)
);

AND2x4_ASAP7_75t_L g4845 ( 
.A(n_4350),
.B(n_3818),
.Y(n_4845)
);

HB1xp67_ASAP7_75t_L g4846 ( 
.A(n_4469),
.Y(n_4846)
);

NAND2x1p5_ASAP7_75t_L g4847 ( 
.A(n_4465),
.B(n_3748),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4360),
.Y(n_4848)
);

HB1xp67_ASAP7_75t_L g4849 ( 
.A(n_4452),
.Y(n_4849)
);

INVx4_ASAP7_75t_L g4850 ( 
.A(n_4487),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4368),
.Y(n_4851)
);

AND2x2_ASAP7_75t_L g4852 ( 
.A(n_4371),
.B(n_3345),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4392),
.Y(n_4853)
);

INVx4_ASAP7_75t_L g4854 ( 
.A(n_4317),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4415),
.Y(n_4855)
);

AND2x2_ASAP7_75t_SL g4856 ( 
.A(n_4178),
.B(n_3928),
.Y(n_4856)
);

AND2x6_ASAP7_75t_L g4857 ( 
.A(n_4430),
.B(n_3361),
.Y(n_4857)
);

INVx2_ASAP7_75t_L g4858 ( 
.A(n_4424),
.Y(n_4858)
);

INVxp33_ASAP7_75t_L g4859 ( 
.A(n_4383),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4100),
.B(n_3818),
.Y(n_4860)
);

INVx3_ASAP7_75t_L g4861 ( 
.A(n_4352),
.Y(n_4861)
);

AND2x2_ASAP7_75t_L g4862 ( 
.A(n_4436),
.B(n_2737),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4447),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4165),
.B(n_3876),
.Y(n_4864)
);

INVx3_ASAP7_75t_L g4865 ( 
.A(n_4352),
.Y(n_4865)
);

AND2x4_ASAP7_75t_L g4866 ( 
.A(n_4486),
.B(n_3876),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4211),
.B(n_2737),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4447),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_SL g4869 ( 
.A(n_4380),
.B(n_2829),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4134),
.Y(n_4870)
);

OR2x2_ASAP7_75t_L g4871 ( 
.A(n_4264),
.B(n_4188),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4395),
.B(n_3876),
.Y(n_4872)
);

AND2x2_ASAP7_75t_L g4873 ( 
.A(n_4164),
.B(n_2737),
.Y(n_4873)
);

HB1xp67_ASAP7_75t_L g4874 ( 
.A(n_4401),
.Y(n_4874)
);

NOR2xp33_ASAP7_75t_L g4875 ( 
.A(n_4162),
.B(n_2650),
.Y(n_4875)
);

NOR2xp33_ASAP7_75t_R g4876 ( 
.A(n_4102),
.B(n_2779),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_4169),
.B(n_2778),
.Y(n_4877)
);

INVxp33_ASAP7_75t_L g4878 ( 
.A(n_4440),
.Y(n_4878)
);

BUFx6f_ASAP7_75t_L g4879 ( 
.A(n_4476),
.Y(n_4879)
);

AND2x2_ASAP7_75t_L g4880 ( 
.A(n_4378),
.B(n_2778),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4179),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4127),
.B(n_4476),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4188),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4275),
.B(n_3887),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4288),
.B(n_3887),
.Y(n_4885)
);

INVx2_ASAP7_75t_L g4886 ( 
.A(n_4471),
.Y(n_4886)
);

HB1xp67_ASAP7_75t_L g4887 ( 
.A(n_4433),
.Y(n_4887)
);

AND2x2_ASAP7_75t_L g4888 ( 
.A(n_4127),
.B(n_2778),
.Y(n_4888)
);

BUFx3_ASAP7_75t_L g4889 ( 
.A(n_4230),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4212),
.Y(n_4890)
);

INVx2_ASAP7_75t_SL g4891 ( 
.A(n_4340),
.Y(n_4891)
);

INVxp67_ASAP7_75t_SL g4892 ( 
.A(n_4212),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4482),
.B(n_3361),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4292),
.B(n_3887),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4482),
.B(n_3362),
.Y(n_4895)
);

AND2x2_ASAP7_75t_L g4896 ( 
.A(n_4484),
.B(n_3362),
.Y(n_4896)
);

INVx3_ASAP7_75t_L g4897 ( 
.A(n_4352),
.Y(n_4897)
);

AND2x2_ASAP7_75t_L g4898 ( 
.A(n_4484),
.B(n_3908),
.Y(n_4898)
);

BUFx3_ASAP7_75t_L g4899 ( 
.A(n_4230),
.Y(n_4899)
);

AND2x4_ASAP7_75t_L g4900 ( 
.A(n_4341),
.B(n_3920),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4214),
.Y(n_4901)
);

NOR2xp33_ASAP7_75t_L g4902 ( 
.A(n_4418),
.B(n_2651),
.Y(n_4902)
);

HB1xp67_ASAP7_75t_L g4903 ( 
.A(n_4320),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4214),
.Y(n_4904)
);

INVx3_ASAP7_75t_L g4905 ( 
.A(n_4352),
.Y(n_4905)
);

HB1xp67_ASAP7_75t_L g4906 ( 
.A(n_4454),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4085),
.B(n_3908),
.Y(n_4907)
);

BUFx6f_ASAP7_75t_L g4908 ( 
.A(n_4216),
.Y(n_4908)
);

NOR2xp33_ASAP7_75t_L g4909 ( 
.A(n_4428),
.B(n_2653),
.Y(n_4909)
);

AND2x4_ASAP7_75t_L g4910 ( 
.A(n_4390),
.B(n_3920),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4197),
.B(n_3920),
.Y(n_4911)
);

HB1xp67_ASAP7_75t_L g4912 ( 
.A(n_4322),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4085),
.B(n_4009),
.Y(n_4913)
);

BUFx2_ASAP7_75t_L g4914 ( 
.A(n_4527),
.Y(n_4914)
);

BUFx6f_ASAP7_75t_L g4915 ( 
.A(n_4495),
.Y(n_4915)
);

NOR3xp33_ASAP7_75t_L g4916 ( 
.A(n_4638),
.B(n_4462),
.C(n_4467),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4835),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_SL g4918 ( 
.A(n_4768),
.B(n_4255),
.Y(n_4918)
);

AOI22xp33_ASAP7_75t_L g4919 ( 
.A1(n_4768),
.A2(n_4449),
.B1(n_4470),
.B2(n_4260),
.Y(n_4919)
);

INVx3_ASAP7_75t_L g4920 ( 
.A(n_4524),
.Y(n_4920)
);

INVx2_ASAP7_75t_L g4921 ( 
.A(n_4835),
.Y(n_4921)
);

BUFx2_ASAP7_75t_L g4922 ( 
.A(n_4527),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4507),
.B(n_4656),
.Y(n_4923)
);

AND2x2_ASAP7_75t_L g4924 ( 
.A(n_4561),
.B(n_4326),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4564),
.B(n_4405),
.Y(n_4925)
);

AOI21xp5_ASAP7_75t_L g4926 ( 
.A1(n_4502),
.A2(n_4161),
.B(n_4300),
.Y(n_4926)
);

AOI21xp5_ASAP7_75t_L g4927 ( 
.A1(n_4664),
.A2(n_4161),
.B(n_4456),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_SL g4928 ( 
.A(n_4583),
.B(n_4168),
.Y(n_4928)
);

AOI21xp5_ASAP7_75t_L g4929 ( 
.A1(n_4664),
.A2(n_3662),
.B(n_3656),
.Y(n_4929)
);

AOI21xp5_ASAP7_75t_L g4930 ( 
.A1(n_4500),
.A2(n_3662),
.B(n_3656),
.Y(n_4930)
);

INVx3_ASAP7_75t_L g4931 ( 
.A(n_4524),
.Y(n_4931)
);

BUFx6f_ASAP7_75t_L g4932 ( 
.A(n_4495),
.Y(n_4932)
);

HB1xp67_ASAP7_75t_L g4933 ( 
.A(n_4692),
.Y(n_4933)
);

A2O1A1Ixp33_ASAP7_75t_L g4934 ( 
.A1(n_4595),
.A2(n_4201),
.B(n_4264),
.C(n_4457),
.Y(n_4934)
);

AND2x6_ASAP7_75t_SL g4935 ( 
.A(n_4721),
.B(n_4429),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4766),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4561),
.B(n_4410),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4739),
.A2(n_3785),
.B(n_3781),
.Y(n_4938)
);

O2A1O1Ixp5_ASAP7_75t_L g4939 ( 
.A1(n_4697),
.A2(n_4763),
.B(n_4772),
.C(n_4733),
.Y(n_4939)
);

AOI33xp33_ASAP7_75t_L g4940 ( 
.A1(n_4530),
.A2(n_1274),
.A3(n_1176),
.B1(n_1198),
.B2(n_1102),
.B3(n_923),
.Y(n_4940)
);

NOR2xp33_ASAP7_75t_L g4941 ( 
.A(n_4878),
.B(n_4391),
.Y(n_4941)
);

AOI21xp5_ASAP7_75t_L g4942 ( 
.A1(n_4739),
.A2(n_4497),
.B(n_4551),
.Y(n_4942)
);

A2O1A1Ixp33_ASAP7_75t_L g4943 ( 
.A1(n_4727),
.A2(n_4416),
.B(n_4459),
.C(n_4434),
.Y(n_4943)
);

A2O1A1Ixp33_ASAP7_75t_L g4944 ( 
.A1(n_4506),
.A2(n_4338),
.B(n_4118),
.C(n_4479),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4844),
.Y(n_4945)
);

NOR2xp33_ASAP7_75t_L g4946 ( 
.A(n_4878),
.B(n_4336),
.Y(n_4946)
);

OR2x2_ASAP7_75t_L g4947 ( 
.A(n_4607),
.B(n_4142),
.Y(n_4947)
);

NAND2x1p5_ASAP7_75t_L g4948 ( 
.A(n_4613),
.B(n_4546),
.Y(n_4948)
);

A2O1A1Ixp33_ASAP7_75t_L g4949 ( 
.A1(n_4909),
.A2(n_4480),
.B(n_4348),
.C(n_4333),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4508),
.B(n_4422),
.Y(n_4950)
);

HB1xp67_ASAP7_75t_L g4951 ( 
.A(n_4685),
.Y(n_4951)
);

AOI21xp5_ASAP7_75t_L g4952 ( 
.A1(n_4497),
.A2(n_3785),
.B(n_3781),
.Y(n_4952)
);

BUFx8_ASAP7_75t_L g4953 ( 
.A(n_4841),
.Y(n_4953)
);

AOI21x1_ASAP7_75t_L g4954 ( 
.A1(n_4496),
.A2(n_3805),
.B(n_3801),
.Y(n_4954)
);

OAI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4799),
.A2(n_3413),
.B(n_3400),
.Y(n_4955)
);

OAI22xp5_ASAP7_75t_L g4956 ( 
.A1(n_4536),
.A2(n_3722),
.B1(n_3892),
.B2(n_3890),
.Y(n_4956)
);

AND2x4_ASAP7_75t_L g4957 ( 
.A(n_4539),
.B(n_3922),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_SL g4958 ( 
.A(n_4774),
.B(n_4397),
.Y(n_4958)
);

AOI21x1_ASAP7_75t_L g4959 ( 
.A1(n_4496),
.A2(n_4867),
.B(n_4520),
.Y(n_4959)
);

AOI21xp5_ASAP7_75t_L g4960 ( 
.A1(n_4691),
.A2(n_3959),
.B(n_3936),
.Y(n_4960)
);

BUFx12f_ASAP7_75t_L g4961 ( 
.A(n_4760),
.Y(n_4961)
);

INVx4_ASAP7_75t_L g4962 ( 
.A(n_4524),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4691),
.A2(n_3991),
.B(n_3996),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4708),
.A2(n_3996),
.B(n_4105),
.Y(n_4964)
);

O2A1O1Ixp33_ASAP7_75t_L g4965 ( 
.A1(n_4700),
.A2(n_1267),
.B(n_1198),
.C(n_1176),
.Y(n_4965)
);

OAI21xp5_ASAP7_75t_L g4966 ( 
.A1(n_4676),
.A2(n_4414),
.B(n_3559),
.Y(n_4966)
);

AOI22xp5_ASAP7_75t_L g4967 ( 
.A1(n_4791),
.A2(n_2875),
.B1(n_2907),
.B2(n_2781),
.Y(n_4967)
);

INVxp67_ASAP7_75t_L g4968 ( 
.A(n_4488),
.Y(n_4968)
);

INVx4_ASAP7_75t_L g4969 ( 
.A(n_4524),
.Y(n_4969)
);

NOR2xp33_ASAP7_75t_L g4970 ( 
.A(n_4859),
.B(n_2653),
.Y(n_4970)
);

OAI22xp5_ASAP7_75t_L g4971 ( 
.A1(n_4859),
.A2(n_3850),
.B1(n_3709),
.B2(n_2707),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4844),
.Y(n_4972)
);

AOI21xp5_ASAP7_75t_L g4973 ( 
.A1(n_4708),
.A2(n_4116),
.B(n_4105),
.Y(n_4973)
);

AOI21xp5_ASAP7_75t_L g4974 ( 
.A1(n_4713),
.A2(n_4122),
.B(n_4116),
.Y(n_4974)
);

A2O1A1Ixp33_ASAP7_75t_L g4975 ( 
.A1(n_4744),
.A2(n_3578),
.B(n_3575),
.C(n_3558),
.Y(n_4975)
);

AOI21xp5_ASAP7_75t_L g4976 ( 
.A1(n_4713),
.A2(n_4575),
.B(n_4613),
.Y(n_4976)
);

AOI21xp5_ASAP7_75t_L g4977 ( 
.A1(n_4613),
.A2(n_4122),
.B(n_3607),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4537),
.B(n_4216),
.Y(n_4978)
);

AO21x1_ASAP7_75t_L g4979 ( 
.A1(n_4761),
.A2(n_4473),
.B(n_4471),
.Y(n_4979)
);

INVx2_ASAP7_75t_L g4980 ( 
.A(n_4848),
.Y(n_4980)
);

AOI21xp5_ASAP7_75t_L g4981 ( 
.A1(n_4786),
.A2(n_3607),
.B(n_3359),
.Y(n_4981)
);

OAI21xp5_ASAP7_75t_L g4982 ( 
.A1(n_4519),
.A2(n_3606),
.B(n_3864),
.Y(n_4982)
);

AOI21xp5_ASAP7_75t_L g4983 ( 
.A1(n_4786),
.A2(n_3607),
.B(n_3336),
.Y(n_4983)
);

OAI22xp5_ASAP7_75t_L g4984 ( 
.A1(n_4863),
.A2(n_4261),
.B1(n_4262),
.B2(n_4259),
.Y(n_4984)
);

OAI21xp5_ASAP7_75t_L g4985 ( 
.A1(n_4745),
.A2(n_3606),
.B(n_3895),
.Y(n_4985)
);

NOR2xp67_ASAP7_75t_L g4986 ( 
.A(n_4891),
.B(n_2837),
.Y(n_4986)
);

CKINVDCx10_ASAP7_75t_R g4987 ( 
.A(n_4526),
.Y(n_4987)
);

AND2x2_ASAP7_75t_L g4988 ( 
.A(n_4517),
.B(n_3922),
.Y(n_4988)
);

O2A1O1Ixp33_ASAP7_75t_SL g4989 ( 
.A1(n_4812),
.A2(n_985),
.B(n_1071),
.C(n_925),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4766),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4537),
.B(n_4259),
.Y(n_4991)
);

AOI21x1_ASAP7_75t_L g4992 ( 
.A1(n_4867),
.A2(n_3085),
.B(n_3910),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4618),
.B(n_4261),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4863),
.A2(n_3246),
.B(n_3194),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4787),
.Y(n_4995)
);

NOR2xp33_ASAP7_75t_L g4996 ( 
.A(n_4698),
.B(n_2661),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4517),
.B(n_3922),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4801),
.B(n_4262),
.Y(n_4998)
);

CKINVDCx5p33_ASAP7_75t_R g4999 ( 
.A(n_4526),
.Y(n_4999)
);

AOI21xp5_ASAP7_75t_L g5000 ( 
.A1(n_4868),
.A2(n_3246),
.B(n_3194),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4553),
.B(n_3924),
.Y(n_5001)
);

INVx1_ASAP7_75t_SL g5002 ( 
.A(n_4802),
.Y(n_5002)
);

A2O1A1Ixp33_ASAP7_75t_L g5003 ( 
.A1(n_4902),
.A2(n_3246),
.B(n_3312),
.C(n_3194),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4868),
.A2(n_3312),
.B(n_3246),
.Y(n_5004)
);

OAI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_4745),
.A2(n_4263),
.B1(n_4268),
.B2(n_4267),
.Y(n_5005)
);

OAI21xp33_ASAP7_75t_L g5006 ( 
.A1(n_4503),
.A2(n_4301),
.B(n_2842),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4788),
.B(n_4263),
.Y(n_5007)
);

AOI21xp5_ASAP7_75t_L g5008 ( 
.A1(n_4511),
.A2(n_3312),
.B(n_3246),
.Y(n_5008)
);

BUFx6f_ASAP7_75t_L g5009 ( 
.A(n_4528),
.Y(n_5009)
);

NAND2x1_ASAP7_75t_L g5010 ( 
.A(n_4491),
.B(n_3848),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4848),
.Y(n_5011)
);

AOI22xp5_ASAP7_75t_L g5012 ( 
.A1(n_4869),
.A2(n_4549),
.B1(n_4663),
.B2(n_4875),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4851),
.Y(n_5013)
);

AOI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_4511),
.A2(n_3312),
.B(n_3748),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_SL g5015 ( 
.A(n_4795),
.B(n_2837),
.Y(n_5015)
);

AOI21xp5_ASAP7_75t_L g5016 ( 
.A1(n_4534),
.A2(n_3312),
.B(n_3748),
.Y(n_5016)
);

NOR2xp33_ASAP7_75t_L g5017 ( 
.A(n_4906),
.B(n_2661),
.Y(n_5017)
);

AOI21xp5_ASAP7_75t_L g5018 ( 
.A1(n_4534),
.A2(n_3765),
.B(n_3748),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4552),
.B(n_4267),
.Y(n_5019)
);

AOI21xp5_ASAP7_75t_L g5020 ( 
.A1(n_4560),
.A2(n_3767),
.B(n_3765),
.Y(n_5020)
);

AND2x2_ASAP7_75t_L g5021 ( 
.A(n_4553),
.B(n_3924),
.Y(n_5021)
);

INVx4_ASAP7_75t_L g5022 ( 
.A(n_4524),
.Y(n_5022)
);

INVx3_ASAP7_75t_L g5023 ( 
.A(n_4816),
.Y(n_5023)
);

NOR2xp33_ASAP7_75t_L g5024 ( 
.A(n_4730),
.B(n_4717),
.Y(n_5024)
);

OAI21x1_ASAP7_75t_L g5025 ( 
.A1(n_4619),
.A2(n_3889),
.B(n_3884),
.Y(n_5025)
);

OAI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_4762),
.A2(n_3431),
.B(n_3418),
.Y(n_5026)
);

OAI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4651),
.A2(n_3432),
.B(n_3471),
.Y(n_5027)
);

OAI21xp5_ASAP7_75t_L g5028 ( 
.A1(n_4873),
.A2(n_3509),
.B(n_4473),
.Y(n_5028)
);

AOI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4560),
.A2(n_3767),
.B(n_3765),
.Y(n_5029)
);

HB1xp67_ASAP7_75t_L g5030 ( 
.A(n_4903),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4571),
.B(n_4268),
.Y(n_5031)
);

OAI22xp5_ASAP7_75t_L g5032 ( 
.A1(n_4571),
.A2(n_4276),
.B1(n_4287),
.B2(n_4270),
.Y(n_5032)
);

HB1xp67_ASAP7_75t_L g5033 ( 
.A(n_4546),
.Y(n_5033)
);

OAI22xp5_ASAP7_75t_L g5034 ( 
.A1(n_4585),
.A2(n_4276),
.B1(n_4287),
.B2(n_4270),
.Y(n_5034)
);

AOI21xp5_ASAP7_75t_L g5035 ( 
.A1(n_4585),
.A2(n_3767),
.B(n_3765),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_SL g5036 ( 
.A(n_4636),
.B(n_2842),
.Y(n_5036)
);

OAI21xp33_ASAP7_75t_L g5037 ( 
.A1(n_4675),
.A2(n_985),
.B(n_925),
.Y(n_5037)
);

AOI22xp5_ASAP7_75t_L g5038 ( 
.A1(n_4789),
.A2(n_2907),
.B1(n_2875),
.B2(n_2781),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4605),
.B(n_4297),
.Y(n_5039)
);

OAI22xp5_ASAP7_75t_L g5040 ( 
.A1(n_4695),
.A2(n_2705),
.B1(n_2708),
.B2(n_2707),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4559),
.B(n_3924),
.Y(n_5041)
);

AO21x1_ASAP7_75t_L g5042 ( 
.A1(n_4731),
.A2(n_923),
.B(n_922),
.Y(n_5042)
);

INVxp67_ASAP7_75t_SL g5043 ( 
.A(n_4490),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4559),
.B(n_3927),
.Y(n_5044)
);

AOI21xp5_ASAP7_75t_L g5045 ( 
.A1(n_4605),
.A2(n_3937),
.B(n_3767),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4525),
.B(n_3927),
.Y(n_5046)
);

O2A1O1Ixp5_ASAP7_75t_L g5047 ( 
.A1(n_4491),
.A2(n_3889),
.B(n_3915),
.C(n_3884),
.Y(n_5047)
);

NOR2xp33_ASAP7_75t_L g5048 ( 
.A(n_4872),
.B(n_2705),
.Y(n_5048)
);

AND2x4_ASAP7_75t_L g5049 ( 
.A(n_4539),
.B(n_3927),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_4851),
.Y(n_5050)
);

AOI21xp5_ASAP7_75t_L g5051 ( 
.A1(n_4805),
.A2(n_3967),
.B(n_3937),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4525),
.B(n_3932),
.Y(n_5052)
);

BUFx3_ASAP7_75t_L g5053 ( 
.A(n_4528),
.Y(n_5053)
);

AOI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4892),
.A2(n_3967),
.B(n_3937),
.Y(n_5054)
);

NOR2xp33_ASAP7_75t_L g5055 ( 
.A(n_4602),
.B(n_2708),
.Y(n_5055)
);

OAI22xp5_ASAP7_75t_L g5056 ( 
.A1(n_4695),
.A2(n_2714),
.B1(n_2783),
.B2(n_2782),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_4839),
.B(n_4297),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4787),
.Y(n_5058)
);

AOI22xp5_ASAP7_75t_L g5059 ( 
.A1(n_4680),
.A2(n_2782),
.B1(n_2783),
.B2(n_2688),
.Y(n_5059)
);

AOI21xp5_ASAP7_75t_L g5060 ( 
.A1(n_4765),
.A2(n_3967),
.B(n_3937),
.Y(n_5060)
);

A2O1A1Ixp33_ASAP7_75t_L g5061 ( 
.A1(n_4574),
.A2(n_925),
.B(n_1071),
.C(n_985),
.Y(n_5061)
);

BUFx3_ASAP7_75t_L g5062 ( 
.A(n_4518),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4881),
.B(n_4448),
.Y(n_5063)
);

AND2x2_ASAP7_75t_L g5064 ( 
.A(n_4532),
.B(n_3932),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4790),
.Y(n_5065)
);

INVx3_ASAP7_75t_L g5066 ( 
.A(n_4816),
.Y(n_5066)
);

OAI21xp5_ASAP7_75t_L g5067 ( 
.A1(n_4873),
.A2(n_3941),
.B(n_3915),
.Y(n_5067)
);

AND2x4_ASAP7_75t_L g5068 ( 
.A(n_4539),
.B(n_3932),
.Y(n_5068)
);

AOI21x1_ASAP7_75t_L g5069 ( 
.A1(n_4877),
.A2(n_3085),
.B(n_4448),
.Y(n_5069)
);

NOR2x1_ASAP7_75t_L g5070 ( 
.A(n_4796),
.B(n_4793),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_4633),
.B(n_4541),
.Y(n_5071)
);

AOI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4765),
.A2(n_4516),
.B(n_3967),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_SL g5073 ( 
.A(n_4833),
.B(n_4775),
.Y(n_5073)
);

NOR2xp33_ASAP7_75t_L g5074 ( 
.A(n_4657),
.B(n_2714),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_SL g5075 ( 
.A(n_4833),
.B(n_3896),
.Y(n_5075)
);

O2A1O1Ixp5_ASAP7_75t_L g5076 ( 
.A1(n_4491),
.A2(n_3947),
.B(n_3950),
.C(n_3941),
.Y(n_5076)
);

AO21x1_ASAP7_75t_L g5077 ( 
.A1(n_4732),
.A2(n_929),
.B(n_924),
.Y(n_5077)
);

INVx2_ASAP7_75t_L g5078 ( 
.A(n_4858),
.Y(n_5078)
);

O2A1O1Ixp33_ASAP7_75t_L g5079 ( 
.A1(n_4811),
.A2(n_1095),
.B(n_1104),
.C(n_1071),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4541),
.B(n_3946),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4545),
.B(n_3946),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4545),
.B(n_3946),
.Y(n_5082)
);

OAI22xp5_ASAP7_75t_L g5083 ( 
.A1(n_4608),
.A2(n_4272),
.B1(n_2982),
.B2(n_2987),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4790),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4808),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4547),
.B(n_4009),
.Y(n_5086)
);

AOI21x1_ASAP7_75t_L g5087 ( 
.A1(n_4877),
.A2(n_3085),
.B(n_3847),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4547),
.B(n_4013),
.Y(n_5088)
);

O2A1O1Ixp33_ASAP7_75t_L g5089 ( 
.A1(n_4912),
.A2(n_1104),
.B(n_1146),
.C(n_1095),
.Y(n_5089)
);

AND2x2_ASAP7_75t_L g5090 ( 
.A(n_4532),
.B(n_4648),
.Y(n_5090)
);

OAI21xp33_ASAP7_75t_L g5091 ( 
.A1(n_4705),
.A2(n_1104),
.B(n_1095),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4765),
.A2(n_3741),
.B(n_3372),
.Y(n_5092)
);

OAI21xp33_ASAP7_75t_L g5093 ( 
.A1(n_4726),
.A2(n_4702),
.B(n_4586),
.Y(n_5093)
);

AOI21xp5_ASAP7_75t_L g5094 ( 
.A1(n_4765),
.A2(n_3741),
.B(n_3372),
.Y(n_5094)
);

AOI21xp5_ASAP7_75t_L g5095 ( 
.A1(n_4516),
.A2(n_3372),
.B(n_3338),
.Y(n_5095)
);

O2A1O1Ixp33_ASAP7_75t_L g5096 ( 
.A1(n_4860),
.A2(n_1146),
.B(n_929),
.C(n_936),
.Y(n_5096)
);

AOI21xp5_ASAP7_75t_L g5097 ( 
.A1(n_4662),
.A2(n_4621),
.B(n_4620),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_4858),
.Y(n_5098)
);

AND2x4_ASAP7_75t_L g5099 ( 
.A(n_4489),
.B(n_4251),
.Y(n_5099)
);

AOI21xp5_ASAP7_75t_L g5100 ( 
.A1(n_4606),
.A2(n_3372),
.B(n_3338),
.Y(n_5100)
);

INVxp67_ASAP7_75t_L g5101 ( 
.A(n_4644),
.Y(n_5101)
);

AND2x2_ASAP7_75t_SL g5102 ( 
.A(n_4617),
.B(n_4113),
.Y(n_5102)
);

BUFx4f_ASAP7_75t_L g5103 ( 
.A(n_4562),
.Y(n_5103)
);

O2A1O1Ixp33_ASAP7_75t_L g5104 ( 
.A1(n_4849),
.A2(n_1146),
.B(n_936),
.C(n_937),
.Y(n_5104)
);

AOI21xp5_ASAP7_75t_L g5105 ( 
.A1(n_4606),
.A2(n_3338),
.B(n_3731),
.Y(n_5105)
);

AOI21xp5_ASAP7_75t_L g5106 ( 
.A1(n_4620),
.A2(n_3338),
.B(n_3731),
.Y(n_5106)
);

AOI21xp5_ASAP7_75t_L g5107 ( 
.A1(n_4621),
.A2(n_3764),
.B(n_3761),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_L g5108 ( 
.A(n_4540),
.B(n_4013),
.Y(n_5108)
);

A2O1A1Ixp33_ASAP7_75t_L g5109 ( 
.A1(n_4550),
.A2(n_937),
.B(n_939),
.C(n_924),
.Y(n_5109)
);

BUFx3_ASAP7_75t_L g5110 ( 
.A(n_4518),
.Y(n_5110)
);

OAI321xp33_ASAP7_75t_L g5111 ( 
.A1(n_4911),
.A2(n_943),
.A3(n_944),
.B1(n_949),
.B2(n_945),
.C(n_939),
.Y(n_5111)
);

O2A1O1Ixp33_ASAP7_75t_L g5112 ( 
.A1(n_4769),
.A2(n_944),
.B(n_945),
.C(n_943),
.Y(n_5112)
);

NOR2xp33_ASAP7_75t_L g5113 ( 
.A(n_4716),
.B(n_2217),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_4540),
.B(n_4022),
.Y(n_5114)
);

AOI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_4629),
.A2(n_3764),
.B(n_3761),
.Y(n_5115)
);

A2O1A1Ixp33_ASAP7_75t_L g5116 ( 
.A1(n_4900),
.A2(n_955),
.B(n_957),
.C(n_949),
.Y(n_5116)
);

NAND2xp5_ASAP7_75t_L g5117 ( 
.A(n_4908),
.B(n_4022),
.Y(n_5117)
);

NAND2xp5_ASAP7_75t_L g5118 ( 
.A(n_4908),
.B(n_4031),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_4908),
.B(n_2688),
.Y(n_5119)
);

AND2x6_ASAP7_75t_SL g5120 ( 
.A(n_4758),
.B(n_4760),
.Y(n_5120)
);

AOI21xp5_ASAP7_75t_L g5121 ( 
.A1(n_4629),
.A2(n_3819),
.B(n_3794),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_4908),
.B(n_2369),
.Y(n_5122)
);

AOI21x1_ASAP7_75t_L g5123 ( 
.A1(n_4880),
.A2(n_3847),
.B(n_3595),
.Y(n_5123)
);

AOI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_4646),
.A2(n_3866),
.B(n_3819),
.Y(n_5124)
);

AOI22xp5_ASAP7_75t_L g5125 ( 
.A1(n_4764),
.A2(n_2691),
.B1(n_2785),
.B2(n_2982),
.Y(n_5125)
);

OAI21xp5_ASAP7_75t_L g5126 ( 
.A1(n_4880),
.A2(n_3950),
.B(n_3947),
.Y(n_5126)
);

NOR2x1_ASAP7_75t_SL g5127 ( 
.A(n_4693),
.B(n_3969),
.Y(n_5127)
);

CKINVDCx10_ASAP7_75t_R g5128 ( 
.A(n_4760),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_SL g5129 ( 
.A(n_4900),
.B(n_3896),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4493),
.Y(n_5130)
);

AOI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_4646),
.A2(n_3866),
.B(n_3794),
.Y(n_5131)
);

INVx3_ASAP7_75t_L g5132 ( 
.A(n_4816),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_4908),
.B(n_2369),
.Y(n_5133)
);

NOR2x1_ASAP7_75t_L g5134 ( 
.A(n_4834),
.B(n_3955),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_SL g5135 ( 
.A(n_4900),
.B(n_3897),
.Y(n_5135)
);

NOR2xp33_ASAP7_75t_L g5136 ( 
.A(n_4813),
.B(n_2691),
.Y(n_5136)
);

AND2x2_ASAP7_75t_SL g5137 ( 
.A(n_4617),
.B(n_3955),
.Y(n_5137)
);

INVx11_ASAP7_75t_L g5138 ( 
.A(n_4857),
.Y(n_5138)
);

AOI21xp5_ASAP7_75t_L g5139 ( 
.A1(n_4647),
.A2(n_3880),
.B(n_3875),
.Y(n_5139)
);

AOI21xp5_ASAP7_75t_L g5140 ( 
.A1(n_4647),
.A2(n_3880),
.B(n_3875),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4808),
.Y(n_5141)
);

AOI21xp5_ASAP7_75t_L g5142 ( 
.A1(n_4678),
.A2(n_3964),
.B(n_3953),
.Y(n_5142)
);

NOR2xp33_ASAP7_75t_L g5143 ( 
.A(n_4577),
.B(n_2691),
.Y(n_5143)
);

AND2x4_ASAP7_75t_L g5144 ( 
.A(n_4489),
.B(n_3832),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_4686),
.B(n_3897),
.Y(n_5145)
);

BUFx6f_ASAP7_75t_L g5146 ( 
.A(n_4562),
.Y(n_5146)
);

O2A1O1Ixp33_ASAP7_75t_L g5147 ( 
.A1(n_4846),
.A2(n_957),
.B(n_960),
.C(n_955),
.Y(n_5147)
);

NAND2x1p5_ASAP7_75t_L g5148 ( 
.A(n_4515),
.B(n_4063),
.Y(n_5148)
);

BUFx6f_ASAP7_75t_L g5149 ( 
.A(n_4562),
.Y(n_5149)
);

OAI21xp5_ASAP7_75t_L g5150 ( 
.A1(n_4660),
.A2(n_3964),
.B(n_3953),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4836),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_4836),
.Y(n_5152)
);

NOR2xp33_ASAP7_75t_L g5153 ( 
.A(n_4582),
.B(n_2785),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_SL g5154 ( 
.A(n_4736),
.B(n_2785),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_4840),
.Y(n_5155)
);

AOI21xp33_ASAP7_75t_L g5156 ( 
.A1(n_4838),
.A2(n_3435),
.B(n_3382),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4568),
.B(n_4901),
.Y(n_5157)
);

AOI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4678),
.A2(n_3998),
.B(n_3971),
.Y(n_5158)
);

BUFx6f_ASAP7_75t_L g5159 ( 
.A(n_4562),
.Y(n_5159)
);

INVx2_ASAP7_75t_L g5160 ( 
.A(n_4493),
.Y(n_5160)
);

AO21x1_ASAP7_75t_L g5161 ( 
.A1(n_4732),
.A2(n_962),
.B(n_960),
.Y(n_5161)
);

AOI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_4707),
.A2(n_3998),
.B(n_3971),
.Y(n_5162)
);

O2A1O1Ixp33_ASAP7_75t_L g5163 ( 
.A1(n_4728),
.A2(n_966),
.B(n_973),
.C(n_962),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4840),
.Y(n_5164)
);

AOI21xp5_ASAP7_75t_L g5165 ( 
.A1(n_4707),
.A2(n_4012),
.B(n_4008),
.Y(n_5165)
);

AOI21xp5_ASAP7_75t_L g5166 ( 
.A1(n_4589),
.A2(n_4012),
.B(n_4008),
.Y(n_5166)
);

AOI21xp5_ASAP7_75t_L g5167 ( 
.A1(n_4522),
.A2(n_4543),
.B(n_4531),
.Y(n_5167)
);

CKINVDCx5p33_ASAP7_75t_R g5168 ( 
.A(n_4645),
.Y(n_5168)
);

AOI21xp5_ASAP7_75t_L g5169 ( 
.A1(n_4522),
.A2(n_3979),
.B(n_3976),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_4531),
.A2(n_3979),
.B(n_3976),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_4686),
.B(n_966),
.Y(n_5171)
);

OAI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_4568),
.A2(n_4035),
.B(n_3854),
.Y(n_5172)
);

A2O1A1Ixp33_ASAP7_75t_L g5173 ( 
.A1(n_4856),
.A2(n_978),
.B(n_981),
.C(n_973),
.Y(n_5173)
);

NAND2x1p5_ASAP7_75t_L g5174 ( 
.A(n_4515),
.B(n_4565),
.Y(n_5174)
);

NOR2xp33_ASAP7_75t_L g5175 ( 
.A(n_4759),
.B(n_2983),
.Y(n_5175)
);

NOR2xp33_ASAP7_75t_L g5176 ( 
.A(n_4780),
.B(n_2983),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4843),
.Y(n_5177)
);

CKINVDCx20_ASAP7_75t_R g5178 ( 
.A(n_4645),
.Y(n_5178)
);

OAI21xp5_ASAP7_75t_L g5179 ( 
.A1(n_4838),
.A2(n_4035),
.B(n_3854),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_4870),
.B(n_4901),
.Y(n_5180)
);

NOR2xp33_ASAP7_75t_L g5181 ( 
.A(n_4556),
.B(n_2987),
.Y(n_5181)
);

AND2x2_ASAP7_75t_L g5182 ( 
.A(n_4783),
.B(n_978),
.Y(n_5182)
);

NAND2xp33_ASAP7_75t_L g5183 ( 
.A(n_4876),
.B(n_2988),
.Y(n_5183)
);

AOI21xp5_ASAP7_75t_L g5184 ( 
.A1(n_4543),
.A2(n_3367),
.B(n_3366),
.Y(n_5184)
);

NOR2xp33_ASAP7_75t_L g5185 ( 
.A(n_4569),
.B(n_2988),
.Y(n_5185)
);

NAND2x1p5_ASAP7_75t_L g5186 ( 
.A(n_4515),
.B(n_4015),
.Y(n_5186)
);

AND2x4_ASAP7_75t_L g5187 ( 
.A(n_4489),
.B(n_3832),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_4870),
.B(n_2369),
.Y(n_5188)
);

CKINVDCx20_ASAP7_75t_R g5189 ( 
.A(n_4757),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_4783),
.B(n_981),
.Y(n_5190)
);

AOI21xp5_ASAP7_75t_L g5191 ( 
.A1(n_4566),
.A2(n_3367),
.B(n_3366),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_4883),
.B(n_2386),
.Y(n_5192)
);

NAND2x1p5_ASAP7_75t_L g5193 ( 
.A(n_4565),
.B(n_3969),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_SL g5194 ( 
.A(n_4736),
.B(n_4420),
.Y(n_5194)
);

O2A1O1Ixp5_ASAP7_75t_L g5195 ( 
.A1(n_4565),
.A2(n_3456),
.B(n_3496),
.C(n_3491),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_4883),
.B(n_2386),
.Y(n_5196)
);

INVxp67_ASAP7_75t_L g5197 ( 
.A(n_4755),
.Y(n_5197)
);

NOR2xp33_ASAP7_75t_L g5198 ( 
.A(n_4588),
.B(n_4616),
.Y(n_5198)
);

OAI22xp33_ASAP7_75t_L g5199 ( 
.A1(n_4841),
.A2(n_2999),
.B1(n_3012),
.B2(n_2989),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_4792),
.B(n_984),
.Y(n_5200)
);

O2A1O1Ixp33_ASAP7_75t_L g5201 ( 
.A1(n_4874),
.A2(n_989),
.B(n_991),
.C(n_984),
.Y(n_5201)
);

NOR2xp67_ASAP7_75t_L g5202 ( 
.A(n_4891),
.B(n_2989),
.Y(n_5202)
);

AOI21xp5_ASAP7_75t_L g5203 ( 
.A1(n_4566),
.A2(n_3373),
.B(n_3370),
.Y(n_5203)
);

OAI21xp5_ASAP7_75t_L g5204 ( 
.A1(n_4505),
.A2(n_4045),
.B(n_4043),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_4567),
.A2(n_3373),
.B(n_3370),
.Y(n_5205)
);

AOI21xp5_ASAP7_75t_L g5206 ( 
.A1(n_4567),
.A2(n_3376),
.B(n_3172),
.Y(n_5206)
);

AOI21xp5_ASAP7_75t_L g5207 ( 
.A1(n_4578),
.A2(n_3376),
.B(n_3172),
.Y(n_5207)
);

BUFx4f_ASAP7_75t_L g5208 ( 
.A(n_4562),
.Y(n_5208)
);

AOI21x1_ASAP7_75t_L g5209 ( 
.A1(n_4888),
.A2(n_4043),
.B(n_4045),
.Y(n_5209)
);

AOI22xp33_ASAP7_75t_L g5210 ( 
.A1(n_4856),
.A2(n_4830),
.B1(n_4824),
.B2(n_4764),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_4890),
.B(n_4904),
.Y(n_5211)
);

HB1xp67_ASAP7_75t_L g5212 ( 
.A(n_4767),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_4890),
.B(n_2386),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_4533),
.B(n_3860),
.Y(n_5214)
);

NAND2xp5_ASAP7_75t_L g5215 ( 
.A(n_4904),
.B(n_2405),
.Y(n_5215)
);

OAI22xp5_ASAP7_75t_L g5216 ( 
.A1(n_4666),
.A2(n_3012),
.B1(n_3019),
.B2(n_2999),
.Y(n_5216)
);

AOI21xp5_ASAP7_75t_L g5217 ( 
.A1(n_4578),
.A2(n_4594),
.B(n_4579),
.Y(n_5217)
);

AOI21xp5_ASAP7_75t_L g5218 ( 
.A1(n_4579),
.A2(n_3172),
.B(n_3113),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_4843),
.Y(n_5219)
);

AOI21xp5_ASAP7_75t_L g5220 ( 
.A1(n_4594),
.A2(n_3172),
.B(n_3113),
.Y(n_5220)
);

AO32x2_ASAP7_75t_L g5221 ( 
.A1(n_4494),
.A2(n_4854),
.A3(n_4815),
.B1(n_4504),
.B2(n_4650),
.Y(n_5221)
);

NOR2xp67_ASAP7_75t_L g5222 ( 
.A(n_4850),
.B(n_3019),
.Y(n_5222)
);

INVx2_ASAP7_75t_L g5223 ( 
.A(n_4498),
.Y(n_5223)
);

OAI22xp5_ASAP7_75t_L g5224 ( 
.A1(n_4871),
.A2(n_3199),
.B1(n_3236),
.B2(n_3113),
.Y(n_5224)
);

BUFx6f_ASAP7_75t_L g5225 ( 
.A(n_4572),
.Y(n_5225)
);

AOI21xp5_ASAP7_75t_L g5226 ( 
.A1(n_4597),
.A2(n_3199),
.B(n_3113),
.Y(n_5226)
);

BUFx8_ASAP7_75t_L g5227 ( 
.A(n_4889),
.Y(n_5227)
);

BUFx3_ASAP7_75t_L g5228 ( 
.A(n_4684),
.Y(n_5228)
);

O2A1O1Ixp33_ASAP7_75t_L g5229 ( 
.A1(n_4887),
.A2(n_991),
.B(n_992),
.C(n_989),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_4641),
.B(n_2405),
.Y(n_5230)
);

NOR2xp33_ASAP7_75t_R g5231 ( 
.A(n_4889),
.B(n_3024),
.Y(n_5231)
);

NOR2xp33_ASAP7_75t_L g5232 ( 
.A(n_4690),
.B(n_3024),
.Y(n_5232)
);

INVx2_ASAP7_75t_SL g5233 ( 
.A(n_4684),
.Y(n_5233)
);

CKINVDCx8_ASAP7_75t_R g5234 ( 
.A(n_4682),
.Y(n_5234)
);

AOI22xp33_ASAP7_75t_L g5235 ( 
.A1(n_4824),
.A2(n_4420),
.B1(n_902),
.B2(n_976),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_4498),
.Y(n_5236)
);

NAND2xp5_ASAP7_75t_L g5237 ( 
.A(n_4898),
.B(n_2405),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_4523),
.Y(n_5238)
);

NOR2xp33_ASAP7_75t_L g5239 ( 
.A(n_4690),
.B(n_1335),
.Y(n_5239)
);

CKINVDCx14_ASAP7_75t_R g5240 ( 
.A(n_4899),
.Y(n_5240)
);

AOI21xp5_ASAP7_75t_L g5241 ( 
.A1(n_4597),
.A2(n_3236),
.B(n_3199),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_L g5242 ( 
.A(n_4898),
.B(n_2270),
.Y(n_5242)
);

BUFx6f_ASAP7_75t_L g5243 ( 
.A(n_4572),
.Y(n_5243)
);

AOI21xp5_ASAP7_75t_L g5244 ( 
.A1(n_4610),
.A2(n_3236),
.B(n_3199),
.Y(n_5244)
);

AOI21xp5_ASAP7_75t_L g5245 ( 
.A1(n_4610),
.A2(n_3236),
.B(n_3667),
.Y(n_5245)
);

AO32x1_ASAP7_75t_L g5246 ( 
.A1(n_4494),
.A2(n_1010),
.A3(n_1012),
.B1(n_1002),
.B2(n_992),
.Y(n_5246)
);

AOI21xp5_ASAP7_75t_L g5247 ( 
.A1(n_4639),
.A2(n_3728),
.B(n_3853),
.Y(n_5247)
);

A2O1A1Ixp33_ASAP7_75t_L g5248 ( 
.A1(n_4830),
.A2(n_1010),
.B(n_1012),
.C(n_1002),
.Y(n_5248)
);

BUFx2_ASAP7_75t_SL g5249 ( 
.A(n_4752),
.Y(n_5249)
);

NOR2xp33_ASAP7_75t_L g5250 ( 
.A(n_4690),
.B(n_4806),
.Y(n_5250)
);

AOI21xp5_ASAP7_75t_L g5251 ( 
.A1(n_4639),
.A2(n_3728),
.B(n_3853),
.Y(n_5251)
);

AOI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_4654),
.A2(n_3859),
.B(n_3598),
.Y(n_5252)
);

NOR2xp67_ASAP7_75t_L g5253 ( 
.A(n_4850),
.B(n_3614),
.Y(n_5253)
);

OAI22xp5_ASAP7_75t_L g5254 ( 
.A1(n_4666),
.A2(n_3593),
.B1(n_3623),
.B2(n_3614),
.Y(n_5254)
);

AOI22x1_ASAP7_75t_L g5255 ( 
.A1(n_4847),
.A2(n_3675),
.B1(n_3679),
.B2(n_3623),
.Y(n_5255)
);

AOI21xp5_ASAP7_75t_L g5256 ( 
.A1(n_4654),
.A2(n_3859),
.B(n_2648),
.Y(n_5256)
);

AOI21xp5_ASAP7_75t_L g5257 ( 
.A1(n_4667),
.A2(n_4061),
.B(n_3417),
.Y(n_5257)
);

AND2x6_ASAP7_75t_SL g5258 ( 
.A(n_4899),
.B(n_1014),
.Y(n_5258)
);

AOI21x1_ASAP7_75t_L g5259 ( 
.A1(n_4888),
.A2(n_4061),
.B(n_3259),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_4882),
.B(n_2292),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_4538),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_4499),
.Y(n_5262)
);

INVx2_ASAP7_75t_SL g5263 ( 
.A(n_4752),
.Y(n_5263)
);

AOI22xp33_ASAP7_75t_L g5264 ( 
.A1(n_4764),
.A2(n_902),
.B1(n_976),
.B2(n_850),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_4882),
.B(n_2295),
.Y(n_5265)
);

NOR2xp67_ASAP7_75t_L g5266 ( 
.A(n_4850),
.B(n_3675),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_4542),
.Y(n_5267)
);

CKINVDCx8_ASAP7_75t_R g5268 ( 
.A(n_4682),
.Y(n_5268)
);

NOR2xp33_ASAP7_75t_L g5269 ( 
.A(n_4690),
.B(n_4807),
.Y(n_5269)
);

OR2x2_ASAP7_75t_L g5270 ( 
.A(n_4871),
.B(n_3382),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_SL g5271 ( 
.A(n_4736),
.B(n_4352),
.Y(n_5271)
);

AOI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_4667),
.A2(n_3496),
.B(n_3491),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_L g5273 ( 
.A(n_4792),
.B(n_2295),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_4825),
.B(n_2310),
.Y(n_5274)
);

OR2x6_ASAP7_75t_L g5275 ( 
.A(n_4693),
.B(n_4754),
.Y(n_5275)
);

INVx2_ASAP7_75t_L g5276 ( 
.A(n_4499),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_SL g5277 ( 
.A(n_4910),
.B(n_4352),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_4672),
.A2(n_3435),
.B(n_3382),
.Y(n_5278)
);

NAND3xp33_ASAP7_75t_L g5279 ( 
.A(n_4734),
.B(n_1018),
.C(n_1014),
.Y(n_5279)
);

INVx1_ASAP7_75t_SL g5280 ( 
.A(n_4615),
.Y(n_5280)
);

OAI22xp5_ASAP7_75t_L g5281 ( 
.A1(n_4689),
.A2(n_1022),
.B1(n_1024),
.B2(n_1018),
.Y(n_5281)
);

AND2x2_ASAP7_75t_SL g5282 ( 
.A(n_4729),
.B(n_1173),
.Y(n_5282)
);

NAND2xp5_ASAP7_75t_L g5283 ( 
.A(n_4825),
.B(n_4907),
.Y(n_5283)
);

BUFx4f_ASAP7_75t_L g5284 ( 
.A(n_4572),
.Y(n_5284)
);

OAI22xp5_ASAP7_75t_L g5285 ( 
.A1(n_4689),
.A2(n_1024),
.B1(n_1032),
.B2(n_1022),
.Y(n_5285)
);

AND2x2_ASAP7_75t_L g5286 ( 
.A(n_4635),
.B(n_1032),
.Y(n_5286)
);

INVxp67_ASAP7_75t_L g5287 ( 
.A(n_4779),
.Y(n_5287)
);

NOR2xp33_ASAP7_75t_R g5288 ( 
.A(n_4572),
.B(n_4599),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_4907),
.B(n_2310),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_SL g5290 ( 
.A(n_4910),
.B(n_3679),
.Y(n_5290)
);

AOI21xp5_ASAP7_75t_L g5291 ( 
.A1(n_4672),
.A2(n_3435),
.B(n_3259),
.Y(n_5291)
);

INVx3_ASAP7_75t_L g5292 ( 
.A(n_4816),
.Y(n_5292)
);

NOR2x1_ASAP7_75t_L g5293 ( 
.A(n_4773),
.B(n_3860),
.Y(n_5293)
);

AOI21xp5_ASAP7_75t_L g5294 ( 
.A1(n_4674),
.A2(n_3259),
.B(n_3254),
.Y(n_5294)
);

NAND2x1p5_ASAP7_75t_L g5295 ( 
.A(n_4592),
.B(n_3981),
.Y(n_5295)
);

INVx2_ASAP7_75t_L g5296 ( 
.A(n_4501),
.Y(n_5296)
);

AND2x4_ASAP7_75t_L g5297 ( 
.A(n_4533),
.B(n_3902),
.Y(n_5297)
);

OAI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_4505),
.A2(n_3865),
.B(n_3848),
.Y(n_5298)
);

AOI21xp5_ASAP7_75t_L g5299 ( 
.A1(n_4674),
.A2(n_3263),
.B(n_3254),
.Y(n_5299)
);

O2A1O1Ixp33_ASAP7_75t_L g5300 ( 
.A1(n_4529),
.A2(n_1038),
.B(n_1041),
.C(n_1033),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_4913),
.B(n_2317),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_4913),
.B(n_2317),
.Y(n_5302)
);

BUFx2_ASAP7_75t_L g5303 ( 
.A(n_4535),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_4521),
.B(n_2337),
.Y(n_5304)
);

INVx2_ASAP7_75t_L g5305 ( 
.A(n_4501),
.Y(n_5305)
);

NOR2xp33_ASAP7_75t_L g5306 ( 
.A(n_4635),
.B(n_1335),
.Y(n_5306)
);

AOI21xp5_ASAP7_75t_L g5307 ( 
.A1(n_4696),
.A2(n_3263),
.B(n_3254),
.Y(n_5307)
);

AO21x1_ASAP7_75t_L g5308 ( 
.A1(n_4732),
.A2(n_1038),
.B(n_1033),
.Y(n_5308)
);

O2A1O1Ixp33_ASAP7_75t_L g5309 ( 
.A1(n_4884),
.A2(n_1044),
.B(n_1047),
.C(n_1041),
.Y(n_5309)
);

AOI21x1_ASAP7_75t_L g5310 ( 
.A1(n_4862),
.A2(n_4822),
.B(n_4619),
.Y(n_5310)
);

O2A1O1Ixp33_ASAP7_75t_L g5311 ( 
.A1(n_4885),
.A2(n_1047),
.B(n_1048),
.C(n_1044),
.Y(n_5311)
);

BUFx3_ASAP7_75t_L g5312 ( 
.A(n_4773),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_4521),
.B(n_2337),
.Y(n_5313)
);

NOR2xp33_ASAP7_75t_L g5314 ( 
.A(n_4635),
.B(n_1335),
.Y(n_5314)
);

AOI22x1_ASAP7_75t_L g5315 ( 
.A1(n_4847),
.A2(n_3803),
.B1(n_3772),
.B2(n_1063),
.Y(n_5315)
);

AOI21xp5_ASAP7_75t_L g5316 ( 
.A1(n_4696),
.A2(n_3265),
.B(n_3263),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4544),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_4596),
.B(n_2338),
.Y(n_5318)
);

OAI22xp5_ASAP7_75t_L g5319 ( 
.A1(n_4548),
.A2(n_1055),
.B1(n_1061),
.B2(n_1048),
.Y(n_5319)
);

NAND2xp5_ASAP7_75t_L g5320 ( 
.A(n_4596),
.B(n_2338),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4576),
.Y(n_5321)
);

AOI21xp5_ASAP7_75t_L g5322 ( 
.A1(n_4699),
.A2(n_3266),
.B(n_3265),
.Y(n_5322)
);

A2O1A1Ixp33_ASAP7_75t_L g5323 ( 
.A1(n_4591),
.A2(n_1061),
.B(n_1064),
.C(n_1055),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_4600),
.B(n_2339),
.Y(n_5324)
);

AOI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_4699),
.A2(n_3266),
.B(n_3265),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_4600),
.B(n_2339),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_SL g5327 ( 
.A(n_4910),
.B(n_3772),
.Y(n_5327)
);

AOI21x1_ASAP7_75t_L g5328 ( 
.A1(n_4862),
.A2(n_3268),
.B(n_3266),
.Y(n_5328)
);

BUFx2_ASAP7_75t_L g5329 ( 
.A(n_4535),
.Y(n_5329)
);

OAI21xp5_ASAP7_75t_L g5330 ( 
.A1(n_4735),
.A2(n_3865),
.B(n_3848),
.Y(n_5330)
);

O2A1O1Ixp33_ASAP7_75t_L g5331 ( 
.A1(n_4894),
.A2(n_1070),
.B(n_1076),
.C(n_1064),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_4652),
.Y(n_5332)
);

AOI21x1_ASAP7_75t_L g5333 ( 
.A1(n_4822),
.A2(n_3272),
.B(n_3268),
.Y(n_5333)
);

AOI21xp5_ASAP7_75t_L g5334 ( 
.A1(n_4703),
.A2(n_3272),
.B(n_3268),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_4669),
.B(n_2342),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4669),
.B(n_2342),
.Y(n_5336)
);

INVx5_ASAP7_75t_L g5337 ( 
.A(n_4509),
.Y(n_5337)
);

A2O1A1Ixp33_ASAP7_75t_L g5338 ( 
.A1(n_4591),
.A2(n_1076),
.B(n_1083),
.C(n_1070),
.Y(n_5338)
);

HB1xp67_ASAP7_75t_L g5339 ( 
.A(n_4615),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_SL g5340 ( 
.A(n_4635),
.B(n_4642),
.Y(n_5340)
);

AOI21xp5_ASAP7_75t_L g5341 ( 
.A1(n_4703),
.A2(n_3277),
.B(n_3272),
.Y(n_5341)
);

AOI21x1_ASAP7_75t_L g5342 ( 
.A1(n_4593),
.A2(n_3278),
.B(n_3277),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_4864),
.B(n_2353),
.Y(n_5343)
);

BUFx4f_ASAP7_75t_L g5344 ( 
.A(n_4572),
.Y(n_5344)
);

AOI22xp33_ASAP7_75t_L g5345 ( 
.A1(n_4635),
.A2(n_902),
.B1(n_976),
.B2(n_850),
.Y(n_5345)
);

NOR2xp33_ASAP7_75t_L g5346 ( 
.A(n_4642),
.B(n_4679),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_SL g5347 ( 
.A(n_4642),
.B(n_3803),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_SL g5348 ( 
.A(n_4642),
.B(n_4047),
.Y(n_5348)
);

NAND2xp5_ASAP7_75t_L g5349 ( 
.A(n_4581),
.B(n_4587),
.Y(n_5349)
);

INVx3_ASAP7_75t_SL g5350 ( 
.A(n_4599),
.Y(n_5350)
);

NAND2xp33_ASAP7_75t_L g5351 ( 
.A(n_4599),
.B(n_3848),
.Y(n_5351)
);

AOI21x1_ASAP7_75t_L g5352 ( 
.A1(n_4593),
.A2(n_3278),
.B(n_3277),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_4624),
.A2(n_3505),
.B1(n_3508),
.B2(n_3504),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4655),
.Y(n_5354)
);

O2A1O1Ixp33_ASAP7_75t_L g5355 ( 
.A1(n_4928),
.A2(n_1087),
.B(n_1090),
.C(n_1083),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_4936),
.Y(n_5356)
);

OR2x2_ASAP7_75t_L g5357 ( 
.A(n_5002),
.B(n_4504),
.Y(n_5357)
);

INVx2_ASAP7_75t_SL g5358 ( 
.A(n_4915),
.Y(n_5358)
);

OAI22xp33_ASAP7_75t_L g5359 ( 
.A1(n_5012),
.A2(n_4624),
.B1(n_4754),
.B2(n_4693),
.Y(n_5359)
);

AOI21xp5_ASAP7_75t_L g5360 ( 
.A1(n_4926),
.A2(n_4743),
.B(n_4729),
.Y(n_5360)
);

INVx2_ASAP7_75t_L g5361 ( 
.A(n_4917),
.Y(n_5361)
);

INVx2_ASAP7_75t_L g5362 ( 
.A(n_4921),
.Y(n_5362)
);

AOI21xp5_ASAP7_75t_L g5363 ( 
.A1(n_4939),
.A2(n_4743),
.B(n_4512),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_5002),
.B(n_4879),
.Y(n_5364)
);

BUFx2_ASAP7_75t_L g5365 ( 
.A(n_4914),
.Y(n_5365)
);

NOR2xp33_ASAP7_75t_L g5366 ( 
.A(n_4923),
.B(n_4642),
.Y(n_5366)
);

INVx2_ASAP7_75t_L g5367 ( 
.A(n_4945),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_4990),
.Y(n_5368)
);

AO21x1_ASAP7_75t_L g5369 ( 
.A1(n_5281),
.A2(n_4661),
.B(n_4658),
.Y(n_5369)
);

NOR2x1_ASAP7_75t_L g5370 ( 
.A(n_5070),
.B(n_4668),
.Y(n_5370)
);

NOR2xp33_ASAP7_75t_SL g5371 ( 
.A(n_5282),
.B(n_5234),
.Y(n_5371)
);

NAND2x1p5_ASAP7_75t_L g5372 ( 
.A(n_5337),
.B(n_4509),
.Y(n_5372)
);

AOI22x1_ASAP7_75t_L g5373 ( 
.A1(n_4942),
.A2(n_4847),
.B1(n_4624),
.B2(n_4681),
.Y(n_5373)
);

AOI21xp5_ASAP7_75t_L g5374 ( 
.A1(n_5097),
.A2(n_4512),
.B(n_4509),
.Y(n_5374)
);

AOI21xp5_ASAP7_75t_L g5375 ( 
.A1(n_5351),
.A2(n_4512),
.B(n_4509),
.Y(n_5375)
);

INVx3_ASAP7_75t_L g5376 ( 
.A(n_5023),
.Y(n_5376)
);

NOR2xp33_ASAP7_75t_R g5377 ( 
.A(n_4987),
.B(n_4599),
.Y(n_5377)
);

BUFx8_ASAP7_75t_L g5378 ( 
.A(n_4961),
.Y(n_5378)
);

HB1xp67_ASAP7_75t_L g5379 ( 
.A(n_5033),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_4995),
.Y(n_5380)
);

AOI21xp5_ASAP7_75t_L g5381 ( 
.A1(n_4976),
.A2(n_4512),
.B(n_4509),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_4972),
.Y(n_5382)
);

NAND2xp5_ASAP7_75t_L g5383 ( 
.A(n_5071),
.B(n_4879),
.Y(n_5383)
);

NAND2xp33_ASAP7_75t_L g5384 ( 
.A(n_4916),
.B(n_4599),
.Y(n_5384)
);

A2O1A1Ixp33_ASAP7_75t_L g5385 ( 
.A1(n_4934),
.A2(n_4693),
.B(n_4754),
.C(n_4533),
.Y(n_5385)
);

NAND2x1_ASAP7_75t_L g5386 ( 
.A(n_5275),
.B(n_4592),
.Y(n_5386)
);

NAND3xp33_ASAP7_75t_SL g5387 ( 
.A(n_5235),
.B(n_4625),
.C(n_4622),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_4951),
.B(n_4879),
.Y(n_5388)
);

A2O1A1Ixp33_ASAP7_75t_L g5389 ( 
.A1(n_4965),
.A2(n_4754),
.B(n_4693),
.C(n_4630),
.Y(n_5389)
);

INVx2_ASAP7_75t_SL g5390 ( 
.A(n_4915),
.Y(n_5390)
);

AOI21xp5_ASAP7_75t_L g5391 ( 
.A1(n_4973),
.A2(n_4512),
.B(n_4710),
.Y(n_5391)
);

OAI21xp5_ASAP7_75t_L g5392 ( 
.A1(n_5279),
.A2(n_4598),
.B(n_4857),
.Y(n_5392)
);

INVx2_ASAP7_75t_L g5393 ( 
.A(n_4980),
.Y(n_5393)
);

AOI21xp5_ASAP7_75t_L g5394 ( 
.A1(n_4974),
.A2(n_4711),
.B(n_4710),
.Y(n_5394)
);

AOI21xp5_ASAP7_75t_L g5395 ( 
.A1(n_5003),
.A2(n_4719),
.B(n_4711),
.Y(n_5395)
);

NAND2x1p5_ASAP7_75t_L g5396 ( 
.A(n_5337),
.B(n_4754),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5011),
.Y(n_5397)
);

O2A1O1Ixp33_ASAP7_75t_L g5398 ( 
.A1(n_5281),
.A2(n_1090),
.B(n_1096),
.C(n_1087),
.Y(n_5398)
);

INVx2_ASAP7_75t_L g5399 ( 
.A(n_5013),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_5058),
.Y(n_5400)
);

NAND2xp5_ASAP7_75t_L g5401 ( 
.A(n_4933),
.B(n_4879),
.Y(n_5401)
);

AOI21xp5_ASAP7_75t_L g5402 ( 
.A1(n_5291),
.A2(n_4977),
.B(n_5092),
.Y(n_5402)
);

AOI21xp5_ASAP7_75t_L g5403 ( 
.A1(n_5094),
.A2(n_4720),
.B(n_4719),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_SL g5404 ( 
.A(n_5093),
.B(n_4919),
.Y(n_5404)
);

AOI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_4994),
.A2(n_4722),
.B(n_4720),
.Y(n_5405)
);

OR2x2_ASAP7_75t_L g5406 ( 
.A(n_5280),
.B(n_4879),
.Y(n_5406)
);

NOR2xp33_ASAP7_75t_L g5407 ( 
.A(n_4996),
.B(n_4679),
.Y(n_5407)
);

NAND2xp5_ASAP7_75t_L g5408 ( 
.A(n_5019),
.B(n_5283),
.Y(n_5408)
);

BUFx10_ASAP7_75t_L g5409 ( 
.A(n_5168),
.Y(n_5409)
);

BUFx6f_ASAP7_75t_L g5410 ( 
.A(n_4915),
.Y(n_5410)
);

INVx6_ASAP7_75t_L g5411 ( 
.A(n_4953),
.Y(n_5411)
);

O2A1O1Ixp33_ASAP7_75t_L g5412 ( 
.A1(n_5285),
.A2(n_1100),
.B(n_1109),
.C(n_1096),
.Y(n_5412)
);

O2A1O1Ixp33_ASAP7_75t_SL g5413 ( 
.A1(n_5173),
.A2(n_1100),
.B(n_1113),
.C(n_1109),
.Y(n_5413)
);

A2O1A1Ixp33_ASAP7_75t_L g5414 ( 
.A1(n_5096),
.A2(n_4630),
.B(n_4592),
.C(n_1116),
.Y(n_5414)
);

OAI22xp5_ASAP7_75t_L g5415 ( 
.A1(n_5210),
.A2(n_4598),
.B1(n_4554),
.B2(n_4679),
.Y(n_5415)
);

A2O1A1Ixp33_ASAP7_75t_L g5416 ( 
.A1(n_4918),
.A2(n_4630),
.B(n_1116),
.C(n_1120),
.Y(n_5416)
);

AOI221xp5_ASAP7_75t_L g5417 ( 
.A1(n_5285),
.A2(n_1069),
.B1(n_1075),
.B2(n_1065),
.C(n_1062),
.Y(n_5417)
);

NAND2xp5_ASAP7_75t_SL g5418 ( 
.A(n_4958),
.B(n_4687),
.Y(n_5418)
);

AOI22xp33_ASAP7_75t_L g5419 ( 
.A1(n_5073),
.A2(n_4679),
.B1(n_1182),
.B2(n_1234),
.Y(n_5419)
);

AOI21xp5_ASAP7_75t_L g5420 ( 
.A1(n_5000),
.A2(n_4724),
.B(n_4722),
.Y(n_5420)
);

INVx4_ASAP7_75t_L g5421 ( 
.A(n_4932),
.Y(n_5421)
);

NAND2xp5_ASAP7_75t_L g5422 ( 
.A(n_4998),
.B(n_4510),
.Y(n_5422)
);

O2A1O1Ixp33_ASAP7_75t_L g5423 ( 
.A1(n_5248),
.A2(n_1120),
.B(n_1126),
.C(n_1124),
.Y(n_5423)
);

AND2x2_ASAP7_75t_L g5424 ( 
.A(n_5090),
.B(n_4510),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_SL g5425 ( 
.A(n_5279),
.B(n_4687),
.Y(n_5425)
);

AOI21xp5_ASAP7_75t_L g5426 ( 
.A1(n_5004),
.A2(n_4725),
.B(n_4724),
.Y(n_5426)
);

NAND2xp5_ASAP7_75t_SL g5427 ( 
.A(n_4944),
.B(n_4687),
.Y(n_5427)
);

NOR2xp33_ASAP7_75t_L g5428 ( 
.A(n_4941),
.B(n_4679),
.Y(n_5428)
);

NOR2xp33_ASAP7_75t_L g5429 ( 
.A(n_4970),
.B(n_4563),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_5198),
.B(n_4671),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5157),
.B(n_4704),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_4978),
.B(n_4991),
.Y(n_5432)
);

AOI22xp5_ASAP7_75t_L g5433 ( 
.A1(n_5216),
.A2(n_1124),
.B1(n_1126),
.B2(n_1113),
.Y(n_5433)
);

NAND3xp33_ASAP7_75t_SL g5434 ( 
.A(n_4940),
.B(n_4627),
.C(n_1078),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5065),
.Y(n_5435)
);

AOI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_5032),
.A2(n_4738),
.B(n_4725),
.Y(n_5436)
);

NAND2xp5_ASAP7_75t_L g5437 ( 
.A(n_5339),
.B(n_4706),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5050),
.Y(n_5438)
);

AOI21xp5_ASAP7_75t_L g5439 ( 
.A1(n_5032),
.A2(n_4738),
.B(n_4746),
.Y(n_5439)
);

NAND2xp5_ASAP7_75t_L g5440 ( 
.A(n_4925),
.B(n_4712),
.Y(n_5440)
);

AOI21xp5_ASAP7_75t_L g5441 ( 
.A1(n_5034),
.A2(n_4747),
.B(n_4746),
.Y(n_5441)
);

AOI21xp5_ASAP7_75t_L g5442 ( 
.A1(n_5034),
.A2(n_4748),
.B(n_4747),
.Y(n_5442)
);

BUFx3_ASAP7_75t_L g5443 ( 
.A(n_4932),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_SL g5444 ( 
.A(n_4943),
.B(n_4701),
.Y(n_5444)
);

NAND2xp5_ASAP7_75t_L g5445 ( 
.A(n_5108),
.B(n_4770),
.Y(n_5445)
);

AOI21xp5_ASAP7_75t_L g5446 ( 
.A1(n_5008),
.A2(n_4750),
.B(n_4748),
.Y(n_5446)
);

O2A1O1Ixp33_ASAP7_75t_L g5447 ( 
.A1(n_5061),
.A2(n_1130),
.B(n_1131),
.C(n_1129),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_SL g5448 ( 
.A(n_4949),
.B(n_4701),
.Y(n_5448)
);

AOI22xp33_ASAP7_75t_SL g5449 ( 
.A1(n_5102),
.A2(n_4609),
.B1(n_4604),
.B2(n_4857),
.Y(n_5449)
);

CKINVDCx14_ASAP7_75t_R g5450 ( 
.A(n_5240),
.Y(n_5450)
);

AOI21xp5_ASAP7_75t_L g5451 ( 
.A1(n_5278),
.A2(n_4756),
.B(n_4750),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_5084),
.Y(n_5452)
);

OAI22xp5_ASAP7_75t_SL g5453 ( 
.A1(n_4967),
.A2(n_4829),
.B1(n_4853),
.B2(n_4819),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5085),
.Y(n_5454)
);

OAI22xp5_ASAP7_75t_L g5455 ( 
.A1(n_5280),
.A2(n_4947),
.B1(n_5264),
.B2(n_5345),
.Y(n_5455)
);

AOI21xp5_ASAP7_75t_L g5456 ( 
.A1(n_5256),
.A2(n_4776),
.B(n_4756),
.Y(n_5456)
);

NOR3xp33_ASAP7_75t_SL g5457 ( 
.A(n_4971),
.B(n_1080),
.C(n_1077),
.Y(n_5457)
);

INVx3_ASAP7_75t_L g5458 ( 
.A(n_5023),
.Y(n_5458)
);

A2O1A1Ixp33_ASAP7_75t_L g5459 ( 
.A1(n_5079),
.A2(n_1130),
.B(n_1131),
.C(n_1129),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5141),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5151),
.Y(n_5461)
);

INVxp67_ASAP7_75t_L g5462 ( 
.A(n_5212),
.Y(n_5462)
);

AOI22xp33_ASAP7_75t_L g5463 ( 
.A1(n_4946),
.A2(n_1182),
.B1(n_1234),
.B2(n_1178),
.Y(n_5463)
);

INVx2_ASAP7_75t_L g5464 ( 
.A(n_5078),
.Y(n_5464)
);

OAI22xp5_ASAP7_75t_L g5465 ( 
.A1(n_5038),
.A2(n_4598),
.B1(n_4554),
.B2(n_4855),
.Y(n_5465)
);

AOI21xp5_ASAP7_75t_L g5466 ( 
.A1(n_5051),
.A2(n_4776),
.B(n_4854),
.Y(n_5466)
);

O2A1O1Ixp33_ASAP7_75t_L g5467 ( 
.A1(n_5112),
.A2(n_1139),
.B(n_1143),
.C(n_1135),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5152),
.Y(n_5468)
);

OAI21x1_ASAP7_75t_L g5469 ( 
.A1(n_5333),
.A2(n_4673),
.B(n_4649),
.Y(n_5469)
);

NOR2xp33_ASAP7_75t_L g5470 ( 
.A(n_5017),
.B(n_4563),
.Y(n_5470)
);

INVx3_ASAP7_75t_L g5471 ( 
.A(n_5066),
.Y(n_5471)
);

NOR2xp33_ASAP7_75t_L g5472 ( 
.A(n_5024),
.B(n_4570),
.Y(n_5472)
);

AND2x6_ASAP7_75t_SL g5473 ( 
.A(n_5136),
.B(n_1135),
.Y(n_5473)
);

INVx2_ASAP7_75t_SL g5474 ( 
.A(n_4932),
.Y(n_5474)
);

A2O1A1Ixp33_ASAP7_75t_L g5475 ( 
.A1(n_5089),
.A2(n_5006),
.B(n_5104),
.C(n_5309),
.Y(n_5475)
);

NAND2x1_ASAP7_75t_L g5476 ( 
.A(n_5275),
.B(n_4857),
.Y(n_5476)
);

O2A1O1Ixp33_ASAP7_75t_L g5477 ( 
.A1(n_5109),
.A2(n_1143),
.B(n_1144),
.C(n_1139),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_5155),
.Y(n_5478)
);

NAND2xp5_ASAP7_75t_L g5479 ( 
.A(n_5114),
.B(n_4893),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5164),
.Y(n_5480)
);

A2O1A1Ixp33_ASAP7_75t_L g5481 ( 
.A1(n_5311),
.A2(n_1147),
.B(n_1148),
.C(n_1144),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_SL g5482 ( 
.A(n_5009),
.B(n_4701),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5030),
.B(n_5043),
.Y(n_5483)
);

OR2x2_ASAP7_75t_L g5484 ( 
.A(n_5270),
.B(n_4492),
.Y(n_5484)
);

OAI22xp5_ASAP7_75t_L g5485 ( 
.A1(n_5059),
.A2(n_4554),
.B1(n_4609),
.B2(n_4604),
.Y(n_5485)
);

OAI22xp5_ASAP7_75t_L g5486 ( 
.A1(n_5125),
.A2(n_4609),
.B1(n_4604),
.B2(n_4781),
.Y(n_5486)
);

INVx2_ASAP7_75t_L g5487 ( 
.A(n_5098),
.Y(n_5487)
);

NOR2xp67_ASAP7_75t_SL g5488 ( 
.A(n_5249),
.B(n_4604),
.Y(n_5488)
);

AOI21xp5_ASAP7_75t_L g5489 ( 
.A1(n_5054),
.A2(n_5060),
.B(n_5247),
.Y(n_5489)
);

AOI21xp5_ASAP7_75t_L g5490 ( 
.A1(n_5251),
.A2(n_4854),
.B(n_4555),
.Y(n_5490)
);

INVx3_ASAP7_75t_L g5491 ( 
.A(n_5066),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_SL g5492 ( 
.A(n_5009),
.B(n_4604),
.Y(n_5492)
);

O2A1O1Ixp5_ASAP7_75t_L g5493 ( 
.A1(n_5042),
.A2(n_4649),
.B(n_4677),
.C(n_4673),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_L g5494 ( 
.A(n_5086),
.B(n_4893),
.Y(n_5494)
);

NOR2xp33_ASAP7_75t_SL g5495 ( 
.A(n_5268),
.B(n_4609),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5088),
.B(n_4895),
.Y(n_5496)
);

AOI22xp5_ASAP7_75t_L g5497 ( 
.A1(n_4950),
.A2(n_1148),
.B1(n_1151),
.B2(n_1147),
.Y(n_5497)
);

O2A1O1Ixp33_ASAP7_75t_L g5498 ( 
.A1(n_5323),
.A2(n_1152),
.B(n_1153),
.C(n_1151),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_SL g5499 ( 
.A(n_5009),
.B(n_4609),
.Y(n_5499)
);

AOI21xp5_ASAP7_75t_L g5500 ( 
.A1(n_5257),
.A2(n_4555),
.B(n_4886),
.Y(n_5500)
);

AOI21xp5_ASAP7_75t_L g5501 ( 
.A1(n_4964),
.A2(n_4886),
.B(n_4492),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_5007),
.B(n_4895),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_5252),
.A2(n_4896),
.B(n_4673),
.Y(n_5503)
);

O2A1O1Ixp33_ASAP7_75t_L g5504 ( 
.A1(n_5338),
.A2(n_1153),
.B(n_1156),
.C(n_1152),
.Y(n_5504)
);

OAI21x1_ASAP7_75t_L g5505 ( 
.A1(n_5310),
.A2(n_4677),
.B(n_4649),
.Y(n_5505)
);

AOI21xp5_ASAP7_75t_L g5506 ( 
.A1(n_4981),
.A2(n_4896),
.B(n_4718),
.Y(n_5506)
);

AND2x2_ASAP7_75t_SL g5507 ( 
.A(n_5137),
.B(n_4866),
.Y(n_5507)
);

NOR2x1_ASAP7_75t_L g5508 ( 
.A(n_5293),
.B(n_4513),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5177),
.Y(n_5509)
);

O2A1O1Ixp33_ASAP7_75t_L g5510 ( 
.A1(n_4989),
.A2(n_1168),
.B(n_1169),
.C(n_1156),
.Y(n_5510)
);

AOI21xp5_ASAP7_75t_L g5511 ( 
.A1(n_4983),
.A2(n_4718),
.B(n_4677),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5219),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5238),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_L g5514 ( 
.A(n_5048),
.B(n_4999),
.Y(n_5514)
);

INVx3_ASAP7_75t_L g5515 ( 
.A(n_5132),
.Y(n_5515)
);

NOR2xp33_ASAP7_75t_L g5516 ( 
.A(n_4935),
.B(n_4570),
.Y(n_5516)
);

INVx5_ASAP7_75t_L g5517 ( 
.A(n_5120),
.Y(n_5517)
);

NAND2xp5_ASAP7_75t_L g5518 ( 
.A(n_4993),
.B(n_4513),
.Y(n_5518)
);

AND2x6_ASAP7_75t_L g5519 ( 
.A(n_4920),
.B(n_4688),
.Y(n_5519)
);

AND2x4_ASAP7_75t_L g5520 ( 
.A(n_5277),
.B(n_4718),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_5261),
.Y(n_5521)
);

OAI22xp5_ASAP7_75t_L g5522 ( 
.A1(n_4968),
.A2(n_4603),
.B1(n_4612),
.B2(n_4601),
.Y(n_5522)
);

NOR2xp33_ASAP7_75t_L g5523 ( 
.A(n_5055),
.B(n_4584),
.Y(n_5523)
);

NOR2xp33_ASAP7_75t_L g5524 ( 
.A(n_5074),
.B(n_4584),
.Y(n_5524)
);

AND2x2_ASAP7_75t_L g5525 ( 
.A(n_4937),
.B(n_4688),
.Y(n_5525)
);

BUFx6f_ASAP7_75t_L g5526 ( 
.A(n_5053),
.Y(n_5526)
);

AOI21xp5_ASAP7_75t_L g5527 ( 
.A1(n_5142),
.A2(n_4740),
.B(n_4737),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5267),
.Y(n_5528)
);

A2O1A1Ixp33_ASAP7_75t_L g5529 ( 
.A1(n_5331),
.A2(n_1168),
.B(n_1169),
.C(n_1159),
.Y(n_5529)
);

INVxp67_ASAP7_75t_L g5530 ( 
.A(n_4922),
.Y(n_5530)
);

BUFx6f_ASAP7_75t_L g5531 ( 
.A(n_5228),
.Y(n_5531)
);

O2A1O1Ixp33_ASAP7_75t_L g5532 ( 
.A1(n_5116),
.A2(n_1177),
.B(n_1179),
.C(n_1159),
.Y(n_5532)
);

AO21x2_ASAP7_75t_L g5533 ( 
.A1(n_5069),
.A2(n_4832),
.B(n_4831),
.Y(n_5533)
);

NAND3xp33_ASAP7_75t_SL g5534 ( 
.A(n_5239),
.B(n_5314),
.C(n_5306),
.Y(n_5534)
);

BUFx6f_ASAP7_75t_L g5535 ( 
.A(n_5312),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_5317),
.Y(n_5536)
);

A2O1A1Ixp33_ASAP7_75t_L g5537 ( 
.A1(n_5037),
.A2(n_1179),
.B(n_1181),
.C(n_1177),
.Y(n_5537)
);

NAND2xp5_ASAP7_75t_L g5538 ( 
.A(n_5057),
.B(n_4777),
.Y(n_5538)
);

OAI22xp5_ASAP7_75t_L g5539 ( 
.A1(n_5101),
.A2(n_4603),
.B1(n_4612),
.B2(n_4601),
.Y(n_5539)
);

INVxp67_ASAP7_75t_L g5540 ( 
.A(n_4988),
.Y(n_5540)
);

O2A1O1Ixp33_ASAP7_75t_L g5541 ( 
.A1(n_5111),
.A2(n_1181),
.B(n_1187),
.C(n_1185),
.Y(n_5541)
);

AOI22xp33_ASAP7_75t_SL g5542 ( 
.A1(n_5254),
.A2(n_4857),
.B1(n_1530),
.B2(n_1577),
.Y(n_5542)
);

NOR2xp33_ASAP7_75t_L g5543 ( 
.A(n_5175),
.B(n_4611),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5321),
.Y(n_5544)
);

BUFx4f_ASAP7_75t_L g5545 ( 
.A(n_5146),
.Y(n_5545)
);

O2A1O1Ixp33_ASAP7_75t_L g5546 ( 
.A1(n_5111),
.A2(n_1187),
.B(n_1190),
.C(n_1185),
.Y(n_5546)
);

NOR2xp33_ASAP7_75t_L g5547 ( 
.A(n_5119),
.B(n_4611),
.Y(n_5547)
);

NAND2xp5_ASAP7_75t_L g5548 ( 
.A(n_5349),
.B(n_4777),
.Y(n_5548)
);

INVx3_ASAP7_75t_L g5549 ( 
.A(n_5132),
.Y(n_5549)
);

O2A1O1Ixp5_ASAP7_75t_L g5550 ( 
.A1(n_4979),
.A2(n_4740),
.B(n_4741),
.C(n_4737),
.Y(n_5550)
);

NOR2xp67_ASAP7_75t_SL g5551 ( 
.A(n_5337),
.B(n_4828),
.Y(n_5551)
);

INVx2_ASAP7_75t_SL g5552 ( 
.A(n_5062),
.Y(n_5552)
);

INVx4_ASAP7_75t_L g5553 ( 
.A(n_5350),
.Y(n_5553)
);

NAND2xp33_ASAP7_75t_SL g5554 ( 
.A(n_5288),
.B(n_4626),
.Y(n_5554)
);

O2A1O1Ixp33_ASAP7_75t_L g5555 ( 
.A1(n_5201),
.A2(n_5229),
.B(n_5163),
.C(n_5147),
.Y(n_5555)
);

NAND2xp5_ASAP7_75t_L g5556 ( 
.A(n_5197),
.B(n_4785),
.Y(n_5556)
);

NAND2xp5_ASAP7_75t_L g5557 ( 
.A(n_4924),
.B(n_4785),
.Y(n_5557)
);

NAND2xp5_ASAP7_75t_L g5558 ( 
.A(n_5118),
.B(n_4809),
.Y(n_5558)
);

AND2x4_ASAP7_75t_L g5559 ( 
.A(n_5275),
.B(n_4737),
.Y(n_5559)
);

NAND2xp5_ASAP7_75t_L g5560 ( 
.A(n_5287),
.B(n_4809),
.Y(n_5560)
);

NAND2xp5_ASAP7_75t_SL g5561 ( 
.A(n_5075),
.B(n_4866),
.Y(n_5561)
);

NOR2xp33_ASAP7_75t_L g5562 ( 
.A(n_5113),
.B(n_5176),
.Y(n_5562)
);

INVx3_ASAP7_75t_L g5563 ( 
.A(n_5292),
.Y(n_5563)
);

BUFx12f_ASAP7_75t_L g5564 ( 
.A(n_5227),
.Y(n_5564)
);

AOI21xp5_ASAP7_75t_L g5565 ( 
.A1(n_5158),
.A2(n_4741),
.B(n_4740),
.Y(n_5565)
);

CKINVDCx14_ASAP7_75t_R g5566 ( 
.A(n_5178),
.Y(n_5566)
);

NAND2xp5_ASAP7_75t_L g5567 ( 
.A(n_5180),
.B(n_5211),
.Y(n_5567)
);

NAND2xp5_ASAP7_75t_L g5568 ( 
.A(n_5080),
.B(n_4810),
.Y(n_5568)
);

O2A1O1Ixp5_ASAP7_75t_L g5569 ( 
.A1(n_5072),
.A2(n_4800),
.B(n_4803),
.C(n_4741),
.Y(n_5569)
);

NAND2xp5_ASAP7_75t_L g5570 ( 
.A(n_5081),
.B(n_5082),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_SL g5571 ( 
.A(n_5233),
.B(n_5263),
.Y(n_5571)
);

INVx3_ASAP7_75t_L g5572 ( 
.A(n_5292),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_L g5573 ( 
.A(n_5117),
.B(n_4810),
.Y(n_5573)
);

OR2x2_ASAP7_75t_L g5574 ( 
.A(n_5332),
.B(n_4821),
.Y(n_5574)
);

BUFx4f_ASAP7_75t_SL g5575 ( 
.A(n_5227),
.Y(n_5575)
);

AOI21xp5_ASAP7_75t_L g5576 ( 
.A1(n_5162),
.A2(n_5165),
.B(n_4927),
.Y(n_5576)
);

A2O1A1Ixp33_ASAP7_75t_L g5577 ( 
.A1(n_5300),
.A2(n_1203),
.B(n_1205),
.C(n_1190),
.Y(n_5577)
);

INVx2_ASAP7_75t_L g5578 ( 
.A(n_5354),
.Y(n_5578)
);

AO21x1_ASAP7_75t_L g5579 ( 
.A1(n_5319),
.A2(n_1205),
.B(n_1203),
.Y(n_5579)
);

NOR3xp33_ASAP7_75t_SL g5580 ( 
.A(n_5040),
.B(n_5199),
.C(n_5083),
.Y(n_5580)
);

NAND2xp5_ASAP7_75t_L g5581 ( 
.A(n_5242),
.B(n_4821),
.Y(n_5581)
);

OAI22xp5_ASAP7_75t_L g5582 ( 
.A1(n_5015),
.A2(n_4817),
.B1(n_4781),
.B2(n_4845),
.Y(n_5582)
);

AOI21xp5_ASAP7_75t_L g5583 ( 
.A1(n_4930),
.A2(n_4803),
.B(n_4800),
.Y(n_5583)
);

O2A1O1Ixp5_ASAP7_75t_SL g5584 ( 
.A1(n_5129),
.A2(n_1208),
.B(n_1216),
.C(n_1206),
.Y(n_5584)
);

BUFx3_ASAP7_75t_L g5585 ( 
.A(n_5110),
.Y(n_5585)
);

O2A1O1Ixp33_ASAP7_75t_L g5586 ( 
.A1(n_4975),
.A2(n_1208),
.B(n_1216),
.C(n_1206),
.Y(n_5586)
);

NOR2xp33_ASAP7_75t_R g5587 ( 
.A(n_5128),
.B(n_4623),
.Y(n_5587)
);

OAI22xp5_ASAP7_75t_L g5588 ( 
.A1(n_5036),
.A2(n_4817),
.B1(n_4845),
.B2(n_4815),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_5130),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5160),
.Y(n_5590)
);

OR2x6_ASAP7_75t_L g5591 ( 
.A(n_4948),
.B(n_4800),
.Y(n_5591)
);

OR2x2_ASAP7_75t_L g5592 ( 
.A(n_5067),
.B(n_5289),
.Y(n_5592)
);

O2A1O1Ixp33_ASAP7_75t_L g5593 ( 
.A1(n_5319),
.A2(n_5091),
.B(n_5183),
.C(n_5135),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_5223),
.Y(n_5594)
);

CKINVDCx5p33_ASAP7_75t_R g5595 ( 
.A(n_5231),
.Y(n_5595)
);

AOI22xp33_ASAP7_75t_L g5596 ( 
.A1(n_4956),
.A2(n_1182),
.B1(n_1234),
.B2(n_1178),
.Y(n_5596)
);

NOR2xp33_ASAP7_75t_L g5597 ( 
.A(n_5269),
.B(n_4623),
.Y(n_5597)
);

A2O1A1Ixp33_ASAP7_75t_L g5598 ( 
.A1(n_5330),
.A2(n_1217),
.B(n_1223),
.C(n_1218),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5236),
.Y(n_5599)
);

NAND3xp33_ASAP7_75t_SL g5600 ( 
.A(n_5189),
.B(n_1084),
.C(n_1082),
.Y(n_5600)
);

AOI21xp5_ASAP7_75t_L g5601 ( 
.A1(n_4984),
.A2(n_4818),
.B(n_4803),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_4953),
.Y(n_5602)
);

NOR2xp33_ASAP7_75t_L g5603 ( 
.A(n_5181),
.B(n_4643),
.Y(n_5603)
);

OA22x2_ASAP7_75t_L g5604 ( 
.A1(n_5194),
.A2(n_4845),
.B1(n_4557),
.B2(n_4558),
.Y(n_5604)
);

NAND2xp5_ASAP7_75t_SL g5605 ( 
.A(n_5260),
.B(n_4866),
.Y(n_5605)
);

BUFx6f_ASAP7_75t_L g5606 ( 
.A(n_5146),
.Y(n_5606)
);

AND2x2_ASAP7_75t_L g5607 ( 
.A(n_4997),
.B(n_5046),
.Y(n_5607)
);

AND2x2_ASAP7_75t_L g5608 ( 
.A(n_5052),
.B(n_4694),
.Y(n_5608)
);

NOR2xp33_ASAP7_75t_L g5609 ( 
.A(n_5185),
.B(n_4643),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_L g5610 ( 
.A(n_5063),
.B(n_4826),
.Y(n_5610)
);

AOI22xp5_ASAP7_75t_L g5611 ( 
.A1(n_5286),
.A2(n_1217),
.B1(n_1223),
.B2(n_1218),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5262),
.Y(n_5612)
);

O2A1O1Ixp5_ASAP7_75t_L g5613 ( 
.A1(n_5077),
.A2(n_4842),
.B(n_4861),
.C(n_4818),
.Y(n_5613)
);

NOR2xp33_ASAP7_75t_L g5614 ( 
.A(n_5056),
.B(n_4816),
.Y(n_5614)
);

AND2x2_ASAP7_75t_L g5615 ( 
.A(n_5064),
.B(n_4694),
.Y(n_5615)
);

AOI21xp5_ASAP7_75t_L g5616 ( 
.A1(n_4984),
.A2(n_4842),
.B(n_4818),
.Y(n_5616)
);

BUFx6f_ASAP7_75t_L g5617 ( 
.A(n_5146),
.Y(n_5617)
);

NOR2xp67_ASAP7_75t_L g5618 ( 
.A(n_4959),
.B(n_4842),
.Y(n_5618)
);

INVxp67_ASAP7_75t_L g5619 ( 
.A(n_5250),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_SL g5620 ( 
.A(n_5265),
.B(n_4709),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_5167),
.A2(n_4865),
.B(n_4861),
.Y(n_5621)
);

NAND2xp5_ASAP7_75t_L g5622 ( 
.A(n_5301),
.B(n_4826),
.Y(n_5622)
);

O2A1O1Ixp33_ASAP7_75t_SL g5623 ( 
.A1(n_5154),
.A2(n_1225),
.B(n_1230),
.C(n_1224),
.Y(n_5623)
);

NAND2xp5_ASAP7_75t_SL g5624 ( 
.A(n_5134),
.B(n_4709),
.Y(n_5624)
);

AND2x2_ASAP7_75t_L g5625 ( 
.A(n_5145),
.B(n_4714),
.Y(n_5625)
);

AOI21xp5_ASAP7_75t_L g5626 ( 
.A1(n_5217),
.A2(n_4865),
.B(n_4861),
.Y(n_5626)
);

BUFx2_ASAP7_75t_L g5627 ( 
.A(n_5303),
.Y(n_5627)
);

OAI21x1_ASAP7_75t_L g5628 ( 
.A1(n_5047),
.A2(n_4897),
.B(n_4865),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5276),
.Y(n_5629)
);

NOR2xp33_ASAP7_75t_L g5630 ( 
.A(n_5143),
.B(n_4823),
.Y(n_5630)
);

O2A1O1Ixp33_ASAP7_75t_L g5631 ( 
.A1(n_4966),
.A2(n_1230),
.B(n_1237),
.C(n_1225),
.Y(n_5631)
);

NAND2xp5_ASAP7_75t_L g5632 ( 
.A(n_5302),
.B(n_4714),
.Y(n_5632)
);

AOI21xp5_ASAP7_75t_L g5633 ( 
.A1(n_5169),
.A2(n_4905),
.B(n_4897),
.Y(n_5633)
);

BUFx2_ASAP7_75t_L g5634 ( 
.A(n_5329),
.Y(n_5634)
);

NAND2x1p5_ASAP7_75t_L g5635 ( 
.A(n_5337),
.B(n_4897),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5296),
.Y(n_5636)
);

AOI21xp5_ASAP7_75t_L g5637 ( 
.A1(n_5170),
.A2(n_4905),
.B(n_4723),
.Y(n_5637)
);

NAND2xp5_ASAP7_75t_L g5638 ( 
.A(n_5031),
.B(n_4857),
.Y(n_5638)
);

AOI21xp5_ASAP7_75t_L g5639 ( 
.A1(n_5014),
.A2(n_4905),
.B(n_4723),
.Y(n_5639)
);

AOI21xp5_ASAP7_75t_L g5640 ( 
.A1(n_5016),
.A2(n_4742),
.B(n_4715),
.Y(n_5640)
);

OAI21xp5_ASAP7_75t_L g5641 ( 
.A1(n_4966),
.A2(n_4742),
.B(n_4715),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_5039),
.B(n_4581),
.Y(n_5642)
);

NOR2x1_ASAP7_75t_L g5643 ( 
.A(n_5335),
.B(n_4650),
.Y(n_5643)
);

AOI21xp5_ASAP7_75t_L g5644 ( 
.A1(n_4960),
.A2(n_4580),
.B(n_4794),
.Y(n_5644)
);

NOR2xp33_ASAP7_75t_SL g5645 ( 
.A(n_4962),
.B(n_4650),
.Y(n_5645)
);

OAI22x1_ASAP7_75t_L g5646 ( 
.A1(n_4948),
.A2(n_1241),
.B1(n_1245),
.B2(n_1237),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_5305),
.Y(n_5647)
);

OAI21xp5_ASAP7_75t_L g5648 ( 
.A1(n_4955),
.A2(n_4590),
.B(n_4587),
.Y(n_5648)
);

NOR2xp33_ASAP7_75t_L g5649 ( 
.A(n_5153),
.B(n_5232),
.Y(n_5649)
);

NAND2xp5_ASAP7_75t_L g5650 ( 
.A(n_5005),
.B(n_4590),
.Y(n_5650)
);

INVx8_ASAP7_75t_L g5651 ( 
.A(n_4957),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_5221),
.Y(n_5652)
);

AOI21xp5_ASAP7_75t_L g5653 ( 
.A1(n_5005),
.A2(n_4797),
.B(n_4794),
.Y(n_5653)
);

AOI21xp5_ASAP7_75t_L g5654 ( 
.A1(n_4955),
.A2(n_4798),
.B(n_4797),
.Y(n_5654)
);

NOR2xp33_ASAP7_75t_L g5655 ( 
.A(n_5001),
.B(n_4823),
.Y(n_5655)
);

NAND2xp5_ASAP7_75t_SL g5656 ( 
.A(n_5099),
.B(n_4823),
.Y(n_5656)
);

AND2x4_ASAP7_75t_SL g5657 ( 
.A(n_5021),
.B(n_4823),
.Y(n_5657)
);

XOR2xp5_ASAP7_75t_L g5658 ( 
.A(n_5099),
.B(n_4823),
.Y(n_5658)
);

O2A1O1Ixp33_ASAP7_75t_L g5659 ( 
.A1(n_5161),
.A2(n_1247),
.B(n_1259),
.C(n_1245),
.Y(n_5659)
);

AOI21xp5_ASAP7_75t_L g5660 ( 
.A1(n_4938),
.A2(n_4798),
.B(n_4628),
.Y(n_5660)
);

AOI21x1_ASAP7_75t_L g5661 ( 
.A1(n_5018),
.A2(n_4628),
.B(n_4626),
.Y(n_5661)
);

INVx2_ASAP7_75t_L g5662 ( 
.A(n_5041),
.Y(n_5662)
);

BUFx4_ASAP7_75t_SL g5663 ( 
.A(n_5258),
.Y(n_5663)
);

INVx2_ASAP7_75t_L g5664 ( 
.A(n_5044),
.Y(n_5664)
);

BUFx2_ASAP7_75t_L g5665 ( 
.A(n_5149),
.Y(n_5665)
);

INVx3_ASAP7_75t_L g5666 ( 
.A(n_5149),
.Y(n_5666)
);

OAI22x1_ASAP7_75t_L g5667 ( 
.A1(n_5174),
.A2(n_1259),
.B1(n_1271),
.B2(n_1247),
.Y(n_5667)
);

O2A1O1Ixp5_ASAP7_75t_SL g5668 ( 
.A1(n_5340),
.A2(n_1241),
.B(n_1271),
.C(n_1224),
.Y(n_5668)
);

BUFx6f_ASAP7_75t_L g5669 ( 
.A(n_5149),
.Y(n_5669)
);

AOI22xp33_ASAP7_75t_L g5670 ( 
.A1(n_5308),
.A2(n_1282),
.B1(n_1178),
.B2(n_1275),
.Y(n_5670)
);

NAND2xp5_ASAP7_75t_SL g5671 ( 
.A(n_5304),
.B(n_4828),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5221),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5221),
.Y(n_5673)
);

AOI21xp5_ASAP7_75t_L g5674 ( 
.A1(n_4929),
.A2(n_4632),
.B(n_4631),
.Y(n_5674)
);

AND2x2_ASAP7_75t_L g5675 ( 
.A(n_5171),
.B(n_4831),
.Y(n_5675)
);

NAND2xp5_ASAP7_75t_L g5676 ( 
.A(n_5182),
.B(n_4832),
.Y(n_5676)
);

AOI21xp5_ASAP7_75t_L g5677 ( 
.A1(n_4952),
.A2(n_4632),
.B(n_4631),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_5190),
.Y(n_5678)
);

NOR3xp33_ASAP7_75t_L g5679 ( 
.A(n_5313),
.B(n_1275),
.C(n_1272),
.Y(n_5679)
);

NAND2x1p5_ASAP7_75t_L g5680 ( 
.A(n_5103),
.B(n_5208),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_5200),
.B(n_4634),
.Y(n_5681)
);

NAND2xp5_ASAP7_75t_SL g5682 ( 
.A(n_5273),
.B(n_5274),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5336),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5259),
.Y(n_5684)
);

AOI21xp5_ASAP7_75t_L g5685 ( 
.A1(n_5020),
.A2(n_4637),
.B(n_4634),
.Y(n_5685)
);

OAI22xp5_ASAP7_75t_L g5686 ( 
.A1(n_5222),
.A2(n_4828),
.B1(n_4640),
.B2(n_4653),
.Y(n_5686)
);

BUFx12f_ASAP7_75t_L g5687 ( 
.A(n_5159),
.Y(n_5687)
);

BUFx6f_ASAP7_75t_L g5688 ( 
.A(n_5159),
.Y(n_5688)
);

INVx2_ASAP7_75t_L g5689 ( 
.A(n_5174),
.Y(n_5689)
);

AOI21xp5_ASAP7_75t_L g5690 ( 
.A1(n_5029),
.A2(n_4640),
.B(n_4637),
.Y(n_5690)
);

INVx2_ASAP7_75t_L g5691 ( 
.A(n_5193),
.Y(n_5691)
);

NAND2xp5_ASAP7_75t_L g5692 ( 
.A(n_5179),
.B(n_4653),
.Y(n_5692)
);

AO22x1_ASAP7_75t_L g5693 ( 
.A1(n_5346),
.A2(n_1278),
.B1(n_1285),
.B2(n_1272),
.Y(n_5693)
);

AOI21xp5_ASAP7_75t_L g5694 ( 
.A1(n_5035),
.A2(n_4665),
.B(n_4659),
.Y(n_5694)
);

NOR2xp33_ASAP7_75t_L g5695 ( 
.A(n_4957),
.B(n_4828),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5193),
.Y(n_5696)
);

CKINVDCx5p33_ASAP7_75t_R g5697 ( 
.A(n_5159),
.Y(n_5697)
);

NAND2xp5_ASAP7_75t_L g5698 ( 
.A(n_5179),
.B(n_4659),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_5067),
.Y(n_5699)
);

HAxp5_ASAP7_75t_L g5700 ( 
.A(n_5202),
.B(n_1270),
.CON(n_5700),
.SN(n_5700)
);

OAI22xp5_ASAP7_75t_L g5701 ( 
.A1(n_4986),
.A2(n_5138),
.B1(n_5330),
.B2(n_5208),
.Y(n_5701)
);

AND2x2_ASAP7_75t_L g5702 ( 
.A(n_5028),
.B(n_4682),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_5295),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5342),
.Y(n_5704)
);

O2A1O1Ixp33_ASAP7_75t_L g5705 ( 
.A1(n_4985),
.A2(n_1286),
.B(n_1290),
.C(n_1278),
.Y(n_5705)
);

BUFx3_ASAP7_75t_L g5706 ( 
.A(n_5225),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_L g5707 ( 
.A(n_5028),
.B(n_4665),
.Y(n_5707)
);

NAND2xp5_ASAP7_75t_L g5708 ( 
.A(n_5343),
.B(n_4670),
.Y(n_5708)
);

OAI22xp5_ASAP7_75t_L g5709 ( 
.A1(n_5103),
.A2(n_4828),
.B1(n_4852),
.B2(n_4837),
.Y(n_5709)
);

BUFx8_ASAP7_75t_SL g5710 ( 
.A(n_5225),
.Y(n_5710)
);

INVx3_ASAP7_75t_L g5711 ( 
.A(n_5225),
.Y(n_5711)
);

NAND2xp5_ASAP7_75t_SL g5712 ( 
.A(n_5318),
.B(n_4670),
.Y(n_5712)
);

BUFx6f_ASAP7_75t_L g5713 ( 
.A(n_5243),
.Y(n_5713)
);

BUFx3_ASAP7_75t_L g5714 ( 
.A(n_5243),
.Y(n_5714)
);

OAI22xp5_ASAP7_75t_L g5715 ( 
.A1(n_5284),
.A2(n_4852),
.B1(n_4837),
.B2(n_4557),
.Y(n_5715)
);

AOI21xp5_ASAP7_75t_L g5716 ( 
.A1(n_5045),
.A2(n_4751),
.B(n_4749),
.Y(n_5716)
);

CKINVDCx8_ASAP7_75t_R g5717 ( 
.A(n_5049),
.Y(n_5717)
);

A2O1A1Ixp33_ASAP7_75t_SL g5718 ( 
.A1(n_4920),
.A2(n_1282),
.B(n_2354),
.C(n_2353),
.Y(n_5718)
);

OA21x2_ASAP7_75t_L g5719 ( 
.A1(n_5076),
.A2(n_4751),
.B(n_4749),
.Y(n_5719)
);

AND2x2_ASAP7_75t_L g5720 ( 
.A(n_5126),
.B(n_4682),
.Y(n_5720)
);

AOI21xp5_ASAP7_75t_L g5721 ( 
.A1(n_4963),
.A2(n_4771),
.B(n_4753),
.Y(n_5721)
);

INVx2_ASAP7_75t_SL g5722 ( 
.A(n_5243),
.Y(n_5722)
);

BUFx3_ASAP7_75t_L g5723 ( 
.A(n_5049),
.Y(n_5723)
);

AOI21xp5_ASAP7_75t_L g5724 ( 
.A1(n_5272),
.A2(n_4771),
.B(n_4753),
.Y(n_5724)
);

BUFx3_ASAP7_75t_L g5725 ( 
.A(n_5068),
.Y(n_5725)
);

AND2x2_ASAP7_75t_L g5726 ( 
.A(n_5126),
.B(n_4682),
.Y(n_5726)
);

A2O1A1Ixp33_ASAP7_75t_L g5727 ( 
.A1(n_5298),
.A2(n_4985),
.B(n_5026),
.C(n_5095),
.Y(n_5727)
);

OR2x6_ASAP7_75t_SL g5728 ( 
.A(n_5320),
.B(n_1086),
.Y(n_5728)
);

AND2x4_ASAP7_75t_L g5729 ( 
.A(n_5271),
.B(n_4683),
.Y(n_5729)
);

OR2x2_ASAP7_75t_L g5730 ( 
.A(n_5237),
.B(n_4778),
.Y(n_5730)
);

INVx2_ASAP7_75t_SL g5731 ( 
.A(n_5284),
.Y(n_5731)
);

INVx2_ASAP7_75t_SL g5732 ( 
.A(n_5344),
.Y(n_5732)
);

AOI21xp5_ASAP7_75t_L g5733 ( 
.A1(n_5245),
.A2(n_4782),
.B(n_4778),
.Y(n_5733)
);

AOI21xp5_ASAP7_75t_L g5734 ( 
.A1(n_5107),
.A2(n_4784),
.B(n_4782),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5352),
.Y(n_5735)
);

NAND2xp5_ASAP7_75t_L g5736 ( 
.A(n_5324),
.B(n_4784),
.Y(n_5736)
);

OAI22xp5_ASAP7_75t_L g5737 ( 
.A1(n_5344),
.A2(n_4558),
.B1(n_4573),
.B2(n_4514),
.Y(n_5737)
);

OAI21xp33_ASAP7_75t_L g5738 ( 
.A1(n_5326),
.A2(n_1286),
.B(n_1285),
.Y(n_5738)
);

OR2x2_ASAP7_75t_L g5739 ( 
.A(n_5204),
.B(n_4804),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5328),
.Y(n_5740)
);

OAI21x1_ASAP7_75t_L g5741 ( 
.A1(n_5195),
.A2(n_4814),
.B(n_4804),
.Y(n_5741)
);

AOI21xp5_ASAP7_75t_L g5742 ( 
.A1(n_5115),
.A2(n_4820),
.B(n_4814),
.Y(n_5742)
);

INVx3_ASAP7_75t_L g5743 ( 
.A(n_4962),
.Y(n_5743)
);

AOI22xp33_ASAP7_75t_L g5744 ( 
.A1(n_5315),
.A2(n_1282),
.B1(n_1296),
.B2(n_1290),
.Y(n_5744)
);

NOR3xp33_ASAP7_75t_L g5745 ( 
.A(n_4969),
.B(n_1296),
.C(n_1089),
.Y(n_5745)
);

NAND3xp33_ASAP7_75t_L g5746 ( 
.A(n_5027),
.B(n_1091),
.C(n_1088),
.Y(n_5746)
);

A2O1A1Ixp33_ASAP7_75t_SL g5747 ( 
.A1(n_4931),
.A2(n_5026),
.B(n_5298),
.C(n_4982),
.Y(n_5747)
);

AOI21xp5_ASAP7_75t_L g5748 ( 
.A1(n_5121),
.A2(n_4827),
.B(n_4820),
.Y(n_5748)
);

BUFx6f_ASAP7_75t_L g5749 ( 
.A(n_5068),
.Y(n_5749)
);

INVx2_ASAP7_75t_SL g5750 ( 
.A(n_4931),
.Y(n_5750)
);

OA22x2_ASAP7_75t_L g5751 ( 
.A1(n_5290),
.A2(n_4573),
.B1(n_4614),
.B2(n_4514),
.Y(n_5751)
);

AOI21xp5_ASAP7_75t_L g5752 ( 
.A1(n_5124),
.A2(n_5139),
.B(n_5131),
.Y(n_5752)
);

HB1xp67_ASAP7_75t_L g5753 ( 
.A(n_4982),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_5140),
.A2(n_4827),
.B(n_3351),
.Y(n_5754)
);

AOI21xp5_ASAP7_75t_L g5755 ( 
.A1(n_5105),
.A2(n_3351),
.B(n_3339),
.Y(n_5755)
);

BUFx6f_ASAP7_75t_L g5756 ( 
.A(n_5144),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5209),
.Y(n_5757)
);

OAI22xp5_ASAP7_75t_L g5758 ( 
.A1(n_5253),
.A2(n_4614),
.B1(n_4683),
.B2(n_1094),
.Y(n_5758)
);

NAND2xp5_ASAP7_75t_L g5759 ( 
.A(n_5150),
.B(n_4683),
.Y(n_5759)
);

OAI22xp5_ASAP7_75t_L g5760 ( 
.A1(n_5266),
.A2(n_4683),
.B1(n_1101),
.B2(n_1103),
.Y(n_5760)
);

OAI22xp5_ASAP7_75t_L g5761 ( 
.A1(n_5224),
.A2(n_1105),
.B1(n_1106),
.B2(n_1093),
.Y(n_5761)
);

OAI21x1_ASAP7_75t_L g5762 ( 
.A1(n_4954),
.A2(n_3354),
.B(n_3339),
.Y(n_5762)
);

AOI21xp5_ASAP7_75t_L g5763 ( 
.A1(n_5106),
.A2(n_3355),
.B(n_3354),
.Y(n_5763)
);

BUFx2_ASAP7_75t_L g5764 ( 
.A(n_4969),
.Y(n_5764)
);

NOR3xp33_ASAP7_75t_L g5765 ( 
.A(n_5022),
.B(n_1110),
.C(n_1107),
.Y(n_5765)
);

AND2x2_ASAP7_75t_L g5766 ( 
.A(n_5144),
.B(n_4683),
.Y(n_5766)
);

O2A1O1Ixp33_ASAP7_75t_SL g5767 ( 
.A1(n_5348),
.A2(n_1097),
.B(n_3505),
.C(n_3504),
.Y(n_5767)
);

OAI21xp5_ASAP7_75t_L g5768 ( 
.A1(n_5027),
.A2(n_3865),
.B(n_3848),
.Y(n_5768)
);

NAND2xp5_ASAP7_75t_L g5769 ( 
.A(n_5150),
.B(n_1111),
.Y(n_5769)
);

INVx4_ASAP7_75t_L g5770 ( 
.A(n_5022),
.Y(n_5770)
);

INVx3_ASAP7_75t_L g5771 ( 
.A(n_5295),
.Y(n_5771)
);

AOI21xp5_ASAP7_75t_L g5772 ( 
.A1(n_5166),
.A2(n_3356),
.B(n_3355),
.Y(n_5772)
);

NOR2xp33_ASAP7_75t_L g5773 ( 
.A(n_5187),
.B(n_1112),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5204),
.Y(n_5774)
);

NAND2xp5_ASAP7_75t_L g5775 ( 
.A(n_5172),
.B(n_1114),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5123),
.Y(n_5776)
);

O2A1O1Ixp5_ASAP7_75t_L g5777 ( 
.A1(n_5010),
.A2(n_3935),
.B(n_3943),
.C(n_3902),
.Y(n_5777)
);

BUFx2_ASAP7_75t_L g5778 ( 
.A(n_5187),
.Y(n_5778)
);

NAND2xp5_ASAP7_75t_L g5779 ( 
.A(n_5432),
.B(n_5156),
.Y(n_5779)
);

O2A1O1Ixp5_ASAP7_75t_L g5780 ( 
.A1(n_5404),
.A2(n_5327),
.B(n_5347),
.C(n_4992),
.Y(n_5780)
);

NAND2xp5_ASAP7_75t_L g5781 ( 
.A(n_5483),
.B(n_5172),
.Y(n_5781)
);

OAI21x1_ASAP7_75t_L g5782 ( 
.A1(n_5752),
.A2(n_5489),
.B(n_5576),
.Y(n_5782)
);

INVx8_ASAP7_75t_L g5783 ( 
.A(n_5564),
.Y(n_5783)
);

NAND2xp5_ASAP7_75t_L g5784 ( 
.A(n_5570),
.B(n_5122),
.Y(n_5784)
);

OAI21x1_ASAP7_75t_L g5785 ( 
.A1(n_5402),
.A2(n_5025),
.B(n_5087),
.Y(n_5785)
);

A2O1A1Ixp33_ASAP7_75t_L g5786 ( 
.A1(n_5555),
.A2(n_5475),
.B(n_5593),
.C(n_5580),
.Y(n_5786)
);

NAND2xp5_ASAP7_75t_L g5787 ( 
.A(n_5408),
.B(n_5133),
.Y(n_5787)
);

AOI21xp5_ASAP7_75t_L g5788 ( 
.A1(n_5394),
.A2(n_5127),
.B(n_5100),
.Y(n_5788)
);

AOI21xp5_ASAP7_75t_SL g5789 ( 
.A1(n_5389),
.A2(n_5353),
.B(n_5230),
.Y(n_5789)
);

CKINVDCx5p33_ASAP7_75t_R g5790 ( 
.A(n_5377),
.Y(n_5790)
);

AO22x2_ASAP7_75t_L g5791 ( 
.A1(n_5774),
.A2(n_5224),
.B1(n_5297),
.B2(n_5214),
.Y(n_5791)
);

AOI21xp5_ASAP7_75t_L g5792 ( 
.A1(n_5374),
.A2(n_5244),
.B(n_5220),
.Y(n_5792)
);

NAND2xp5_ASAP7_75t_L g5793 ( 
.A(n_5462),
.B(n_5297),
.Y(n_5793)
);

AO31x2_ASAP7_75t_L g5794 ( 
.A1(n_5369),
.A2(n_5192),
.A3(n_5196),
.B(n_5188),
.Y(n_5794)
);

INVx2_ASAP7_75t_L g5795 ( 
.A(n_5513),
.Y(n_5795)
);

OAI21x1_ASAP7_75t_L g5796 ( 
.A1(n_5661),
.A2(n_5255),
.B(n_5207),
.Y(n_5796)
);

OAI21x1_ASAP7_75t_SL g5797 ( 
.A1(n_5363),
.A2(n_5226),
.B(n_5218),
.Y(n_5797)
);

HB1xp67_ASAP7_75t_L g5798 ( 
.A(n_5379),
.Y(n_5798)
);

OAI21x1_ASAP7_75t_L g5799 ( 
.A1(n_5505),
.A2(n_5206),
.B(n_5334),
.Y(n_5799)
);

NAND2xp5_ASAP7_75t_L g5800 ( 
.A(n_5383),
.B(n_5214),
.Y(n_5800)
);

NAND2xp5_ASAP7_75t_L g5801 ( 
.A(n_5364),
.B(n_5213),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5356),
.Y(n_5802)
);

AOI221xp5_ASAP7_75t_SL g5803 ( 
.A1(n_5453),
.A2(n_976),
.B1(n_1158),
.B2(n_902),
.C(n_850),
.Y(n_5803)
);

OAI21x1_ASAP7_75t_L g5804 ( 
.A1(n_5373),
.A2(n_5299),
.B(n_5294),
.Y(n_5804)
);

AOI21xp5_ASAP7_75t_L g5805 ( 
.A1(n_5391),
.A2(n_5241),
.B(n_5307),
.Y(n_5805)
);

NAND2xp5_ASAP7_75t_L g5806 ( 
.A(n_5422),
.B(n_5215),
.Y(n_5806)
);

OAI21xp33_ASAP7_75t_SL g5807 ( 
.A1(n_5604),
.A2(n_5246),
.B(n_5316),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5368),
.Y(n_5808)
);

INVx6_ASAP7_75t_L g5809 ( 
.A(n_5409),
.Y(n_5809)
);

NAND3xp33_ASAP7_75t_L g5810 ( 
.A(n_5746),
.B(n_1122),
.C(n_1118),
.Y(n_5810)
);

AO31x2_ASAP7_75t_L g5811 ( 
.A1(n_5684),
.A2(n_5325),
.A3(n_5341),
.B(n_5322),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_5628),
.A2(n_5191),
.B(n_5184),
.Y(n_5812)
);

OAI21x1_ASAP7_75t_L g5813 ( 
.A1(n_5640),
.A2(n_5205),
.B(n_5203),
.Y(n_5813)
);

BUFx6f_ASAP7_75t_L g5814 ( 
.A(n_5526),
.Y(n_5814)
);

OAI21xp5_ASAP7_75t_L g5815 ( 
.A1(n_5746),
.A2(n_5186),
.B(n_5148),
.Y(n_5815)
);

AOI21xp5_ASAP7_75t_L g5816 ( 
.A1(n_5371),
.A2(n_5246),
.B(n_5186),
.Y(n_5816)
);

NAND2xp5_ASAP7_75t_SL g5817 ( 
.A(n_5517),
.B(n_5148),
.Y(n_5817)
);

AND2x4_ASAP7_75t_L g5818 ( 
.A(n_5520),
.B(n_5689),
.Y(n_5818)
);

OAI21x1_ASAP7_75t_L g5819 ( 
.A1(n_5639),
.A2(n_5550),
.B(n_5469),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_SL g5820 ( 
.A(n_5517),
.B(n_1582),
.Y(n_5820)
);

AOI21xp5_ASAP7_75t_L g5821 ( 
.A1(n_5371),
.A2(n_5246),
.B(n_3278),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5380),
.Y(n_5822)
);

NAND2x1_ASAP7_75t_L g5823 ( 
.A(n_5370),
.B(n_3865),
.Y(n_5823)
);

AOI21xp5_ASAP7_75t_L g5824 ( 
.A1(n_5448),
.A2(n_3229),
.B(n_3226),
.Y(n_5824)
);

OAI21x1_ASAP7_75t_L g5825 ( 
.A1(n_5381),
.A2(n_3358),
.B(n_3356),
.Y(n_5825)
);

OAI21x1_ASAP7_75t_L g5826 ( 
.A1(n_5527),
.A2(n_3358),
.B(n_3935),
.Y(n_5826)
);

NAND2xp5_ASAP7_75t_L g5827 ( 
.A(n_5388),
.B(n_1678),
.Y(n_5827)
);

INVx1_ASAP7_75t_SL g5828 ( 
.A(n_5585),
.Y(n_5828)
);

INVx3_ASAP7_75t_L g5829 ( 
.A(n_5386),
.Y(n_5829)
);

NAND2xp5_ASAP7_75t_L g5830 ( 
.A(n_5401),
.B(n_1678),
.Y(n_5830)
);

AOI31xp67_ASAP7_75t_L g5831 ( 
.A1(n_5751),
.A2(n_2358),
.A3(n_2361),
.B(n_2354),
.Y(n_5831)
);

AOI31xp67_ASAP7_75t_L g5832 ( 
.A1(n_5425),
.A2(n_2361),
.A3(n_2362),
.B(n_2358),
.Y(n_5832)
);

NAND2xp5_ASAP7_75t_L g5833 ( 
.A(n_5567),
.B(n_1678),
.Y(n_5833)
);

A2O1A1Ixp33_ASAP7_75t_L g5834 ( 
.A1(n_5586),
.A2(n_1157),
.B(n_1171),
.C(n_1138),
.Y(n_5834)
);

AOI21xp5_ASAP7_75t_L g5835 ( 
.A1(n_5395),
.A2(n_5442),
.B(n_5441),
.Y(n_5835)
);

NOR2xp33_ASAP7_75t_L g5836 ( 
.A(n_5562),
.B(n_1582),
.Y(n_5836)
);

OAI21x1_ASAP7_75t_L g5837 ( 
.A1(n_5565),
.A2(n_3949),
.B(n_3943),
.Y(n_5837)
);

AOI21xp5_ASAP7_75t_L g5838 ( 
.A1(n_5439),
.A2(n_3229),
.B(n_3226),
.Y(n_5838)
);

OAI21x1_ASAP7_75t_L g5839 ( 
.A1(n_5613),
.A2(n_3961),
.B(n_3949),
.Y(n_5839)
);

AOI221x1_ASAP7_75t_L g5840 ( 
.A1(n_5646),
.A2(n_1638),
.B1(n_1758),
.B2(n_1626),
.C(n_1586),
.Y(n_5840)
);

BUFx12f_ASAP7_75t_L g5841 ( 
.A(n_5378),
.Y(n_5841)
);

OAI21x1_ASAP7_75t_L g5842 ( 
.A1(n_5511),
.A2(n_3986),
.B(n_3961),
.Y(n_5842)
);

INVx2_ASAP7_75t_SL g5843 ( 
.A(n_5526),
.Y(n_5843)
);

AO32x2_ASAP7_75t_L g5844 ( 
.A1(n_5522),
.A2(n_1191),
.A3(n_1195),
.B1(n_1158),
.B2(n_850),
.Y(n_5844)
);

OAI21x1_ASAP7_75t_L g5845 ( 
.A1(n_5569),
.A2(n_3988),
.B(n_3986),
.Y(n_5845)
);

AO21x1_ASAP7_75t_L g5846 ( 
.A1(n_5554),
.A2(n_1191),
.B(n_1158),
.Y(n_5846)
);

INVx2_ASAP7_75t_L g5847 ( 
.A(n_5521),
.Y(n_5847)
);

OAI21x1_ASAP7_75t_L g5848 ( 
.A1(n_5466),
.A2(n_4002),
.B(n_3988),
.Y(n_5848)
);

O2A1O1Ixp5_ASAP7_75t_SL g5849 ( 
.A1(n_5757),
.A2(n_4032),
.B(n_4010),
.C(n_4002),
.Y(n_5849)
);

INVx6_ASAP7_75t_L g5850 ( 
.A(n_5409),
.Y(n_5850)
);

OAI21xp5_ASAP7_75t_L g5851 ( 
.A1(n_5775),
.A2(n_3865),
.B(n_1128),
.Y(n_5851)
);

AOI221x1_ASAP7_75t_L g5852 ( 
.A1(n_5516),
.A2(n_1638),
.B1(n_1758),
.B2(n_1626),
.C(n_1586),
.Y(n_5852)
);

NAND2xp5_ASAP7_75t_L g5853 ( 
.A(n_5502),
.B(n_1586),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_5424),
.B(n_1586),
.Y(n_5854)
);

AOI221x1_ASAP7_75t_L g5855 ( 
.A1(n_5453),
.A2(n_5455),
.B1(n_5534),
.B2(n_5667),
.C(n_5644),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_L g5856 ( 
.A(n_5592),
.B(n_1586),
.Y(n_5856)
);

OAI21xp5_ASAP7_75t_L g5857 ( 
.A1(n_5631),
.A2(n_5769),
.B(n_5705),
.Y(n_5857)
);

AOI21xp5_ASAP7_75t_L g5858 ( 
.A1(n_5403),
.A2(n_3238),
.B(n_3234),
.Y(n_5858)
);

AO31x2_ASAP7_75t_L g5859 ( 
.A1(n_5776),
.A2(n_3238),
.A3(n_3242),
.B(n_3234),
.Y(n_5859)
);

OAI21x1_ASAP7_75t_L g5860 ( 
.A1(n_5493),
.A2(n_5583),
.B(n_5762),
.Y(n_5860)
);

INVx2_ASAP7_75t_SL g5861 ( 
.A(n_5526),
.Y(n_5861)
);

OAI21xp5_ASAP7_75t_L g5862 ( 
.A1(n_5745),
.A2(n_1132),
.B(n_1127),
.Y(n_5862)
);

NAND2xp5_ASAP7_75t_L g5863 ( 
.A(n_5440),
.B(n_1626),
.Y(n_5863)
);

AOI21xp5_ASAP7_75t_SL g5864 ( 
.A1(n_5385),
.A2(n_3975),
.B(n_3969),
.Y(n_5864)
);

OAI21x1_ASAP7_75t_SL g5865 ( 
.A1(n_5701),
.A2(n_2368),
.B(n_2362),
.Y(n_5865)
);

OR2x2_ASAP7_75t_L g5866 ( 
.A(n_5484),
.B(n_1626),
.Y(n_5866)
);

NAND2xp5_ASAP7_75t_L g5867 ( 
.A(n_5479),
.B(n_1626),
.Y(n_5867)
);

OAI21xp5_ASAP7_75t_L g5868 ( 
.A1(n_5459),
.A2(n_1134),
.B(n_1133),
.Y(n_5868)
);

AOI21xp5_ASAP7_75t_L g5869 ( 
.A1(n_5436),
.A2(n_3245),
.B(n_3242),
.Y(n_5869)
);

OAI21x1_ASAP7_75t_L g5870 ( 
.A1(n_5633),
.A2(n_4032),
.B(n_4010),
.Y(n_5870)
);

INVx2_ASAP7_75t_L g5871 ( 
.A(n_5536),
.Y(n_5871)
);

OAI21xp5_ASAP7_75t_L g5872 ( 
.A1(n_5434),
.A2(n_1141),
.B(n_1140),
.Y(n_5872)
);

OAI21x1_ASAP7_75t_L g5873 ( 
.A1(n_5392),
.A2(n_3248),
.B(n_3245),
.Y(n_5873)
);

NAND2xp5_ASAP7_75t_L g5874 ( 
.A(n_5494),
.B(n_1638),
.Y(n_5874)
);

OAI21xp5_ASAP7_75t_L g5875 ( 
.A1(n_5497),
.A2(n_1145),
.B(n_1142),
.Y(n_5875)
);

NAND2xp5_ASAP7_75t_L g5876 ( 
.A(n_5496),
.B(n_1638),
.Y(n_5876)
);

AND2x2_ASAP7_75t_L g5877 ( 
.A(n_5365),
.B(n_1638),
.Y(n_5877)
);

OAI21xp5_ASAP7_75t_L g5878 ( 
.A1(n_5497),
.A2(n_1150),
.B(n_1149),
.Y(n_5878)
);

NAND2xp5_ASAP7_75t_L g5879 ( 
.A(n_5445),
.B(n_5430),
.Y(n_5879)
);

OAI21x1_ASAP7_75t_L g5880 ( 
.A1(n_5392),
.A2(n_3248),
.B(n_3487),
.Y(n_5880)
);

AO31x2_ASAP7_75t_L g5881 ( 
.A1(n_5740),
.A2(n_3520),
.A3(n_3522),
.B(n_3508),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_L g5882 ( 
.A(n_5692),
.B(n_1758),
.Y(n_5882)
);

AO31x2_ASAP7_75t_L g5883 ( 
.A1(n_5704),
.A2(n_5735),
.A3(n_5727),
.B(n_5616),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_5698),
.B(n_1758),
.Y(n_5884)
);

BUFx3_ASAP7_75t_L g5885 ( 
.A(n_5531),
.Y(n_5885)
);

NAND2xp5_ASAP7_75t_L g5886 ( 
.A(n_5699),
.B(n_1758),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5578),
.Y(n_5887)
);

OAI21x1_ASAP7_75t_L g5888 ( 
.A1(n_5621),
.A2(n_3488),
.B(n_3487),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_L g5889 ( 
.A(n_5753),
.B(n_1154),
.Y(n_5889)
);

INVx2_ASAP7_75t_L g5890 ( 
.A(n_5528),
.Y(n_5890)
);

OAI21x1_ASAP7_75t_L g5891 ( 
.A1(n_5626),
.A2(n_3488),
.B(n_3487),
.Y(n_5891)
);

OAI21x1_ASAP7_75t_L g5892 ( 
.A1(n_5601),
.A2(n_3502),
.B(n_3488),
.Y(n_5892)
);

NAND2xp5_ASAP7_75t_L g5893 ( 
.A(n_5707),
.B(n_1160),
.Y(n_5893)
);

OAI21x1_ASAP7_75t_L g5894 ( 
.A1(n_5754),
.A2(n_3502),
.B(n_3488),
.Y(n_5894)
);

HB1xp67_ASAP7_75t_L g5895 ( 
.A(n_5627),
.Y(n_5895)
);

AOI21xp5_ASAP7_75t_L g5896 ( 
.A1(n_5444),
.A2(n_2935),
.B(n_3796),
.Y(n_5896)
);

AOI221x1_ASAP7_75t_L g5897 ( 
.A1(n_5455),
.A2(n_5416),
.B1(n_5678),
.B2(n_5465),
.C(n_5387),
.Y(n_5897)
);

INVx2_ASAP7_75t_SL g5898 ( 
.A(n_5531),
.Y(n_5898)
);

NAND2xp5_ASAP7_75t_SL g5899 ( 
.A(n_5517),
.B(n_1489),
.Y(n_5899)
);

OAI21x1_ASAP7_75t_L g5900 ( 
.A1(n_5637),
.A2(n_3540),
.B(n_3502),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5634),
.B(n_1158),
.Y(n_5901)
);

OR2x2_ASAP7_75t_L g5902 ( 
.A(n_5357),
.B(n_7),
.Y(n_5902)
);

INVx4_ASAP7_75t_L g5903 ( 
.A(n_5411),
.Y(n_5903)
);

AND2x2_ASAP7_75t_L g5904 ( 
.A(n_5540),
.B(n_5607),
.Y(n_5904)
);

NAND2xp5_ASAP7_75t_L g5905 ( 
.A(n_5573),
.B(n_1163),
.Y(n_5905)
);

NOR2xp33_ASAP7_75t_L g5906 ( 
.A(n_5619),
.B(n_1165),
.Y(n_5906)
);

NAND2xp5_ASAP7_75t_L g5907 ( 
.A(n_5683),
.B(n_1166),
.Y(n_5907)
);

INVx3_ASAP7_75t_L g5908 ( 
.A(n_5421),
.Y(n_5908)
);

INVx2_ASAP7_75t_L g5909 ( 
.A(n_5544),
.Y(n_5909)
);

OAI21x1_ASAP7_75t_L g5910 ( 
.A1(n_5490),
.A2(n_3540),
.B(n_3502),
.Y(n_5910)
);

AOI22x1_ASAP7_75t_L g5911 ( 
.A1(n_5595),
.A2(n_1167),
.B1(n_1172),
.B2(n_1170),
.Y(n_5911)
);

OAI21x1_ASAP7_75t_L g5912 ( 
.A1(n_5716),
.A2(n_3565),
.B(n_3540),
.Y(n_5912)
);

OAI21x1_ASAP7_75t_L g5913 ( 
.A1(n_5777),
.A2(n_3565),
.B(n_3540),
.Y(n_5913)
);

AO221x2_ASAP7_75t_L g5914 ( 
.A1(n_5359),
.A2(n_12),
.B1(n_8),
.B2(n_10),
.C(n_13),
.Y(n_5914)
);

OAI21x1_ASAP7_75t_L g5915 ( 
.A1(n_5685),
.A2(n_5694),
.B(n_5690),
.Y(n_5915)
);

NAND2xp5_ASAP7_75t_L g5916 ( 
.A(n_5638),
.B(n_1174),
.Y(n_5916)
);

OAI21x1_ASAP7_75t_L g5917 ( 
.A1(n_5506),
.A2(n_3597),
.B(n_3565),
.Y(n_5917)
);

NAND2xp5_ASAP7_75t_L g5918 ( 
.A(n_5431),
.B(n_1175),
.Y(n_5918)
);

INVx2_ASAP7_75t_L g5919 ( 
.A(n_5400),
.Y(n_5919)
);

OAI21x1_ASAP7_75t_L g5920 ( 
.A1(n_5446),
.A2(n_3597),
.B(n_3565),
.Y(n_5920)
);

AOI21xp5_ASAP7_75t_L g5921 ( 
.A1(n_5500),
.A2(n_3821),
.B(n_3796),
.Y(n_5921)
);

OAI21xp5_ASAP7_75t_L g5922 ( 
.A1(n_5467),
.A2(n_1183),
.B(n_1180),
.Y(n_5922)
);

OAI22x1_ASAP7_75t_L g5923 ( 
.A1(n_5530),
.A2(n_1189),
.B1(n_1192),
.B2(n_1188),
.Y(n_5923)
);

A2O1A1Ixp33_ASAP7_75t_L g5924 ( 
.A1(n_5457),
.A2(n_1220),
.B(n_1236),
.C(n_1202),
.Y(n_5924)
);

OAI21x1_ASAP7_75t_SL g5925 ( 
.A1(n_5677),
.A2(n_2373),
.B(n_2368),
.Y(n_5925)
);

NAND2xp5_ASAP7_75t_L g5926 ( 
.A(n_5568),
.B(n_1193),
.Y(n_5926)
);

AOI21xp5_ASAP7_75t_L g5927 ( 
.A1(n_5456),
.A2(n_3821),
.B(n_3796),
.Y(n_5927)
);

NAND2xp5_ASAP7_75t_L g5928 ( 
.A(n_5558),
.B(n_5525),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_L g5929 ( 
.A(n_5557),
.B(n_1194),
.Y(n_5929)
);

OR2x6_ASAP7_75t_L g5930 ( 
.A(n_5360),
.B(n_3975),
.Y(n_5930)
);

NAND2xp5_ASAP7_75t_L g5931 ( 
.A(n_5437),
.B(n_5556),
.Y(n_5931)
);

INVx4_ASAP7_75t_L g5932 ( 
.A(n_5411),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5435),
.Y(n_5933)
);

NOR2xp33_ASAP7_75t_SL g5934 ( 
.A(n_5575),
.B(n_3697),
.Y(n_5934)
);

OAI21xp5_ASAP7_75t_L g5935 ( 
.A1(n_5481),
.A2(n_1197),
.B(n_1196),
.Y(n_5935)
);

NAND2xp33_ASAP7_75t_L g5936 ( 
.A(n_5679),
.B(n_1199),
.Y(n_5936)
);

AOI22xp5_ASAP7_75t_L g5937 ( 
.A1(n_5418),
.A2(n_1204),
.B1(n_1207),
.B2(n_1200),
.Y(n_5937)
);

CKINVDCx14_ASAP7_75t_R g5938 ( 
.A(n_5450),
.Y(n_5938)
);

BUFx6f_ASAP7_75t_L g5939 ( 
.A(n_5531),
.Y(n_5939)
);

AOI21x1_ASAP7_75t_SL g5940 ( 
.A1(n_5729),
.A2(n_1097),
.B(n_8),
.Y(n_5940)
);

INVx4_ASAP7_75t_L g5941 ( 
.A(n_5535),
.Y(n_5941)
);

OAI21xp5_ASAP7_75t_L g5942 ( 
.A1(n_5529),
.A2(n_1212),
.B(n_1209),
.Y(n_5942)
);

CKINVDCx5p33_ASAP7_75t_R g5943 ( 
.A(n_5566),
.Y(n_5943)
);

AOI21xp5_ASAP7_75t_L g5944 ( 
.A1(n_5405),
.A2(n_3930),
.B(n_3821),
.Y(n_5944)
);

NOR2x1_ASAP7_75t_L g5945 ( 
.A(n_5618),
.B(n_3975),
.Y(n_5945)
);

AOI21x1_ASAP7_75t_L g5946 ( 
.A1(n_5693),
.A2(n_2375),
.B(n_2373),
.Y(n_5946)
);

CKINVDCx14_ASAP7_75t_R g5947 ( 
.A(n_5587),
.Y(n_5947)
);

OAI21xp5_ASAP7_75t_SL g5948 ( 
.A1(n_5433),
.A2(n_1195),
.B(n_1191),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5560),
.B(n_1213),
.Y(n_5949)
);

AOI21xp5_ASAP7_75t_L g5950 ( 
.A1(n_5420),
.A2(n_4047),
.B(n_3930),
.Y(n_5950)
);

AND2x2_ASAP7_75t_SL g5951 ( 
.A(n_5507),
.B(n_3981),
.Y(n_5951)
);

INVx2_ASAP7_75t_L g5952 ( 
.A(n_5452),
.Y(n_5952)
);

NOR2xp67_ASAP7_75t_L g5953 ( 
.A(n_5618),
.B(n_5454),
.Y(n_5953)
);

NOR2xp33_ASAP7_75t_L g5954 ( 
.A(n_5649),
.B(n_1215),
.Y(n_5954)
);

AOI221x1_ASAP7_75t_L g5955 ( 
.A1(n_5582),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.C(n_15),
.Y(n_5955)
);

OAI21x1_ASAP7_75t_L g5956 ( 
.A1(n_5451),
.A2(n_3605),
.B(n_3597),
.Y(n_5956)
);

OAI21x1_ASAP7_75t_L g5957 ( 
.A1(n_5426),
.A2(n_3605),
.B(n_3597),
.Y(n_5957)
);

OAI21x1_ASAP7_75t_L g5958 ( 
.A1(n_5768),
.A2(n_3605),
.B(n_3468),
.Y(n_5958)
);

OA21x2_ASAP7_75t_L g5959 ( 
.A1(n_5674),
.A2(n_1221),
.B(n_1219),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_L g5960 ( 
.A(n_5518),
.B(n_1222),
.Y(n_5960)
);

OAI21xp5_ASAP7_75t_L g5961 ( 
.A1(n_5577),
.A2(n_1228),
.B(n_1227),
.Y(n_5961)
);

OAI21xp5_ASAP7_75t_L g5962 ( 
.A1(n_5447),
.A2(n_1233),
.B(n_1229),
.Y(n_5962)
);

AOI21xp33_ASAP7_75t_L g5963 ( 
.A1(n_5747),
.A2(n_1244),
.B(n_1235),
.Y(n_5963)
);

OAI21x1_ASAP7_75t_L g5964 ( 
.A1(n_5768),
.A2(n_3605),
.B(n_3468),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5460),
.Y(n_5965)
);

AND2x4_ASAP7_75t_L g5966 ( 
.A(n_5520),
.B(n_3930),
.Y(n_5966)
);

AND2x2_ASAP7_75t_L g5967 ( 
.A(n_5625),
.B(n_1191),
.Y(n_5967)
);

NAND2xp5_ASAP7_75t_L g5968 ( 
.A(n_5650),
.B(n_1246),
.Y(n_5968)
);

OAI21xp33_ASAP7_75t_L g5969 ( 
.A1(n_5433),
.A2(n_1249),
.B(n_1248),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5461),
.Y(n_5970)
);

OAI21x1_ASAP7_75t_L g5971 ( 
.A1(n_5734),
.A2(n_3468),
.B(n_3464),
.Y(n_5971)
);

INVx2_ASAP7_75t_SL g5972 ( 
.A(n_5535),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5366),
.B(n_5548),
.Y(n_5973)
);

AND2x2_ASAP7_75t_L g5974 ( 
.A(n_5662),
.B(n_1195),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_5664),
.B(n_5642),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_SL g5976 ( 
.A(n_5535),
.B(n_1489),
.Y(n_5976)
);

OAI21x1_ASAP7_75t_L g5977 ( 
.A1(n_5742),
.A2(n_3474),
.B(n_3464),
.Y(n_5977)
);

OAI21xp5_ASAP7_75t_L g5978 ( 
.A1(n_5598),
.A2(n_1252),
.B(n_1251),
.Y(n_5978)
);

OAI21xp5_ASAP7_75t_L g5979 ( 
.A1(n_5414),
.A2(n_5542),
.B(n_5355),
.Y(n_5979)
);

INVx6_ASAP7_75t_L g5980 ( 
.A(n_5378),
.Y(n_5980)
);

INVxp67_ASAP7_75t_SL g5981 ( 
.A(n_5508),
.Y(n_5981)
);

AOI21x1_ASAP7_75t_SL g5982 ( 
.A1(n_5729),
.A2(n_5759),
.B(n_5538),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5468),
.Y(n_5983)
);

BUFx6f_ASAP7_75t_L g5984 ( 
.A(n_5410),
.Y(n_5984)
);

AND2x4_ASAP7_75t_L g5985 ( 
.A(n_5591),
.B(n_4047),
.Y(n_5985)
);

NAND2xp5_ASAP7_75t_L g5986 ( 
.A(n_5702),
.B(n_1253),
.Y(n_5986)
);

AO31x2_ASAP7_75t_L g5987 ( 
.A1(n_5652),
.A2(n_3522),
.A3(n_3523),
.B(n_3520),
.Y(n_5987)
);

INVx2_ASAP7_75t_L g5988 ( 
.A(n_5478),
.Y(n_5988)
);

AOI21xp5_ASAP7_75t_L g5989 ( 
.A1(n_5654),
.A2(n_3528),
.B(n_3523),
.Y(n_5989)
);

A2O1A1Ixp33_ASAP7_75t_L g5990 ( 
.A1(n_5423),
.A2(n_1289),
.B(n_1260),
.C(n_1258),
.Y(n_5990)
);

INVx2_ASAP7_75t_L g5991 ( 
.A(n_5480),
.Y(n_5991)
);

A2O1A1Ixp33_ASAP7_75t_L g5992 ( 
.A1(n_5384),
.A2(n_1276),
.B(n_1295),
.C(n_1263),
.Y(n_5992)
);

OAI21x1_ASAP7_75t_L g5993 ( 
.A1(n_5748),
.A2(n_3474),
.B(n_3464),
.Y(n_5993)
);

NOR2xp33_ASAP7_75t_SL g5994 ( 
.A(n_5602),
.B(n_3697),
.Y(n_5994)
);

OAI21x1_ASAP7_75t_L g5995 ( 
.A1(n_5772),
.A2(n_3475),
.B(n_3474),
.Y(n_5995)
);

AO31x2_ASAP7_75t_L g5996 ( 
.A1(n_5672),
.A2(n_3529),
.A3(n_3531),
.B(n_3528),
.Y(n_5996)
);

OAI21x1_ASAP7_75t_SL g5997 ( 
.A1(n_5375),
.A2(n_2384),
.B(n_2375),
.Y(n_5997)
);

NAND2xp5_ASAP7_75t_L g5998 ( 
.A(n_5632),
.B(n_5641),
.Y(n_5998)
);

OAI21x1_ASAP7_75t_L g5999 ( 
.A1(n_5503),
.A2(n_3482),
.B(n_3475),
.Y(n_5999)
);

NAND2xp5_ASAP7_75t_L g6000 ( 
.A(n_5641),
.B(n_1254),
.Y(n_6000)
);

OAI21xp5_ASAP7_75t_L g6001 ( 
.A1(n_5477),
.A2(n_1264),
.B(n_1261),
.Y(n_6001)
);

OAI21x1_ASAP7_75t_L g6002 ( 
.A1(n_5660),
.A2(n_3482),
.B(n_3475),
.Y(n_6002)
);

OAI21xp5_ASAP7_75t_L g6003 ( 
.A1(n_5765),
.A2(n_1266),
.B(n_1265),
.Y(n_6003)
);

AOI21xp5_ASAP7_75t_L g6004 ( 
.A1(n_5501),
.A2(n_3531),
.B(n_3529),
.Y(n_6004)
);

INVx3_ASAP7_75t_L g6005 ( 
.A(n_5421),
.Y(n_6005)
);

OAI21x1_ASAP7_75t_L g6006 ( 
.A1(n_5721),
.A2(n_3484),
.B(n_3482),
.Y(n_6006)
);

AO31x2_ASAP7_75t_L g6007 ( 
.A1(n_5673),
.A2(n_3549),
.A3(n_3553),
.B(n_3547),
.Y(n_6007)
);

OA21x2_ASAP7_75t_L g6008 ( 
.A1(n_5653),
.A2(n_1269),
.B(n_1268),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_5648),
.B(n_1273),
.Y(n_6009)
);

INVx2_ASAP7_75t_L g6010 ( 
.A(n_5509),
.Y(n_6010)
);

AOI21xp5_ASAP7_75t_L g6011 ( 
.A1(n_5427),
.A2(n_3549),
.B(n_3547),
.Y(n_6011)
);

OA21x2_ASAP7_75t_L g6012 ( 
.A1(n_5733),
.A2(n_1280),
.B(n_1277),
.Y(n_6012)
);

NAND2xp5_ASAP7_75t_L g6013 ( 
.A(n_5648),
.B(n_1284),
.Y(n_6013)
);

NAND3xp33_ASAP7_75t_L g6014 ( 
.A(n_5463),
.B(n_1288),
.C(n_1287),
.Y(n_6014)
);

OAI21xp5_ASAP7_75t_L g6015 ( 
.A1(n_5659),
.A2(n_1294),
.B(n_1292),
.Y(n_6015)
);

A2O1A1Ixp33_ASAP7_75t_L g6016 ( 
.A1(n_5510),
.A2(n_1300),
.B(n_1297),
.C(n_1240),
.Y(n_6016)
);

OR2x2_ASAP7_75t_L g6017 ( 
.A(n_5406),
.B(n_15),
.Y(n_6017)
);

NAND3xp33_ASAP7_75t_L g6018 ( 
.A(n_5596),
.B(n_2390),
.C(n_2384),
.Y(n_6018)
);

AND2x2_ASAP7_75t_L g6019 ( 
.A(n_5608),
.B(n_5615),
.Y(n_6019)
);

INVx3_ASAP7_75t_L g6020 ( 
.A(n_5410),
.Y(n_6020)
);

OAI21x1_ASAP7_75t_L g6021 ( 
.A1(n_5476),
.A2(n_3484),
.B(n_3553),
.Y(n_6021)
);

NOR2xp33_ASAP7_75t_L g6022 ( 
.A(n_5728),
.B(n_17),
.Y(n_6022)
);

BUFx6f_ASAP7_75t_L g6023 ( 
.A(n_5410),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_5589),
.B(n_18),
.Y(n_6024)
);

NAND2xp5_ASAP7_75t_L g6025 ( 
.A(n_5590),
.B(n_19),
.Y(n_6025)
);

OAI21xp5_ASAP7_75t_L g6026 ( 
.A1(n_5398),
.A2(n_2414),
.B(n_2390),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_5512),
.Y(n_6027)
);

NAND2xp5_ASAP7_75t_L g6028 ( 
.A(n_5599),
.B(n_20),
.Y(n_6028)
);

AOI21x1_ASAP7_75t_L g6029 ( 
.A1(n_5488),
.A2(n_2420),
.B(n_2414),
.Y(n_6029)
);

NAND2xp5_ASAP7_75t_L g6030 ( 
.A(n_5629),
.B(n_5636),
.Y(n_6030)
);

OAI21xp5_ASAP7_75t_L g6031 ( 
.A1(n_5412),
.A2(n_2420),
.B(n_3816),
.Y(n_6031)
);

AND2x2_ASAP7_75t_L g6032 ( 
.A(n_5778),
.B(n_1195),
.Y(n_6032)
);

OAI21x1_ASAP7_75t_L g6033 ( 
.A1(n_5755),
.A2(n_3484),
.B(n_3556),
.Y(n_6033)
);

NOR2xp33_ASAP7_75t_L g6034 ( 
.A(n_5514),
.B(n_21),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_5720),
.B(n_22),
.Y(n_6035)
);

NAND2xp5_ASAP7_75t_L g6036 ( 
.A(n_5726),
.B(n_23),
.Y(n_6036)
);

NAND2xp5_ASAP7_75t_L g6037 ( 
.A(n_5610),
.B(n_25),
.Y(n_6037)
);

NOR2x1_ASAP7_75t_SL g6038 ( 
.A(n_5591),
.B(n_3981),
.Y(n_6038)
);

OAI21x1_ASAP7_75t_L g6039 ( 
.A1(n_5763),
.A2(n_3564),
.B(n_3556),
.Y(n_6039)
);

AO32x2_ASAP7_75t_L g6040 ( 
.A1(n_5522),
.A2(n_1270),
.A3(n_1242),
.B1(n_1240),
.B2(n_1489),
.Y(n_6040)
);

BUFx6f_ASAP7_75t_L g6041 ( 
.A(n_5606),
.Y(n_6041)
);

NAND2xp5_ASAP7_75t_L g6042 ( 
.A(n_5361),
.B(n_5362),
.Y(n_6042)
);

NAND2xp5_ASAP7_75t_L g6043 ( 
.A(n_5367),
.B(n_25),
.Y(n_6043)
);

INVx3_ASAP7_75t_L g6044 ( 
.A(n_5443),
.Y(n_6044)
);

O2A1O1Ixp33_ASAP7_75t_L g6045 ( 
.A1(n_5623),
.A2(n_1242),
.B(n_1270),
.C(n_1240),
.Y(n_6045)
);

AO21x1_ASAP7_75t_L g6046 ( 
.A1(n_5571),
.A2(n_1242),
.B(n_1240),
.Y(n_6046)
);

AND2x4_ASAP7_75t_L g6047 ( 
.A(n_5591),
.B(n_3990),
.Y(n_6047)
);

NAND2xp5_ASAP7_75t_L g6048 ( 
.A(n_5382),
.B(n_26),
.Y(n_6048)
);

OAI21x1_ASAP7_75t_SL g6049 ( 
.A1(n_5486),
.A2(n_3571),
.B(n_3564),
.Y(n_6049)
);

BUFx10_ASAP7_75t_L g6050 ( 
.A(n_5773),
.Y(n_6050)
);

BUFx3_ASAP7_75t_L g6051 ( 
.A(n_5552),
.Y(n_6051)
);

AO31x2_ASAP7_75t_L g6052 ( 
.A1(n_5485),
.A2(n_3573),
.A3(n_3571),
.B(n_3322),
.Y(n_6052)
);

OAI21x1_ASAP7_75t_SL g6053 ( 
.A1(n_5658),
.A2(n_3573),
.B(n_3322),
.Y(n_6053)
);

OAI21xp5_ASAP7_75t_L g6054 ( 
.A1(n_5498),
.A2(n_3816),
.B(n_3714),
.Y(n_6054)
);

OAI21x1_ASAP7_75t_L g6055 ( 
.A1(n_5741),
.A2(n_3470),
.B(n_3469),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5574),
.Y(n_6056)
);

A2O1A1Ixp33_ASAP7_75t_L g6057 ( 
.A1(n_5504),
.A2(n_1270),
.B(n_1242),
.C(n_1530),
.Y(n_6057)
);

OAI21xp5_ASAP7_75t_L g6058 ( 
.A1(n_5532),
.A2(n_3816),
.B(n_3714),
.Y(n_6058)
);

OAI21x1_ASAP7_75t_L g6059 ( 
.A1(n_5724),
.A2(n_3470),
.B(n_3469),
.Y(n_6059)
);

NAND2xp5_ASAP7_75t_SL g6060 ( 
.A(n_5588),
.B(n_1530),
.Y(n_6060)
);

OAI21x1_ASAP7_75t_L g6061 ( 
.A1(n_5635),
.A2(n_3477),
.B(n_3473),
.Y(n_6061)
);

OAI21x1_ASAP7_75t_L g6062 ( 
.A1(n_5643),
.A2(n_3477),
.B(n_3473),
.Y(n_6062)
);

BUFx6f_ASAP7_75t_L g6063 ( 
.A(n_5606),
.Y(n_6063)
);

AOI21xp5_ASAP7_75t_SL g6064 ( 
.A1(n_5680),
.A2(n_4004),
.B(n_3990),
.Y(n_6064)
);

NAND2xp5_ASAP7_75t_L g6065 ( 
.A(n_5393),
.B(n_26),
.Y(n_6065)
);

OAI21x1_ASAP7_75t_L g6066 ( 
.A1(n_5686),
.A2(n_3479),
.B(n_3478),
.Y(n_6066)
);

OAI21x1_ASAP7_75t_L g6067 ( 
.A1(n_5668),
.A2(n_3479),
.B(n_3478),
.Y(n_6067)
);

OAI22xp5_ASAP7_75t_L g6068 ( 
.A1(n_5449),
.A2(n_4004),
.B1(n_4007),
.B2(n_3990),
.Y(n_6068)
);

OA21x2_ASAP7_75t_L g6069 ( 
.A1(n_5624),
.A2(n_3092),
.B(n_3090),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5397),
.Y(n_6070)
);

OAI21x1_ASAP7_75t_L g6071 ( 
.A1(n_5415),
.A2(n_3485),
.B(n_3324),
.Y(n_6071)
);

BUFx10_ASAP7_75t_L g6072 ( 
.A(n_5473),
.Y(n_6072)
);

CKINVDCx5p33_ASAP7_75t_R g6073 ( 
.A(n_5663),
.Y(n_6073)
);

AND2x4_ASAP7_75t_L g6074 ( 
.A(n_5559),
.B(n_4004),
.Y(n_6074)
);

INVx2_ASAP7_75t_SL g6075 ( 
.A(n_5358),
.Y(n_6075)
);

NAND2x1p5_ASAP7_75t_L g6076 ( 
.A(n_5551),
.B(n_4007),
.Y(n_6076)
);

NAND2xp5_ASAP7_75t_SL g6077 ( 
.A(n_5756),
.B(n_1577),
.Y(n_6077)
);

OAI21x1_ASAP7_75t_L g6078 ( 
.A1(n_5584),
.A2(n_3485),
.B(n_3324),
.Y(n_6078)
);

NAND2xp5_ASAP7_75t_L g6079 ( 
.A(n_5399),
.B(n_28),
.Y(n_6079)
);

A2O1A1Ixp33_ASAP7_75t_L g6080 ( 
.A1(n_5541),
.A2(n_1577),
.B(n_32),
.C(n_29),
.Y(n_6080)
);

INVx3_ASAP7_75t_L g6081 ( 
.A(n_5376),
.Y(n_6081)
);

NAND2xp5_ASAP7_75t_L g6082 ( 
.A(n_5438),
.B(n_30),
.Y(n_6082)
);

AND2x2_ASAP7_75t_L g6083 ( 
.A(n_5428),
.B(n_30),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5464),
.Y(n_6084)
);

A2O1A1Ixp33_ASAP7_75t_L g6085 ( 
.A1(n_5546),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_5487),
.B(n_34),
.Y(n_6086)
);

BUFx6f_ASAP7_75t_L g6087 ( 
.A(n_5606),
.Y(n_6087)
);

NAND2xp5_ASAP7_75t_L g6088 ( 
.A(n_5675),
.B(n_38),
.Y(n_6088)
);

INVx3_ASAP7_75t_L g6089 ( 
.A(n_5376),
.Y(n_6089)
);

OAI21x1_ASAP7_75t_L g6090 ( 
.A1(n_5372),
.A2(n_3333),
.B(n_3318),
.Y(n_6090)
);

OAI21x1_ASAP7_75t_L g6091 ( 
.A1(n_5396),
.A2(n_3333),
.B(n_3318),
.Y(n_6091)
);

OAI21x1_ASAP7_75t_L g6092 ( 
.A1(n_5671),
.A2(n_5743),
.B(n_5499),
.Y(n_6092)
);

AO21x1_ASAP7_75t_L g6093 ( 
.A1(n_5761),
.A2(n_39),
.B(n_40),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_5620),
.B(n_40),
.Y(n_6094)
);

AOI21xp5_ASAP7_75t_L g6095 ( 
.A1(n_5495),
.A2(n_4015),
.B(n_4007),
.Y(n_6095)
);

O2A1O1Ixp33_ASAP7_75t_L g6096 ( 
.A1(n_5413),
.A2(n_3092),
.B(n_3101),
.C(n_3090),
.Y(n_6096)
);

OAI21xp33_ASAP7_75t_L g6097 ( 
.A1(n_5611),
.A2(n_2466),
.B(n_3101),
.Y(n_6097)
);

BUFx2_ASAP7_75t_L g6098 ( 
.A(n_5519),
.Y(n_6098)
);

OAI21x1_ASAP7_75t_L g6099 ( 
.A1(n_5743),
.A2(n_5492),
.B(n_5709),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_5594),
.Y(n_6100)
);

AO22x2_ASAP7_75t_L g6101 ( 
.A1(n_5539),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_6101)
);

OAI21xp5_ASAP7_75t_L g6102 ( 
.A1(n_5611),
.A2(n_5537),
.B(n_5744),
.Y(n_6102)
);

AND2x4_ASAP7_75t_L g6103 ( 
.A(n_5559),
.B(n_4015),
.Y(n_6103)
);

NOR2xp33_ASAP7_75t_SL g6104 ( 
.A(n_5553),
.B(n_3697),
.Y(n_6104)
);

AOI22xp5_ASAP7_75t_L g6105 ( 
.A1(n_5561),
.A2(n_3697),
.B1(n_3724),
.B2(n_3714),
.Y(n_6105)
);

NOR2x1_ASAP7_75t_SL g6106 ( 
.A(n_5533),
.B(n_4063),
.Y(n_6106)
);

NAND2xp5_ASAP7_75t_L g6107 ( 
.A(n_5708),
.B(n_41),
.Y(n_6107)
);

OAI21x1_ASAP7_75t_L g6108 ( 
.A1(n_5715),
.A2(n_3106),
.B(n_3104),
.Y(n_6108)
);

AOI21xp5_ASAP7_75t_L g6109 ( 
.A1(n_5495),
.A2(n_4063),
.B(n_3106),
.Y(n_6109)
);

BUFx2_ASAP7_75t_L g6110 ( 
.A(n_5519),
.Y(n_6110)
);

O2A1O1Ixp5_ASAP7_75t_L g6111 ( 
.A1(n_5579),
.A2(n_3110),
.B(n_3112),
.C(n_3104),
.Y(n_6111)
);

NOR2xp33_ASAP7_75t_SL g6112 ( 
.A(n_5553),
.B(n_3697),
.Y(n_6112)
);

OAI21x1_ASAP7_75t_L g6113 ( 
.A1(n_5458),
.A2(n_3112),
.B(n_3110),
.Y(n_6113)
);

AOI21xp5_ASAP7_75t_L g6114 ( 
.A1(n_5645),
.A2(n_3120),
.B(n_3114),
.Y(n_6114)
);

OAI21x1_ASAP7_75t_L g6115 ( 
.A1(n_5458),
.A2(n_3120),
.B(n_3114),
.Y(n_6115)
);

AOI21x1_ASAP7_75t_L g6116 ( 
.A1(n_5761),
.A2(n_3125),
.B(n_3123),
.Y(n_6116)
);

AOI21xp5_ASAP7_75t_L g6117 ( 
.A1(n_5645),
.A2(n_3125),
.B(n_3123),
.Y(n_6117)
);

NAND2xp5_ASAP7_75t_L g6118 ( 
.A(n_5739),
.B(n_44),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5612),
.Y(n_6119)
);

AND2x6_ASAP7_75t_L g6120 ( 
.A(n_5771),
.B(n_3126),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_L g6121 ( 
.A(n_5581),
.B(n_44),
.Y(n_6121)
);

OAI21x1_ASAP7_75t_L g6122 ( 
.A1(n_5471),
.A2(n_3138),
.B(n_3126),
.Y(n_6122)
);

AOI21x1_ASAP7_75t_SL g6123 ( 
.A1(n_5681),
.A2(n_45),
.B(n_46),
.Y(n_6123)
);

NAND2xp5_ASAP7_75t_L g6124 ( 
.A(n_5622),
.B(n_46),
.Y(n_6124)
);

OAI21xp5_ASAP7_75t_L g6125 ( 
.A1(n_5670),
.A2(n_3816),
.B(n_3724),
.Y(n_6125)
);

NOR2x1_ASAP7_75t_L g6126 ( 
.A(n_5471),
.B(n_3138),
.Y(n_6126)
);

NAND2xp5_ASAP7_75t_L g6127 ( 
.A(n_5647),
.B(n_47),
.Y(n_6127)
);

HB1xp67_ASAP7_75t_L g6128 ( 
.A(n_5719),
.Y(n_6128)
);

CKINVDCx5p33_ASAP7_75t_R g6129 ( 
.A(n_5710),
.Y(n_6129)
);

OAI21xp5_ASAP7_75t_L g6130 ( 
.A1(n_5600),
.A2(n_3816),
.B(n_3724),
.Y(n_6130)
);

OAI21xp33_ASAP7_75t_L g6131 ( 
.A1(n_5738),
.A2(n_2466),
.B(n_3147),
.Y(n_6131)
);

BUFx5_ASAP7_75t_L g6132 ( 
.A(n_5519),
.Y(n_6132)
);

BUFx4_ASAP7_75t_SL g6133 ( 
.A(n_5473),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_5533),
.Y(n_6134)
);

OAI22xp5_ASAP7_75t_L g6135 ( 
.A1(n_5419),
.A2(n_3147),
.B1(n_3150),
.B2(n_3148),
.Y(n_6135)
);

OAI21x1_ASAP7_75t_L g6136 ( 
.A1(n_5491),
.A2(n_5549),
.B(n_5515),
.Y(n_6136)
);

NAND2xp5_ASAP7_75t_L g6137 ( 
.A(n_5730),
.B(n_47),
.Y(n_6137)
);

INVx2_ASAP7_75t_L g6138 ( 
.A(n_5890),
.Y(n_6138)
);

NOR2x1_ASAP7_75t_L g6139 ( 
.A(n_5953),
.B(n_5491),
.Y(n_6139)
);

AO21x2_ASAP7_75t_L g6140 ( 
.A1(n_6134),
.A2(n_5482),
.B(n_5682),
.Y(n_6140)
);

INVx8_ASAP7_75t_L g6141 ( 
.A(n_5783),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_5802),
.Y(n_6142)
);

INVx3_ASAP7_75t_L g6143 ( 
.A(n_5829),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_5802),
.Y(n_6144)
);

NAND2xp5_ASAP7_75t_SL g6145 ( 
.A(n_5835),
.B(n_5764),
.Y(n_6145)
);

OA21x2_ASAP7_75t_L g6146 ( 
.A1(n_5819),
.A2(n_5656),
.B(n_5665),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_5808),
.Y(n_6147)
);

AOI22x1_ASAP7_75t_L g6148 ( 
.A1(n_6101),
.A2(n_5697),
.B1(n_5770),
.B2(n_5474),
.Y(n_6148)
);

BUFx3_ASAP7_75t_L g6149 ( 
.A(n_5841),
.Y(n_6149)
);

INVx1_ASAP7_75t_L g6150 ( 
.A(n_5808),
.Y(n_6150)
);

OAI21x1_ASAP7_75t_L g6151 ( 
.A1(n_5860),
.A2(n_5539),
.B(n_5515),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5822),
.Y(n_6152)
);

HB1xp67_ASAP7_75t_L g6153 ( 
.A(n_6128),
.Y(n_6153)
);

BUFx6f_ASAP7_75t_L g6154 ( 
.A(n_5980),
.Y(n_6154)
);

INVx3_ASAP7_75t_L g6155 ( 
.A(n_5829),
.Y(n_6155)
);

OAI21x1_ASAP7_75t_SL g6156 ( 
.A1(n_5846),
.A2(n_6046),
.B(n_6038),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_5909),
.Y(n_6157)
);

AO21x2_ASAP7_75t_L g6158 ( 
.A1(n_6134),
.A2(n_5718),
.B(n_5696),
.Y(n_6158)
);

NAND2xp5_ASAP7_75t_L g6159 ( 
.A(n_6056),
.B(n_5719),
.Y(n_6159)
);

CKINVDCx5p33_ASAP7_75t_R g6160 ( 
.A(n_5943),
.Y(n_6160)
);

INVx3_ASAP7_75t_L g6161 ( 
.A(n_5818),
.Y(n_6161)
);

AO21x2_ASAP7_75t_L g6162 ( 
.A1(n_5953),
.A2(n_5703),
.B(n_5691),
.Y(n_6162)
);

AOI22xp33_ASAP7_75t_L g6163 ( 
.A1(n_5857),
.A2(n_5738),
.B1(n_5614),
.B2(n_5417),
.Y(n_6163)
);

INVx3_ASAP7_75t_L g6164 ( 
.A(n_5818),
.Y(n_6164)
);

AND2x4_ASAP7_75t_L g6165 ( 
.A(n_6098),
.B(n_5549),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5822),
.Y(n_6166)
);

AO21x1_ASAP7_75t_L g6167 ( 
.A1(n_5981),
.A2(n_5472),
.B(n_5597),
.Y(n_6167)
);

OAI21x1_ASAP7_75t_L g6168 ( 
.A1(n_5782),
.A2(n_5572),
.B(n_5563),
.Y(n_6168)
);

INVx8_ASAP7_75t_L g6169 ( 
.A(n_5783),
.Y(n_6169)
);

OAI21x1_ASAP7_75t_L g6170 ( 
.A1(n_5792),
.A2(n_5572),
.B(n_5563),
.Y(n_6170)
);

BUFx12f_ASAP7_75t_L g6171 ( 
.A(n_6073),
.Y(n_6171)
);

BUFx3_ASAP7_75t_L g6172 ( 
.A(n_5980),
.Y(n_6172)
);

INVx5_ASAP7_75t_L g6173 ( 
.A(n_5809),
.Y(n_6173)
);

OR2x6_ASAP7_75t_L g6174 ( 
.A(n_5915),
.B(n_5651),
.Y(n_6174)
);

INVx2_ASAP7_75t_SL g6175 ( 
.A(n_5809),
.Y(n_6175)
);

BUFx12f_ASAP7_75t_L g6176 ( 
.A(n_5790),
.Y(n_6176)
);

INVx1_ASAP7_75t_SL g6177 ( 
.A(n_5895),
.Y(n_6177)
);

INVx2_ASAP7_75t_L g6178 ( 
.A(n_6084),
.Y(n_6178)
);

NAND2x1p5_ASAP7_75t_L g6179 ( 
.A(n_6069),
.B(n_5770),
.Y(n_6179)
);

AO21x2_ASAP7_75t_L g6180 ( 
.A1(n_6106),
.A2(n_5712),
.B(n_5605),
.Y(n_6180)
);

AO21x1_ASAP7_75t_SL g6181 ( 
.A1(n_5781),
.A2(n_5736),
.B(n_5676),
.Y(n_6181)
);

INVx2_ASAP7_75t_L g6182 ( 
.A(n_6084),
.Y(n_6182)
);

BUFx3_ASAP7_75t_L g6183 ( 
.A(n_6129),
.Y(n_6183)
);

BUFx3_ASAP7_75t_L g6184 ( 
.A(n_5850),
.Y(n_6184)
);

BUFx2_ASAP7_75t_R g6185 ( 
.A(n_5899),
.Y(n_6185)
);

OR2x2_ASAP7_75t_L g6186 ( 
.A(n_5798),
.B(n_5655),
.Y(n_6186)
);

BUFx3_ASAP7_75t_L g6187 ( 
.A(n_5850),
.Y(n_6187)
);

BUFx6f_ASAP7_75t_L g6188 ( 
.A(n_5814),
.Y(n_6188)
);

INVx2_ASAP7_75t_L g6189 ( 
.A(n_6100),
.Y(n_6189)
);

OA21x2_ASAP7_75t_L g6190 ( 
.A1(n_6092),
.A2(n_5630),
.B(n_5547),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5933),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_5933),
.Y(n_6192)
);

INVx3_ASAP7_75t_L g6193 ( 
.A(n_6136),
.Y(n_6193)
);

HB1xp67_ASAP7_75t_L g6194 ( 
.A(n_5965),
.Y(n_6194)
);

NOR2xp33_ASAP7_75t_L g6195 ( 
.A(n_5889),
.B(n_5429),
.Y(n_6195)
);

BUFx3_ASAP7_75t_L g6196 ( 
.A(n_5814),
.Y(n_6196)
);

INVx2_ASAP7_75t_L g6197 ( 
.A(n_6100),
.Y(n_6197)
);

BUFx2_ASAP7_75t_R g6198 ( 
.A(n_6133),
.Y(n_6198)
);

BUFx3_ASAP7_75t_L g6199 ( 
.A(n_6051),
.Y(n_6199)
);

OAI21x1_ASAP7_75t_SL g6200 ( 
.A1(n_6093),
.A2(n_5390),
.B(n_5750),
.Y(n_6200)
);

CKINVDCx6p67_ASAP7_75t_R g6201 ( 
.A(n_6072),
.Y(n_6201)
);

OAI21x1_ASAP7_75t_L g6202 ( 
.A1(n_5785),
.A2(n_5771),
.B(n_5711),
.Y(n_6202)
);

OR2x6_ASAP7_75t_L g6203 ( 
.A(n_5864),
.B(n_5651),
.Y(n_6203)
);

INVx3_ASAP7_75t_L g6204 ( 
.A(n_5941),
.Y(n_6204)
);

INVx2_ASAP7_75t_L g6205 ( 
.A(n_6119),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5965),
.Y(n_6206)
);

BUFx6f_ASAP7_75t_L g6207 ( 
.A(n_5814),
.Y(n_6207)
);

INVx2_ASAP7_75t_SL g6208 ( 
.A(n_5939),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_5970),
.Y(n_6209)
);

AO21x2_ASAP7_75t_L g6210 ( 
.A1(n_5886),
.A2(n_5737),
.B(n_5767),
.Y(n_6210)
);

INVx4_ASAP7_75t_L g6211 ( 
.A(n_5903),
.Y(n_6211)
);

AND2x4_ASAP7_75t_L g6212 ( 
.A(n_6110),
.B(n_5519),
.Y(n_6212)
);

INVx5_ASAP7_75t_L g6213 ( 
.A(n_5930),
.Y(n_6213)
);

NOR2xp33_ASAP7_75t_L g6214 ( 
.A(n_5786),
.B(n_5916),
.Y(n_6214)
);

INVx2_ASAP7_75t_L g6215 ( 
.A(n_6119),
.Y(n_6215)
);

BUFx6f_ASAP7_75t_L g6216 ( 
.A(n_5939),
.Y(n_6216)
);

BUFx3_ASAP7_75t_L g6217 ( 
.A(n_5885),
.Y(n_6217)
);

INVx8_ASAP7_75t_L g6218 ( 
.A(n_5877),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_5970),
.Y(n_6219)
);

OAI21x1_ASAP7_75t_SL g6220 ( 
.A1(n_5903),
.A2(n_5722),
.B(n_5731),
.Y(n_6220)
);

BUFx6f_ASAP7_75t_L g6221 ( 
.A(n_5939),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_5983),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5983),
.Y(n_6223)
);

AOI22xp5_ASAP7_75t_L g6224 ( 
.A1(n_5948),
.A2(n_5407),
.B1(n_5470),
.B2(n_5543),
.Y(n_6224)
);

INVx2_ASAP7_75t_SL g6225 ( 
.A(n_5843),
.Y(n_6225)
);

INVx3_ASAP7_75t_L g6226 ( 
.A(n_5941),
.Y(n_6226)
);

AND2x2_ASAP7_75t_L g6227 ( 
.A(n_5904),
.B(n_5766),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_6056),
.B(n_5666),
.Y(n_6228)
);

INVx1_ASAP7_75t_SL g6229 ( 
.A(n_6081),
.Y(n_6229)
);

BUFx12f_ASAP7_75t_L g6230 ( 
.A(n_6050),
.Y(n_6230)
);

INVx2_ASAP7_75t_L g6231 ( 
.A(n_5919),
.Y(n_6231)
);

AO21x2_ASAP7_75t_L g6232 ( 
.A1(n_5925),
.A2(n_5760),
.B(n_5524),
.Y(n_6232)
);

BUFx2_ASAP7_75t_R g6233 ( 
.A(n_5817),
.Y(n_6233)
);

INVx8_ASAP7_75t_L g6234 ( 
.A(n_6120),
.Y(n_6234)
);

INVx2_ASAP7_75t_L g6235 ( 
.A(n_5952),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_6027),
.Y(n_6236)
);

INVx3_ASAP7_75t_L g6237 ( 
.A(n_6081),
.Y(n_6237)
);

INVx5_ASAP7_75t_L g6238 ( 
.A(n_5930),
.Y(n_6238)
);

BUFx4_ASAP7_75t_SL g6239 ( 
.A(n_5947),
.Y(n_6239)
);

OA21x2_ASAP7_75t_L g6240 ( 
.A1(n_6099),
.A2(n_5695),
.B(n_5523),
.Y(n_6240)
);

BUFx12f_ASAP7_75t_L g6241 ( 
.A(n_6050),
.Y(n_6241)
);

AND2x4_ASAP7_75t_L g6242 ( 
.A(n_6089),
.B(n_5706),
.Y(n_6242)
);

OAI21x1_ASAP7_75t_L g6243 ( 
.A1(n_5796),
.A2(n_5711),
.B(n_5666),
.Y(n_6243)
);

BUFx6f_ASAP7_75t_L g6244 ( 
.A(n_5984),
.Y(n_6244)
);

BUFx2_ASAP7_75t_L g6245 ( 
.A(n_5908),
.Y(n_6245)
);

OR2x6_ASAP7_75t_L g6246 ( 
.A(n_5921),
.B(n_5651),
.Y(n_6246)
);

AOI22x1_ASAP7_75t_L g6247 ( 
.A1(n_6101),
.A2(n_5700),
.B1(n_5687),
.B2(n_5732),
.Y(n_6247)
);

BUFx3_ASAP7_75t_L g6248 ( 
.A(n_5861),
.Y(n_6248)
);

AND2x2_ASAP7_75t_L g6249 ( 
.A(n_6019),
.B(n_5657),
.Y(n_6249)
);

AO21x2_ASAP7_75t_L g6250 ( 
.A1(n_5797),
.A2(n_5758),
.B(n_5609),
.Y(n_6250)
);

AND2x4_ASAP7_75t_L g6251 ( 
.A(n_6089),
.B(n_5714),
.Y(n_6251)
);

INVx6_ASAP7_75t_SL g6252 ( 
.A(n_6072),
.Y(n_6252)
);

AOI21x1_ASAP7_75t_L g6253 ( 
.A1(n_5968),
.A2(n_3150),
.B(n_3148),
.Y(n_6253)
);

INVx2_ASAP7_75t_L g6254 ( 
.A(n_5988),
.Y(n_6254)
);

INVx3_ASAP7_75t_L g6255 ( 
.A(n_5908),
.Y(n_6255)
);

INVx6_ASAP7_75t_SL g6256 ( 
.A(n_6074),
.Y(n_6256)
);

NAND2xp5_ASAP7_75t_L g6257 ( 
.A(n_5779),
.B(n_5617),
.Y(n_6257)
);

OAI21x1_ASAP7_75t_L g6258 ( 
.A1(n_5788),
.A2(n_5805),
.B(n_5945),
.Y(n_6258)
);

BUFx3_ASAP7_75t_L g6259 ( 
.A(n_5898),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_6027),
.Y(n_6260)
);

HB1xp67_ASAP7_75t_L g6261 ( 
.A(n_5991),
.Y(n_6261)
);

INVx2_ASAP7_75t_L g6262 ( 
.A(n_6010),
.Y(n_6262)
);

AND2x4_ASAP7_75t_L g6263 ( 
.A(n_6005),
.B(n_5723),
.Y(n_6263)
);

OAI21x1_ASAP7_75t_L g6264 ( 
.A1(n_5945),
.A2(n_5603),
.B(n_5717),
.Y(n_6264)
);

AOI22xp33_ASAP7_75t_L g6265 ( 
.A1(n_5914),
.A2(n_5725),
.B1(n_5756),
.B2(n_5749),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_5795),
.Y(n_6266)
);

INVx3_ASAP7_75t_L g6267 ( 
.A(n_6005),
.Y(n_6267)
);

OAI21x1_ASAP7_75t_L g6268 ( 
.A1(n_5812),
.A2(n_3399),
.B(n_3389),
.Y(n_6268)
);

AND2x4_ASAP7_75t_L g6269 ( 
.A(n_6044),
.B(n_5756),
.Y(n_6269)
);

OAI21xp5_ASAP7_75t_L g6270 ( 
.A1(n_5855),
.A2(n_5897),
.B(n_5803),
.Y(n_6270)
);

BUFx3_ASAP7_75t_L g6271 ( 
.A(n_5972),
.Y(n_6271)
);

BUFx3_ASAP7_75t_L g6272 ( 
.A(n_6044),
.Y(n_6272)
);

INVx2_ASAP7_75t_L g6273 ( 
.A(n_5847),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5871),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5887),
.Y(n_6275)
);

OAI21x1_ASAP7_75t_L g6276 ( 
.A1(n_6004),
.A2(n_5892),
.B(n_5989),
.Y(n_6276)
);

OAI21x1_ASAP7_75t_L g6277 ( 
.A1(n_5799),
.A2(n_3399),
.B(n_3389),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_6030),
.Y(n_6278)
);

OAI21x1_ASAP7_75t_L g6279 ( 
.A1(n_5910),
.A2(n_3399),
.B(n_3389),
.Y(n_6279)
);

AO21x2_ASAP7_75t_L g6280 ( 
.A1(n_5882),
.A2(n_3160),
.B(n_3153),
.Y(n_6280)
);

INVx3_ASAP7_75t_L g6281 ( 
.A(n_5932),
.Y(n_6281)
);

OAI21xp5_ASAP7_75t_L g6282 ( 
.A1(n_5955),
.A2(n_5959),
.B(n_6008),
.Y(n_6282)
);

BUFx10_ASAP7_75t_L g6283 ( 
.A(n_6022),
.Y(n_6283)
);

NAND2x1p5_ASAP7_75t_L g6284 ( 
.A(n_6069),
.B(n_5545),
.Y(n_6284)
);

AO21x2_ASAP7_75t_L g6285 ( 
.A1(n_5884),
.A2(n_3160),
.B(n_3153),
.Y(n_6285)
);

INVx4_ASAP7_75t_L g6286 ( 
.A(n_5932),
.Y(n_6286)
);

HB1xp67_ASAP7_75t_L g6287 ( 
.A(n_5987),
.Y(n_6287)
);

OAI21xp5_ASAP7_75t_L g6288 ( 
.A1(n_5959),
.A2(n_5545),
.B(n_3724),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6070),
.Y(n_6289)
);

OAI21x1_ASAP7_75t_L g6290 ( 
.A1(n_6055),
.A2(n_3399),
.B(n_3389),
.Y(n_6290)
);

AO21x2_ASAP7_75t_L g6291 ( 
.A1(n_5856),
.A2(n_3166),
.B(n_3164),
.Y(n_6291)
);

NOR2xp33_ASAP7_75t_L g6292 ( 
.A(n_5986),
.B(n_5749),
.Y(n_6292)
);

AND2x4_ASAP7_75t_L g6293 ( 
.A(n_6075),
.B(n_5617),
.Y(n_6293)
);

AND2x4_ASAP7_75t_L g6294 ( 
.A(n_5985),
.B(n_5617),
.Y(n_6294)
);

AOI21x1_ASAP7_75t_L g6295 ( 
.A1(n_5893),
.A2(n_3166),
.B(n_3164),
.Y(n_6295)
);

BUFx3_ASAP7_75t_L g6296 ( 
.A(n_5984),
.Y(n_6296)
);

OAI21x1_ASAP7_75t_L g6297 ( 
.A1(n_5917),
.A2(n_3419),
.B(n_3408),
.Y(n_6297)
);

AO21x2_ASAP7_75t_L g6298 ( 
.A1(n_5997),
.A2(n_3170),
.B(n_3169),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6042),
.Y(n_6299)
);

INVx6_ASAP7_75t_L g6300 ( 
.A(n_5984),
.Y(n_6300)
);

CKINVDCx5p33_ASAP7_75t_R g6301 ( 
.A(n_5938),
.Y(n_6301)
);

INVx2_ASAP7_75t_L g6302 ( 
.A(n_5866),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_5975),
.Y(n_6303)
);

BUFx2_ASAP7_75t_SL g6304 ( 
.A(n_5828),
.Y(n_6304)
);

BUFx12f_ASAP7_75t_L g6305 ( 
.A(n_5967),
.Y(n_6305)
);

OAI21xp5_ASAP7_75t_L g6306 ( 
.A1(n_6008),
.A2(n_3724),
.B(n_3714),
.Y(n_6306)
);

AOI22x1_ASAP7_75t_L g6307 ( 
.A1(n_5923),
.A2(n_5749),
.B1(n_5688),
.B2(n_5713),
.Y(n_6307)
);

CKINVDCx20_ASAP7_75t_R g6308 ( 
.A(n_6083),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_5931),
.Y(n_6309)
);

BUFx6f_ASAP7_75t_L g6310 ( 
.A(n_6023),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_5928),
.Y(n_6311)
);

BUFx6f_ASAP7_75t_L g6312 ( 
.A(n_6023),
.Y(n_6312)
);

AO21x2_ASAP7_75t_L g6313 ( 
.A1(n_5827),
.A2(n_3170),
.B(n_3169),
.Y(n_6313)
);

AO21x1_ASAP7_75t_L g6314 ( 
.A1(n_6034),
.A2(n_48),
.B(n_49),
.Y(n_6314)
);

NAND2x1p5_ASAP7_75t_L g6315 ( 
.A(n_5823),
.B(n_5669),
.Y(n_6315)
);

NAND2xp5_ASAP7_75t_L g6316 ( 
.A(n_5879),
.B(n_5669),
.Y(n_6316)
);

BUFx2_ASAP7_75t_L g6317 ( 
.A(n_6020),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_5987),
.Y(n_6318)
);

INVx5_ASAP7_75t_L g6319 ( 
.A(n_6120),
.Y(n_6319)
);

INVx3_ASAP7_75t_L g6320 ( 
.A(n_6020),
.Y(n_6320)
);

OAI21xp5_ASAP7_75t_L g6321 ( 
.A1(n_6012),
.A2(n_3714),
.B(n_3175),
.Y(n_6321)
);

OAI21x1_ASAP7_75t_L g6322 ( 
.A1(n_5804),
.A2(n_3419),
.B(n_3408),
.Y(n_6322)
);

OAI21x1_ASAP7_75t_L g6323 ( 
.A1(n_5813),
.A2(n_3419),
.B(n_3408),
.Y(n_6323)
);

BUFx5_ASAP7_75t_L g6324 ( 
.A(n_6120),
.Y(n_6324)
);

OAI21xp5_ASAP7_75t_L g6325 ( 
.A1(n_6012),
.A2(n_3175),
.B(n_3171),
.Y(n_6325)
);

CKINVDCx16_ASAP7_75t_R g6326 ( 
.A(n_5966),
.Y(n_6326)
);

OR2x2_ASAP7_75t_L g6327 ( 
.A(n_5973),
.B(n_5669),
.Y(n_6327)
);

OAI21x1_ASAP7_75t_L g6328 ( 
.A1(n_5880),
.A2(n_3419),
.B(n_3408),
.Y(n_6328)
);

NAND2x1p5_ASAP7_75t_L g6329 ( 
.A(n_6126),
.B(n_5688),
.Y(n_6329)
);

INVx8_ASAP7_75t_L g6330 ( 
.A(n_6120),
.Y(n_6330)
);

AO21x2_ASAP7_75t_L g6331 ( 
.A1(n_5830),
.A2(n_3176),
.B(n_3171),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_5793),
.Y(n_6332)
);

BUFx4_ASAP7_75t_R g6333 ( 
.A(n_6132),
.Y(n_6333)
);

INVx3_ASAP7_75t_L g6334 ( 
.A(n_6023),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_5987),
.Y(n_6335)
);

INVx2_ASAP7_75t_L g6336 ( 
.A(n_5883),
.Y(n_6336)
);

BUFx3_ASAP7_75t_L g6337 ( 
.A(n_6041),
.Y(n_6337)
);

BUFx2_ASAP7_75t_SL g6338 ( 
.A(n_5901),
.Y(n_6338)
);

OAI21xp33_ASAP7_75t_L g6339 ( 
.A1(n_6080),
.A2(n_48),
.B(n_50),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_5996),
.Y(n_6340)
);

INVx2_ASAP7_75t_L g6341 ( 
.A(n_5883),
.Y(n_6341)
);

CKINVDCx14_ASAP7_75t_R g6342 ( 
.A(n_6032),
.Y(n_6342)
);

OAI21x1_ASAP7_75t_L g6343 ( 
.A1(n_5900),
.A2(n_3466),
.B(n_3182),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_5996),
.Y(n_6344)
);

BUFx4_ASAP7_75t_SL g6345 ( 
.A(n_5902),
.Y(n_6345)
);

BUFx12f_ASAP7_75t_L g6346 ( 
.A(n_6017),
.Y(n_6346)
);

INVx3_ASAP7_75t_L g6347 ( 
.A(n_6041),
.Y(n_6347)
);

NAND2x1p5_ASAP7_75t_L g6348 ( 
.A(n_6126),
.B(n_5688),
.Y(n_6348)
);

BUFx6f_ASAP7_75t_L g6349 ( 
.A(n_6041),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_5996),
.Y(n_6350)
);

AOI21xp5_ASAP7_75t_L g6351 ( 
.A1(n_6114),
.A2(n_5713),
.B(n_2721),
.Y(n_6351)
);

OAI21x1_ASAP7_75t_L g6352 ( 
.A1(n_5780),
.A2(n_3466),
.B(n_3182),
.Y(n_6352)
);

NAND2x1p5_ASAP7_75t_L g6353 ( 
.A(n_5985),
.B(n_5713),
.Y(n_6353)
);

OAI21x1_ASAP7_75t_L g6354 ( 
.A1(n_5842),
.A2(n_3466),
.B(n_3187),
.Y(n_6354)
);

NAND2x1p5_ASAP7_75t_L g6355 ( 
.A(n_5912),
.B(n_2628),
.Y(n_6355)
);

BUFx3_ASAP7_75t_L g6356 ( 
.A(n_6063),
.Y(n_6356)
);

OAI21x1_ASAP7_75t_L g6357 ( 
.A1(n_5888),
.A2(n_3466),
.B(n_3187),
.Y(n_6357)
);

INVx2_ASAP7_75t_SL g6358 ( 
.A(n_6063),
.Y(n_6358)
);

BUFx3_ASAP7_75t_L g6359 ( 
.A(n_6063),
.Y(n_6359)
);

BUFx2_ASAP7_75t_L g6360 ( 
.A(n_6132),
.Y(n_6360)
);

BUFx3_ASAP7_75t_L g6361 ( 
.A(n_6087),
.Y(n_6361)
);

BUFx12f_ASAP7_75t_L g6362 ( 
.A(n_5974),
.Y(n_6362)
);

BUFx2_ASAP7_75t_SL g6363 ( 
.A(n_6132),
.Y(n_6363)
);

INVxp67_ASAP7_75t_SL g6364 ( 
.A(n_5863),
.Y(n_6364)
);

OAI21x1_ASAP7_75t_L g6365 ( 
.A1(n_5891),
.A2(n_3188),
.B(n_3176),
.Y(n_6365)
);

OAI21x1_ASAP7_75t_L g6366 ( 
.A1(n_5837),
.A2(n_3192),
.B(n_3188),
.Y(n_6366)
);

OAI21x1_ASAP7_75t_L g6367 ( 
.A1(n_5870),
.A2(n_3208),
.B(n_3192),
.Y(n_6367)
);

INVx2_ASAP7_75t_R g6368 ( 
.A(n_6132),
.Y(n_6368)
);

AO21x2_ASAP7_75t_L g6369 ( 
.A1(n_6118),
.A2(n_3209),
.B(n_3208),
.Y(n_6369)
);

NAND2x1p5_ASAP7_75t_L g6370 ( 
.A(n_5951),
.B(n_2628),
.Y(n_6370)
);

CKINVDCx16_ASAP7_75t_R g6371 ( 
.A(n_5966),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6007),
.Y(n_6372)
);

OAI21x1_ASAP7_75t_L g6373 ( 
.A1(n_6021),
.A2(n_3219),
.B(n_3209),
.Y(n_6373)
);

INVx1_ASAP7_75t_SL g6374 ( 
.A(n_5854),
.Y(n_6374)
);

BUFx3_ASAP7_75t_L g6375 ( 
.A(n_6087),
.Y(n_6375)
);

OR3x4_ASAP7_75t_SL g6376 ( 
.A(n_5914),
.B(n_50),
.C(n_51),
.Y(n_6376)
);

AO21x2_ASAP7_75t_L g6377 ( 
.A1(n_5867),
.A2(n_3221),
.B(n_3219),
.Y(n_6377)
);

AND2x4_ASAP7_75t_L g6378 ( 
.A(n_5800),
.B(n_51),
.Y(n_6378)
);

AOI21xp5_ASAP7_75t_L g6379 ( 
.A1(n_6117),
.A2(n_2723),
.B(n_2721),
.Y(n_6379)
);

BUFx3_ASAP7_75t_L g6380 ( 
.A(n_6087),
.Y(n_6380)
);

BUFx6f_ASAP7_75t_L g6381 ( 
.A(n_6074),
.Y(n_6381)
);

NAND2x1p5_ASAP7_75t_L g6382 ( 
.A(n_6095),
.B(n_2721),
.Y(n_6382)
);

AND2x4_ASAP7_75t_L g6383 ( 
.A(n_6047),
.B(n_52),
.Y(n_6383)
);

AO21x2_ASAP7_75t_L g6384 ( 
.A1(n_5874),
.A2(n_3221),
.B(n_3220),
.Y(n_6384)
);

OAI21x1_ASAP7_75t_L g6385 ( 
.A1(n_5944),
.A2(n_5950),
.B(n_5848),
.Y(n_6385)
);

INVx3_ASAP7_75t_L g6386 ( 
.A(n_6132),
.Y(n_6386)
);

OAI21x1_ASAP7_75t_L g6387 ( 
.A1(n_5849),
.A2(n_5873),
.B(n_5927),
.Y(n_6387)
);

OAI21x1_ASAP7_75t_L g6388 ( 
.A1(n_5956),
.A2(n_3220),
.B(n_3214),
.Y(n_6388)
);

OAI21xp5_ASAP7_75t_L g6389 ( 
.A1(n_5979),
.A2(n_2426),
.B(n_2247),
.Y(n_6389)
);

OR2x2_ASAP7_75t_L g6390 ( 
.A(n_5801),
.B(n_52),
.Y(n_6390)
);

OAI21x1_ASAP7_75t_L g6391 ( 
.A1(n_5920),
.A2(n_2279),
.B(n_2234),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_5883),
.Y(n_6392)
);

OAI21x1_ASAP7_75t_L g6393 ( 
.A1(n_5957),
.A2(n_2279),
.B(n_2234),
.Y(n_6393)
);

AND2x2_ASAP7_75t_L g6394 ( 
.A(n_5998),
.B(n_53),
.Y(n_6394)
);

AOI21x1_ASAP7_75t_L g6395 ( 
.A1(n_6060),
.A2(n_1505),
.B(n_53),
.Y(n_6395)
);

OAI21x1_ASAP7_75t_L g6396 ( 
.A1(n_5982),
.A2(n_6071),
.B(n_5845),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_6007),
.Y(n_6397)
);

NOR2x1_ASAP7_75t_SL g6398 ( 
.A(n_6068),
.B(n_5976),
.Y(n_6398)
);

OAI21x1_ASAP7_75t_L g6399 ( 
.A1(n_5826),
.A2(n_2279),
.B(n_2234),
.Y(n_6399)
);

INVx2_ASAP7_75t_L g6400 ( 
.A(n_5791),
.Y(n_6400)
);

AOI22x1_ASAP7_75t_L g6401 ( 
.A1(n_6011),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_6401)
);

BUFx8_ASAP7_75t_L g6402 ( 
.A(n_6040),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_6007),
.Y(n_6403)
);

INVx2_ASAP7_75t_L g6404 ( 
.A(n_5791),
.Y(n_6404)
);

BUFx2_ASAP7_75t_SL g6405 ( 
.A(n_6103),
.Y(n_6405)
);

INVx5_ASAP7_75t_L g6406 ( 
.A(n_6047),
.Y(n_6406)
);

OAI21xp5_ASAP7_75t_L g6407 ( 
.A1(n_5810),
.A2(n_2426),
.B(n_2247),
.Y(n_6407)
);

AO21x1_ASAP7_75t_L g6408 ( 
.A1(n_5954),
.A2(n_54),
.B(n_56),
.Y(n_6408)
);

OAI21xp5_ASAP7_75t_L g6409 ( 
.A1(n_5851),
.A2(n_2247),
.B(n_2166),
.Y(n_6409)
);

BUFx3_ASAP7_75t_L g6410 ( 
.A(n_6103),
.Y(n_6410)
);

OR2x6_ASAP7_75t_L g6411 ( 
.A(n_6064),
.B(n_2466),
.Y(n_6411)
);

OAI21x1_ASAP7_75t_L g6412 ( 
.A1(n_5958),
.A2(n_2319),
.B(n_2187),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_6052),
.Y(n_6413)
);

AOI22x1_ASAP7_75t_L g6414 ( 
.A1(n_5872),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_6414)
);

INVx5_ASAP7_75t_L g6415 ( 
.A(n_5940),
.Y(n_6415)
);

BUFx12f_ASAP7_75t_L g6416 ( 
.A(n_6076),
.Y(n_6416)
);

OR2x2_ASAP7_75t_L g6417 ( 
.A(n_5784),
.B(n_60),
.Y(n_6417)
);

INVx3_ASAP7_75t_L g6418 ( 
.A(n_6061),
.Y(n_6418)
);

NAND2x1p5_ASAP7_75t_L g6419 ( 
.A(n_6109),
.B(n_2723),
.Y(n_6419)
);

INVx2_ASAP7_75t_SL g6420 ( 
.A(n_6024),
.Y(n_6420)
);

CKINVDCx20_ASAP7_75t_R g6421 ( 
.A(n_6088),
.Y(n_6421)
);

NAND2x1p5_ASAP7_75t_L g6422 ( 
.A(n_5964),
.B(n_2723),
.Y(n_6422)
);

INVx2_ASAP7_75t_SL g6423 ( 
.A(n_6025),
.Y(n_6423)
);

OAI21x1_ASAP7_75t_SL g6424 ( 
.A1(n_6053),
.A2(n_61),
.B(n_62),
.Y(n_6424)
);

BUFx3_ASAP7_75t_L g6425 ( 
.A(n_6035),
.Y(n_6425)
);

INVx3_ASAP7_75t_L g6426 ( 
.A(n_6113),
.Y(n_6426)
);

OAI21x1_ASAP7_75t_L g6427 ( 
.A1(n_5894),
.A2(n_6002),
.B(n_6066),
.Y(n_6427)
);

OAI21x1_ASAP7_75t_L g6428 ( 
.A1(n_5999),
.A2(n_2319),
.B(n_2187),
.Y(n_6428)
);

BUFx3_ASAP7_75t_L g6429 ( 
.A(n_6036),
.Y(n_6429)
);

BUFx3_ASAP7_75t_L g6430 ( 
.A(n_5906),
.Y(n_6430)
);

AO21x2_ASAP7_75t_L g6431 ( 
.A1(n_5876),
.A2(n_72),
.B(n_62),
.Y(n_6431)
);

AO21x2_ASAP7_75t_L g6432 ( 
.A1(n_5853),
.A2(n_73),
.B(n_63),
.Y(n_6432)
);

INVx3_ASAP7_75t_SL g6433 ( 
.A(n_6077),
.Y(n_6433)
);

INVx2_ASAP7_75t_L g6434 ( 
.A(n_6052),
.Y(n_6434)
);

AOI22xp33_ASAP7_75t_L g6435 ( 
.A1(n_6214),
.A2(n_6102),
.B1(n_5936),
.B2(n_5969),
.Y(n_6435)
);

CKINVDCx20_ASAP7_75t_R g6436 ( 
.A(n_6301),
.Y(n_6436)
);

BUFx6f_ASAP7_75t_L g6437 ( 
.A(n_6154),
.Y(n_6437)
);

OR2x6_ASAP7_75t_L g6438 ( 
.A(n_6304),
.B(n_5789),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6194),
.Y(n_6439)
);

AND2x4_ASAP7_75t_L g6440 ( 
.A(n_6173),
.B(n_6052),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6194),
.Y(n_6441)
);

NAND3xp33_ASAP7_75t_L g6442 ( 
.A(n_6270),
.B(n_5836),
.C(n_5963),
.Y(n_6442)
);

CKINVDCx20_ASAP7_75t_R g6443 ( 
.A(n_6301),
.Y(n_6443)
);

A2O1A1Ixp33_ASAP7_75t_L g6444 ( 
.A1(n_6270),
.A2(n_6214),
.B(n_6339),
.C(n_6282),
.Y(n_6444)
);

AND2x4_ASAP7_75t_L g6445 ( 
.A(n_6173),
.B(n_6028),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_6161),
.B(n_5787),
.Y(n_6446)
);

AO21x2_ASAP7_75t_L g6447 ( 
.A1(n_6153),
.A2(n_6137),
.B(n_6037),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_6142),
.Y(n_6448)
);

AND2x4_ASAP7_75t_L g6449 ( 
.A(n_6173),
.B(n_6108),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6144),
.Y(n_6450)
);

CKINVDCx5p33_ASAP7_75t_R g6451 ( 
.A(n_6239),
.Y(n_6451)
);

INVx2_ASAP7_75t_L g6452 ( 
.A(n_6162),
.Y(n_6452)
);

NAND2x1p5_ASAP7_75t_L g6453 ( 
.A(n_6319),
.B(n_6062),
.Y(n_6453)
);

A2O1A1Ixp33_ASAP7_75t_L g6454 ( 
.A1(n_6339),
.A2(n_6045),
.B(n_6057),
.C(n_6085),
.Y(n_6454)
);

INVx4_ASAP7_75t_L g6455 ( 
.A(n_6141),
.Y(n_6455)
);

NOR2xp33_ASAP7_75t_L g6456 ( 
.A(n_6201),
.B(n_6107),
.Y(n_6456)
);

OAI22xp5_ASAP7_75t_L g6457 ( 
.A1(n_6265),
.A2(n_6105),
.B1(n_5816),
.B2(n_6013),
.Y(n_6457)
);

NOR2x1_ASAP7_75t_SL g6458 ( 
.A(n_6162),
.B(n_5820),
.Y(n_6458)
);

OA21x2_ASAP7_75t_L g6459 ( 
.A1(n_6159),
.A2(n_5821),
.B(n_5852),
.Y(n_6459)
);

OAI21x1_ASAP7_75t_L g6460 ( 
.A1(n_6151),
.A2(n_6049),
.B(n_6006),
.Y(n_6460)
);

O2A1O1Ixp33_ASAP7_75t_SL g6461 ( 
.A1(n_6376),
.A2(n_5992),
.B(n_6000),
.C(n_6009),
.Y(n_6461)
);

NOR2xp67_ASAP7_75t_L g6462 ( 
.A(n_6173),
.B(n_5807),
.Y(n_6462)
);

AOI21x1_ASAP7_75t_L g6463 ( 
.A1(n_6167),
.A2(n_5949),
.B(n_5918),
.Y(n_6463)
);

INVx2_ASAP7_75t_L g6464 ( 
.A(n_6178),
.Y(n_6464)
);

OAI21x1_ASAP7_75t_L g6465 ( 
.A1(n_6243),
.A2(n_6202),
.B(n_6168),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6147),
.Y(n_6466)
);

OAI21x1_ASAP7_75t_L g6467 ( 
.A1(n_6139),
.A2(n_6029),
.B(n_5825),
.Y(n_6467)
);

INVx2_ASAP7_75t_SL g6468 ( 
.A(n_6141),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_6150),
.Y(n_6469)
);

NAND3xp33_ASAP7_75t_L g6470 ( 
.A(n_6402),
.B(n_6016),
.C(n_6094),
.Y(n_6470)
);

OAI21xp5_ASAP7_75t_L g6471 ( 
.A1(n_6145),
.A2(n_5926),
.B(n_5960),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_6309),
.B(n_5806),
.Y(n_6472)
);

AOI22xp33_ASAP7_75t_L g6473 ( 
.A1(n_6402),
.A2(n_5865),
.B1(n_6014),
.B2(n_6130),
.Y(n_6473)
);

OAI221xp5_ASAP7_75t_L g6474 ( 
.A1(n_6163),
.A2(n_5862),
.B1(n_5875),
.B2(n_5878),
.C(n_6003),
.Y(n_6474)
);

OAI21x1_ASAP7_75t_SL g6475 ( 
.A1(n_6398),
.A2(n_6048),
.B(n_6043),
.Y(n_6475)
);

OAI21x1_ASAP7_75t_L g6476 ( 
.A1(n_6139),
.A2(n_6122),
.B(n_6115),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6152),
.Y(n_6477)
);

BUFx6f_ASAP7_75t_L g6478 ( 
.A(n_6154),
.Y(n_6478)
);

OA21x2_ASAP7_75t_L g6479 ( 
.A1(n_6159),
.A2(n_6079),
.B(n_6065),
.Y(n_6479)
);

HB1xp67_ASAP7_75t_L g6480 ( 
.A(n_6261),
.Y(n_6480)
);

INVx6_ASAP7_75t_L g6481 ( 
.A(n_6171),
.Y(n_6481)
);

INVx8_ASAP7_75t_L g6482 ( 
.A(n_6141),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6161),
.B(n_5794),
.Y(n_6483)
);

AOI22xp33_ASAP7_75t_L g6484 ( 
.A1(n_6163),
.A2(n_6015),
.B1(n_5896),
.B2(n_6058),
.Y(n_6484)
);

INVx2_ASAP7_75t_L g6485 ( 
.A(n_6182),
.Y(n_6485)
);

AO32x2_ASAP7_75t_L g6486 ( 
.A1(n_6420),
.A2(n_5807),
.A3(n_5844),
.B1(n_6040),
.B2(n_5831),
.Y(n_6486)
);

OAI21x1_ASAP7_75t_L g6487 ( 
.A1(n_6170),
.A2(n_5977),
.B(n_5971),
.Y(n_6487)
);

NAND2x1p5_ASAP7_75t_L g6488 ( 
.A(n_6319),
.B(n_6213),
.Y(n_6488)
);

INVx1_ASAP7_75t_L g6489 ( 
.A(n_6166),
.Y(n_6489)
);

BUFx3_ASAP7_75t_L g6490 ( 
.A(n_6149),
.Y(n_6490)
);

INVx3_ASAP7_75t_L g6491 ( 
.A(n_6211),
.Y(n_6491)
);

OAI221xp5_ASAP7_75t_L g6492 ( 
.A1(n_6282),
.A2(n_6433),
.B1(n_6247),
.B2(n_6145),
.C(n_6265),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6303),
.B(n_6121),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_6191),
.Y(n_6494)
);

OA21x2_ASAP7_75t_L g6495 ( 
.A1(n_6400),
.A2(n_6086),
.B(n_6082),
.Y(n_6495)
);

NOR2x1_ASAP7_75t_SL g6496 ( 
.A(n_6181),
.B(n_5946),
.Y(n_6496)
);

AOI22xp33_ASAP7_75t_L g6497 ( 
.A1(n_6414),
.A2(n_6054),
.B1(n_5978),
.B2(n_6125),
.Y(n_6497)
);

INVx2_ASAP7_75t_L g6498 ( 
.A(n_6189),
.Y(n_6498)
);

OAI221xp5_ASAP7_75t_L g6499 ( 
.A1(n_6433),
.A2(n_5929),
.B1(n_5911),
.B2(n_5905),
.C(n_6124),
.Y(n_6499)
);

AND2x4_ASAP7_75t_L g6500 ( 
.A(n_6212),
.B(n_5881),
.Y(n_6500)
);

OAI21x1_ASAP7_75t_L g6501 ( 
.A1(n_6258),
.A2(n_6179),
.B(n_6193),
.Y(n_6501)
);

CKINVDCx5p33_ASAP7_75t_R g6502 ( 
.A(n_6239),
.Y(n_6502)
);

AOI22xp33_ASAP7_75t_L g6503 ( 
.A1(n_6415),
.A2(n_5815),
.B1(n_6001),
.B2(n_5922),
.Y(n_6503)
);

OAI22xp5_ASAP7_75t_L g6504 ( 
.A1(n_6233),
.A2(n_5937),
.B1(n_6127),
.B2(n_5834),
.Y(n_6504)
);

A2O1A1Ixp33_ASAP7_75t_L g6505 ( 
.A1(n_6415),
.A2(n_6376),
.B(n_6288),
.C(n_6195),
.Y(n_6505)
);

INVx1_ASAP7_75t_L g6506 ( 
.A(n_6192),
.Y(n_6506)
);

NAND2xp5_ASAP7_75t_L g6507 ( 
.A(n_6311),
.B(n_5794),
.Y(n_6507)
);

AND2x2_ASAP7_75t_L g6508 ( 
.A(n_6164),
.B(n_5794),
.Y(n_6508)
);

OAI21x1_ASAP7_75t_L g6509 ( 
.A1(n_6179),
.A2(n_5993),
.B(n_6059),
.Y(n_6509)
);

AOI222xp33_ASAP7_75t_L g6510 ( 
.A1(n_6415),
.A2(n_5962),
.B1(n_5868),
.B2(n_5961),
.C1(n_5942),
.C2(n_5935),
.Y(n_6510)
);

BUFx4f_ASAP7_75t_SL g6511 ( 
.A(n_6252),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6206),
.Y(n_6512)
);

AND2x2_ASAP7_75t_L g6513 ( 
.A(n_6164),
.B(n_5881),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_6209),
.Y(n_6514)
);

OAI21x1_ASAP7_75t_L g6515 ( 
.A1(n_6193),
.A2(n_6116),
.B(n_5833),
.Y(n_6515)
);

AO21x2_ASAP7_75t_L g6516 ( 
.A1(n_6153),
.A2(n_5907),
.B(n_5869),
.Y(n_6516)
);

OA21x2_ASAP7_75t_L g6517 ( 
.A1(n_6404),
.A2(n_5840),
.B(n_5913),
.Y(n_6517)
);

AND2x4_ASAP7_75t_L g6518 ( 
.A(n_6212),
.B(n_5881),
.Y(n_6518)
);

INVx2_ASAP7_75t_L g6519 ( 
.A(n_6197),
.Y(n_6519)
);

NOR2x1_ASAP7_75t_R g6520 ( 
.A(n_6230),
.B(n_5911),
.Y(n_6520)
);

AND2x2_ASAP7_75t_L g6521 ( 
.A(n_6272),
.B(n_5811),
.Y(n_6521)
);

HB1xp67_ASAP7_75t_L g6522 ( 
.A(n_6261),
.Y(n_6522)
);

OAI21x1_ASAP7_75t_L g6523 ( 
.A1(n_6336),
.A2(n_6392),
.B(n_6341),
.Y(n_6523)
);

OA21x2_ASAP7_75t_L g6524 ( 
.A1(n_6360),
.A2(n_6111),
.B(n_6090),
.Y(n_6524)
);

AO31x2_ASAP7_75t_L g6525 ( 
.A1(n_6314),
.A2(n_5838),
.A3(n_5824),
.B(n_5858),
.Y(n_6525)
);

NAND2xp5_ASAP7_75t_L g6526 ( 
.A(n_6278),
.B(n_5811),
.Y(n_6526)
);

AOI21xp5_ASAP7_75t_L g6527 ( 
.A1(n_6288),
.A2(n_6112),
.B(n_6104),
.Y(n_6527)
);

OAI221xp5_ASAP7_75t_L g6528 ( 
.A1(n_6174),
.A2(n_6148),
.B1(n_6224),
.B2(n_6307),
.C(n_6415),
.Y(n_6528)
);

A2O1A1Ixp33_ASAP7_75t_L g6529 ( 
.A1(n_6195),
.A2(n_5924),
.B(n_5990),
.C(n_6097),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6219),
.Y(n_6530)
);

INVx2_ASAP7_75t_L g6531 ( 
.A(n_6205),
.Y(n_6531)
);

AO22x2_ASAP7_75t_L g6532 ( 
.A1(n_6177),
.A2(n_6200),
.B1(n_6338),
.B2(n_6423),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_L g6533 ( 
.A(n_6374),
.B(n_5811),
.Y(n_6533)
);

OAI21x1_ASAP7_75t_L g6534 ( 
.A1(n_6386),
.A2(n_5839),
.B(n_6123),
.Y(n_6534)
);

AND2x4_ASAP7_75t_L g6535 ( 
.A(n_6143),
.B(n_6091),
.Y(n_6535)
);

O2A1O1Ixp33_ASAP7_75t_SL g6536 ( 
.A1(n_6185),
.A2(n_6040),
.B(n_5844),
.C(n_6131),
.Y(n_6536)
);

AND2x2_ASAP7_75t_L g6537 ( 
.A(n_6165),
.B(n_6177),
.Y(n_6537)
);

A2O1A1Ixp33_ASAP7_75t_L g6538 ( 
.A1(n_6342),
.A2(n_5844),
.B(n_6031),
.C(n_5994),
.Y(n_6538)
);

OR2x6_ASAP7_75t_L g6539 ( 
.A(n_6169),
.B(n_5832),
.Y(n_6539)
);

AOI22xp33_ASAP7_75t_SL g6540 ( 
.A1(n_6342),
.A2(n_6156),
.B1(n_6250),
.B2(n_6283),
.Y(n_6540)
);

AOI21xp5_ASAP7_75t_L g6541 ( 
.A1(n_6306),
.A2(n_5934),
.B(n_6018),
.Y(n_6541)
);

AND2x2_ASAP7_75t_L g6542 ( 
.A(n_6165),
.B(n_5859),
.Y(n_6542)
);

INVxp33_ASAP7_75t_SL g6543 ( 
.A(n_6160),
.Y(n_6543)
);

AND2x4_ASAP7_75t_L g6544 ( 
.A(n_6143),
.B(n_6155),
.Y(n_6544)
);

OR2x2_ASAP7_75t_L g6545 ( 
.A(n_6302),
.B(n_5859),
.Y(n_6545)
);

AO21x1_ASAP7_75t_L g6546 ( 
.A1(n_6284),
.A2(n_6096),
.B(n_6039),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_6215),
.Y(n_6547)
);

AO31x2_ASAP7_75t_L g6548 ( 
.A1(n_6408),
.A2(n_6135),
.A3(n_5859),
.B(n_65),
.Y(n_6548)
);

AND2x4_ASAP7_75t_L g6549 ( 
.A(n_6155),
.B(n_6033),
.Y(n_6549)
);

BUFx6f_ASAP7_75t_L g6550 ( 
.A(n_6154),
.Y(n_6550)
);

OAI21xp5_ASAP7_75t_L g6551 ( 
.A1(n_6264),
.A2(n_6026),
.B(n_5995),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_6374),
.B(n_6067),
.Y(n_6552)
);

OAI21x1_ASAP7_75t_L g6553 ( 
.A1(n_6386),
.A2(n_6396),
.B(n_6284),
.Y(n_6553)
);

BUFx2_ASAP7_75t_L g6554 ( 
.A(n_6252),
.Y(n_6554)
);

INVx2_ASAP7_75t_L g6555 ( 
.A(n_6222),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6223),
.Y(n_6556)
);

AOI22xp33_ASAP7_75t_L g6557 ( 
.A1(n_6250),
.A2(n_2466),
.B1(n_2383),
.B2(n_2392),
.Y(n_6557)
);

BUFx3_ASAP7_75t_L g6558 ( 
.A(n_6176),
.Y(n_6558)
);

NOR2xp33_ASAP7_75t_SL g6559 ( 
.A(n_6198),
.B(n_3862),
.Y(n_6559)
);

AO21x2_ASAP7_75t_L g6560 ( 
.A1(n_6140),
.A2(n_6078),
.B(n_63),
.Y(n_6560)
);

INVx2_ASAP7_75t_L g6561 ( 
.A(n_6236),
.Y(n_6561)
);

OAI21x1_ASAP7_75t_L g6562 ( 
.A1(n_6426),
.A2(n_2319),
.B(n_64),
.Y(n_6562)
);

OAI21x1_ASAP7_75t_L g6563 ( 
.A1(n_6426),
.A2(n_64),
.B(n_65),
.Y(n_6563)
);

BUFx2_ASAP7_75t_L g6564 ( 
.A(n_6241),
.Y(n_6564)
);

BUFx6f_ASAP7_75t_L g6565 ( 
.A(n_6172),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_6260),
.Y(n_6566)
);

OAI21x1_ASAP7_75t_L g6567 ( 
.A1(n_6418),
.A2(n_67),
.B(n_68),
.Y(n_6567)
);

INVx2_ASAP7_75t_L g6568 ( 
.A(n_6237),
.Y(n_6568)
);

OR2x4_ASAP7_75t_L g6569 ( 
.A(n_6417),
.B(n_67),
.Y(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_6257),
.B(n_70),
.Y(n_6570)
);

OAI21x1_ASAP7_75t_L g6571 ( 
.A1(n_6418),
.A2(n_70),
.B(n_71),
.Y(n_6571)
);

INVx2_ASAP7_75t_L g6572 ( 
.A(n_6237),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6228),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_6228),
.Y(n_6574)
);

AO31x2_ASAP7_75t_L g6575 ( 
.A1(n_6413),
.A2(n_73),
.A3(n_71),
.B(n_72),
.Y(n_6575)
);

NAND2xp5_ASAP7_75t_L g6576 ( 
.A(n_6257),
.B(n_75),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6299),
.Y(n_6577)
);

AOI21xp5_ASAP7_75t_L g6578 ( 
.A1(n_6306),
.A2(n_2383),
.B(n_2320),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6266),
.Y(n_6579)
);

NAND2xp5_ASAP7_75t_L g6580 ( 
.A(n_6332),
.B(n_6316),
.Y(n_6580)
);

INVx2_ASAP7_75t_L g6581 ( 
.A(n_6245),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6274),
.Y(n_6582)
);

AND2x4_ASAP7_75t_L g6583 ( 
.A(n_6406),
.B(n_75),
.Y(n_6583)
);

AO21x2_ASAP7_75t_L g6584 ( 
.A1(n_6140),
.A2(n_76),
.B(n_77),
.Y(n_6584)
);

INVx1_ASAP7_75t_L g6585 ( 
.A(n_6275),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_6289),
.Y(n_6586)
);

OAI21x1_ASAP7_75t_L g6587 ( 
.A1(n_6434),
.A2(n_77),
.B(n_78),
.Y(n_6587)
);

OAI22xp33_ASAP7_75t_L g6588 ( 
.A1(n_6203),
.A2(n_84),
.B1(n_78),
.B2(n_82),
.Y(n_6588)
);

NAND2x1p5_ASAP7_75t_L g6589 ( 
.A(n_6319),
.B(n_2723),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6255),
.Y(n_6590)
);

INVx1_ASAP7_75t_L g6591 ( 
.A(n_6138),
.Y(n_6591)
);

CKINVDCx5p33_ASAP7_75t_R g6592 ( 
.A(n_6160),
.Y(n_6592)
);

OAI21x1_ASAP7_75t_L g6593 ( 
.A1(n_6146),
.A2(n_82),
.B(n_85),
.Y(n_6593)
);

A2O1A1Ixp33_ASAP7_75t_L g6594 ( 
.A1(n_6224),
.A2(n_96),
.B(n_108),
.C(n_87),
.Y(n_6594)
);

NOR2xp33_ASAP7_75t_L g6595 ( 
.A(n_6198),
.B(n_88),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6157),
.Y(n_6596)
);

NOR2xp33_ASAP7_75t_L g6597 ( 
.A(n_6172),
.B(n_88),
.Y(n_6597)
);

AND2x4_ASAP7_75t_L g6598 ( 
.A(n_6406),
.B(n_89),
.Y(n_6598)
);

BUFx6f_ASAP7_75t_L g6599 ( 
.A(n_6169),
.Y(n_6599)
);

INVx2_ASAP7_75t_L g6600 ( 
.A(n_6255),
.Y(n_6600)
);

HB1xp67_ASAP7_75t_L g6601 ( 
.A(n_6180),
.Y(n_6601)
);

INVxp33_ASAP7_75t_L g6602 ( 
.A(n_6292),
.Y(n_6602)
);

OAI21x1_ASAP7_75t_SL g6603 ( 
.A1(n_6220),
.A2(n_89),
.B(n_90),
.Y(n_6603)
);

OAI21x1_ASAP7_75t_L g6604 ( 
.A1(n_6146),
.A2(n_6348),
.B(n_6329),
.Y(n_6604)
);

INVx1_ASAP7_75t_L g6605 ( 
.A(n_6231),
.Y(n_6605)
);

OA21x2_ASAP7_75t_L g6606 ( 
.A1(n_6318),
.A2(n_91),
.B(n_93),
.Y(n_6606)
);

AOI21x1_ASAP7_75t_L g6607 ( 
.A1(n_6240),
.A2(n_93),
.B(n_94),
.Y(n_6607)
);

INVx2_ASAP7_75t_L g6608 ( 
.A(n_6267),
.Y(n_6608)
);

NOR2xp33_ASAP7_75t_L g6609 ( 
.A(n_6185),
.B(n_95),
.Y(n_6609)
);

CKINVDCx6p67_ASAP7_75t_R g6610 ( 
.A(n_6169),
.Y(n_6610)
);

HB1xp67_ASAP7_75t_L g6611 ( 
.A(n_6180),
.Y(n_6611)
);

BUFx6f_ASAP7_75t_L g6612 ( 
.A(n_6188),
.Y(n_6612)
);

AO31x2_ASAP7_75t_L g6613 ( 
.A1(n_6335),
.A2(n_98),
.A3(n_95),
.B(n_97),
.Y(n_6613)
);

AOI21xp33_ASAP7_75t_L g6614 ( 
.A1(n_6240),
.A2(n_99),
.B(n_100),
.Y(n_6614)
);

AO31x2_ASAP7_75t_L g6615 ( 
.A1(n_6340),
.A2(n_105),
.A3(n_100),
.B(n_101),
.Y(n_6615)
);

BUFx6f_ASAP7_75t_L g6616 ( 
.A(n_6188),
.Y(n_6616)
);

NAND2xp5_ASAP7_75t_L g6617 ( 
.A(n_6316),
.B(n_101),
.Y(n_6617)
);

HB1xp67_ASAP7_75t_L g6618 ( 
.A(n_6235),
.Y(n_6618)
);

OA21x2_ASAP7_75t_L g6619 ( 
.A1(n_6344),
.A2(n_105),
.B(n_107),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6254),
.Y(n_6620)
);

AO31x2_ASAP7_75t_L g6621 ( 
.A1(n_6350),
.A2(n_110),
.A3(n_107),
.B(n_109),
.Y(n_6621)
);

NAND3xp33_ASAP7_75t_L g6622 ( 
.A(n_6190),
.B(n_2383),
.C(n_2320),
.Y(n_6622)
);

OAI21x1_ASAP7_75t_L g6623 ( 
.A1(n_6329),
.A2(n_110),
.B(n_112),
.Y(n_6623)
);

OAI21x1_ASAP7_75t_L g6624 ( 
.A1(n_6348),
.A2(n_113),
.B(n_114),
.Y(n_6624)
);

AOI22xp33_ASAP7_75t_L g6625 ( 
.A1(n_6283),
.A2(n_2383),
.B1(n_2392),
.B2(n_2320),
.Y(n_6625)
);

OAI21x1_ASAP7_75t_L g6626 ( 
.A1(n_6385),
.A2(n_116),
.B(n_117),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6262),
.Y(n_6627)
);

OAI221xp5_ASAP7_75t_L g6628 ( 
.A1(n_6174),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.C(n_119),
.Y(n_6628)
);

OAI21x1_ASAP7_75t_L g6629 ( 
.A1(n_6322),
.A2(n_118),
.B(n_120),
.Y(n_6629)
);

NAND2xp5_ASAP7_75t_L g6630 ( 
.A(n_6364),
.B(n_120),
.Y(n_6630)
);

OAI21x1_ASAP7_75t_L g6631 ( 
.A1(n_6372),
.A2(n_123),
.B(n_124),
.Y(n_6631)
);

AOI21x1_ASAP7_75t_L g6632 ( 
.A1(n_6394),
.A2(n_123),
.B(n_125),
.Y(n_6632)
);

OAI21xp5_ASAP7_75t_L g6633 ( 
.A1(n_6321),
.A2(n_126),
.B(n_127),
.Y(n_6633)
);

OAI22xp5_ASAP7_75t_L g6634 ( 
.A1(n_6233),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6273),
.Y(n_6635)
);

BUFx6f_ASAP7_75t_L g6636 ( 
.A(n_6188),
.Y(n_6636)
);

AOI21xp5_ASAP7_75t_L g6637 ( 
.A1(n_6321),
.A2(n_2392),
.B(n_2320),
.Y(n_6637)
);

OAI21x1_ASAP7_75t_L g6638 ( 
.A1(n_6397),
.A2(n_128),
.B(n_129),
.Y(n_6638)
);

A2O1A1Ixp33_ASAP7_75t_L g6639 ( 
.A1(n_6389),
.A2(n_142),
.B(n_151),
.C(n_130),
.Y(n_6639)
);

OAI21x1_ASAP7_75t_L g6640 ( 
.A1(n_6403),
.A2(n_131),
.B(n_132),
.Y(n_6640)
);

OAI21x1_ASAP7_75t_L g6641 ( 
.A1(n_6268),
.A2(n_132),
.B(n_134),
.Y(n_6641)
);

INVx2_ASAP7_75t_SL g6642 ( 
.A(n_6184),
.Y(n_6642)
);

OAI22xp33_ASAP7_75t_L g6643 ( 
.A1(n_6203),
.A2(n_138),
.B1(n_134),
.B2(n_137),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_6364),
.Y(n_6644)
);

AO21x2_ASAP7_75t_L g6645 ( 
.A1(n_6287),
.A2(n_138),
.B(n_139),
.Y(n_6645)
);

OAI22xp5_ASAP7_75t_L g6646 ( 
.A1(n_6203),
.A2(n_144),
.B1(n_140),
.B2(n_143),
.Y(n_6646)
);

OAI22xp5_ASAP7_75t_SL g6647 ( 
.A1(n_6308),
.A2(n_145),
.B1(n_140),
.B2(n_144),
.Y(n_6647)
);

AND2x4_ASAP7_75t_L g6648 ( 
.A(n_6406),
.B(n_145),
.Y(n_6648)
);

OAI21x1_ASAP7_75t_L g6649 ( 
.A1(n_6427),
.A2(n_146),
.B(n_147),
.Y(n_6649)
);

OAI21x1_ASAP7_75t_L g6650 ( 
.A1(n_6323),
.A2(n_146),
.B(n_147),
.Y(n_6650)
);

OAI211xp5_ASAP7_75t_SL g6651 ( 
.A1(n_6390),
.A2(n_152),
.B(n_148),
.C(n_149),
.Y(n_6651)
);

AOI21x1_ASAP7_75t_L g6652 ( 
.A1(n_6287),
.A2(n_152),
.B(n_153),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_6327),
.Y(n_6653)
);

BUFx6f_ASAP7_75t_L g6654 ( 
.A(n_6207),
.Y(n_6654)
);

AND2x4_ASAP7_75t_L g6655 ( 
.A(n_6406),
.B(n_154),
.Y(n_6655)
);

AO21x1_ASAP7_75t_L g6656 ( 
.A1(n_6211),
.A2(n_154),
.B(n_155),
.Y(n_6656)
);

OAI21x1_ASAP7_75t_L g6657 ( 
.A1(n_6277),
.A2(n_6267),
.B(n_6190),
.Y(n_6657)
);

INVx3_ASAP7_75t_L g6658 ( 
.A(n_6286),
.Y(n_6658)
);

OAI21x1_ASAP7_75t_L g6659 ( 
.A1(n_6276),
.A2(n_155),
.B(n_156),
.Y(n_6659)
);

AO21x2_ASAP7_75t_L g6660 ( 
.A1(n_6158),
.A2(n_157),
.B(n_159),
.Y(n_6660)
);

NAND2x1p5_ASAP7_75t_L g6661 ( 
.A(n_6319),
.B(n_2733),
.Y(n_6661)
);

HB1xp67_ASAP7_75t_L g6662 ( 
.A(n_6229),
.Y(n_6662)
);

OAI21x1_ASAP7_75t_L g6663 ( 
.A1(n_6204),
.A2(n_157),
.B(n_160),
.Y(n_6663)
);

OR2x6_ASAP7_75t_L g6664 ( 
.A(n_6286),
.B(n_2733),
.Y(n_6664)
);

AOI22xp33_ASAP7_75t_L g6665 ( 
.A1(n_6305),
.A2(n_2408),
.B1(n_2413),
.B2(n_2392),
.Y(n_6665)
);

AOI21x1_ASAP7_75t_L g6666 ( 
.A1(n_6295),
.A2(n_161),
.B(n_162),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_6186),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_6317),
.Y(n_6668)
);

OAI21x1_ASAP7_75t_L g6669 ( 
.A1(n_6204),
.A2(n_162),
.B(n_163),
.Y(n_6669)
);

HB1xp67_ASAP7_75t_L g6670 ( 
.A(n_6229),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_6227),
.Y(n_6671)
);

BUFx6f_ASAP7_75t_L g6672 ( 
.A(n_6207),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6320),
.Y(n_6673)
);

HB1xp67_ASAP7_75t_L g6674 ( 
.A(n_6345),
.Y(n_6674)
);

AOI21xp5_ASAP7_75t_L g6675 ( 
.A1(n_6325),
.A2(n_2413),
.B(n_2408),
.Y(n_6675)
);

OAI21x1_ASAP7_75t_L g6676 ( 
.A1(n_6226),
.A2(n_164),
.B(n_165),
.Y(n_6676)
);

OAI21x1_ASAP7_75t_L g6677 ( 
.A1(n_6226),
.A2(n_6320),
.B(n_6290),
.Y(n_6677)
);

OAI21x1_ASAP7_75t_L g6678 ( 
.A1(n_6387),
.A2(n_6328),
.B(n_6379),
.Y(n_6678)
);

BUFx2_ASAP7_75t_L g6679 ( 
.A(n_6256),
.Y(n_6679)
);

INVx2_ASAP7_75t_L g6680 ( 
.A(n_6300),
.Y(n_6680)
);

INVx2_ASAP7_75t_L g6681 ( 
.A(n_6300),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6300),
.Y(n_6682)
);

CKINVDCx5p33_ASAP7_75t_R g6683 ( 
.A(n_6183),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6369),
.Y(n_6684)
);

BUFx2_ASAP7_75t_L g6685 ( 
.A(n_6256),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6242),
.B(n_164),
.Y(n_6686)
);

NAND2x1p5_ASAP7_75t_L g6687 ( 
.A(n_6213),
.B(n_2733),
.Y(n_6687)
);

HB1xp67_ASAP7_75t_L g6688 ( 
.A(n_6345),
.Y(n_6688)
);

BUFx12f_ASAP7_75t_L g6689 ( 
.A(n_6362),
.Y(n_6689)
);

NOR2xp67_ASAP7_75t_L g6690 ( 
.A(n_6281),
.B(n_166),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6369),
.Y(n_6691)
);

OAI21xp5_ASAP7_75t_L g6692 ( 
.A1(n_6292),
.A2(n_166),
.B(n_167),
.Y(n_6692)
);

OA21x2_ASAP7_75t_L g6693 ( 
.A1(n_6501),
.A2(n_6325),
.B(n_6379),
.Y(n_6693)
);

INVx1_ASAP7_75t_L g6694 ( 
.A(n_6448),
.Y(n_6694)
);

AO21x2_ASAP7_75t_L g6695 ( 
.A1(n_6607),
.A2(n_6158),
.B(n_6431),
.Y(n_6695)
);

NAND2x1p5_ASAP7_75t_L g6696 ( 
.A(n_6449),
.B(n_6213),
.Y(n_6696)
);

INVxp33_ASAP7_75t_L g6697 ( 
.A(n_6520),
.Y(n_6697)
);

OAI21xp5_ASAP7_75t_L g6698 ( 
.A1(n_6444),
.A2(n_6174),
.B(n_6395),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_6450),
.Y(n_6699)
);

AO21x2_ASAP7_75t_L g6700 ( 
.A1(n_6607),
.A2(n_6614),
.B(n_6458),
.Y(n_6700)
);

A2O1A1Ixp33_ASAP7_75t_L g6701 ( 
.A1(n_6505),
.A2(n_6389),
.B(n_6430),
.C(n_6378),
.Y(n_6701)
);

OAI21x1_ASAP7_75t_L g6702 ( 
.A1(n_6604),
.A2(n_6553),
.B(n_6465),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6466),
.Y(n_6703)
);

OAI21x1_ASAP7_75t_L g6704 ( 
.A1(n_6657),
.A2(n_6281),
.B(n_6334),
.Y(n_6704)
);

OA21x2_ASAP7_75t_L g6705 ( 
.A1(n_6452),
.A2(n_6175),
.B(n_6351),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6469),
.Y(n_6706)
);

OA21x2_ASAP7_75t_L g6707 ( 
.A1(n_6523),
.A2(n_6351),
.B(n_6352),
.Y(n_6707)
);

OAI21x1_ASAP7_75t_L g6708 ( 
.A1(n_6488),
.A2(n_6347),
.B(n_6334),
.Y(n_6708)
);

OAI21xp5_ASAP7_75t_L g6709 ( 
.A1(n_6540),
.A2(n_6378),
.B(n_6401),
.Y(n_6709)
);

A2O1A1Ixp33_ASAP7_75t_L g6710 ( 
.A1(n_6609),
.A2(n_6492),
.B(n_6454),
.C(n_6470),
.Y(n_6710)
);

NAND2xp5_ASAP7_75t_L g6711 ( 
.A(n_6447),
.B(n_6425),
.Y(n_6711)
);

INVx2_ASAP7_75t_L g6712 ( 
.A(n_6612),
.Y(n_6712)
);

AND2x2_ASAP7_75t_SL g6713 ( 
.A(n_6674),
.B(n_6326),
.Y(n_6713)
);

AOI21xp5_ASAP7_75t_L g6714 ( 
.A1(n_6461),
.A2(n_6536),
.B(n_6438),
.Y(n_6714)
);

OA21x2_ASAP7_75t_L g6715 ( 
.A1(n_6507),
.A2(n_6393),
.B(n_6391),
.Y(n_6715)
);

BUFx2_ASAP7_75t_SL g6716 ( 
.A(n_6436),
.Y(n_6716)
);

BUFx3_ASAP7_75t_L g6717 ( 
.A(n_6443),
.Y(n_6717)
);

NAND2xp5_ASAP7_75t_SL g6718 ( 
.A(n_6463),
.B(n_6187),
.Y(n_6718)
);

AO31x2_ASAP7_75t_L g6719 ( 
.A1(n_6458),
.A2(n_6333),
.A3(n_6368),
.B(n_6431),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6477),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6489),
.Y(n_6721)
);

AND2x2_ASAP7_75t_L g6722 ( 
.A(n_6537),
.B(n_6269),
.Y(n_6722)
);

OAI21x1_ASAP7_75t_L g6723 ( 
.A1(n_6677),
.A2(n_6347),
.B(n_6353),
.Y(n_6723)
);

AOI21x1_ASAP7_75t_L g6724 ( 
.A1(n_6554),
.A2(n_6564),
.B(n_6688),
.Y(n_6724)
);

OAI21x1_ASAP7_75t_SL g6725 ( 
.A1(n_6463),
.A2(n_6424),
.B(n_6253),
.Y(n_6725)
);

INVx1_ASAP7_75t_L g6726 ( 
.A(n_6494),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6506),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_6667),
.B(n_6495),
.Y(n_6728)
);

AOI21xp5_ASAP7_75t_L g6729 ( 
.A1(n_6438),
.A2(n_6232),
.B(n_6234),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6512),
.Y(n_6730)
);

AND2x4_ASAP7_75t_L g6731 ( 
.A(n_6491),
.B(n_6213),
.Y(n_6731)
);

AOI22xp5_ASAP7_75t_L g6732 ( 
.A1(n_6634),
.A2(n_6232),
.B1(n_6246),
.B2(n_6371),
.Y(n_6732)
);

AOI21x1_ASAP7_75t_L g6733 ( 
.A1(n_6532),
.A2(n_6652),
.B(n_6611),
.Y(n_6733)
);

NAND2x1p5_ASAP7_75t_L g6734 ( 
.A(n_6449),
.B(n_6238),
.Y(n_6734)
);

BUFx6f_ASAP7_75t_L g6735 ( 
.A(n_6490),
.Y(n_6735)
);

AO31x2_ASAP7_75t_L g6736 ( 
.A1(n_6546),
.A2(n_6333),
.A3(n_6368),
.B(n_6432),
.Y(n_6736)
);

AO31x2_ASAP7_75t_L g6737 ( 
.A1(n_6656),
.A2(n_6432),
.A3(n_6196),
.B(n_6363),
.Y(n_6737)
);

BUFx12f_ASAP7_75t_L g6738 ( 
.A(n_6451),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_6514),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6530),
.Y(n_6740)
);

A2O1A1Ixp33_ASAP7_75t_L g6741 ( 
.A1(n_6594),
.A2(n_6429),
.B(n_6383),
.C(n_6234),
.Y(n_6741)
);

AO21x2_ASAP7_75t_L g6742 ( 
.A1(n_6601),
.A2(n_6584),
.B(n_6622),
.Y(n_6742)
);

OAI21x1_ASAP7_75t_L g6743 ( 
.A1(n_6593),
.A2(n_6353),
.B(n_6422),
.Y(n_6743)
);

INVxp33_ASAP7_75t_L g6744 ( 
.A(n_6595),
.Y(n_6744)
);

AOI22xp33_ASAP7_75t_L g6745 ( 
.A1(n_6442),
.A2(n_6346),
.B1(n_6218),
.B2(n_6246),
.Y(n_6745)
);

INVx3_ASAP7_75t_L g6746 ( 
.A(n_6565),
.Y(n_6746)
);

BUFx2_ASAP7_75t_L g6747 ( 
.A(n_6532),
.Y(n_6747)
);

OR2x2_ASAP7_75t_L g6748 ( 
.A(n_6479),
.B(n_6218),
.Y(n_6748)
);

INVx2_ASAP7_75t_L g6749 ( 
.A(n_6612),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_L g6750 ( 
.A(n_6495),
.B(n_6218),
.Y(n_6750)
);

AND2x2_ASAP7_75t_L g6751 ( 
.A(n_6679),
.B(n_6269),
.Y(n_6751)
);

BUFx4f_ASAP7_75t_SL g6752 ( 
.A(n_6689),
.Y(n_6752)
);

AO21x2_ASAP7_75t_L g6753 ( 
.A1(n_6660),
.A2(n_6251),
.B(n_6242),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6612),
.Y(n_6754)
);

OAI21x1_ASAP7_75t_L g6755 ( 
.A1(n_6526),
.A2(n_6422),
.B(n_6355),
.Y(n_6755)
);

A2O1A1Ixp33_ASAP7_75t_L g6756 ( 
.A1(n_6538),
.A2(n_6383),
.B(n_6330),
.C(n_6234),
.Y(n_6756)
);

OA21x2_ASAP7_75t_L g6757 ( 
.A1(n_6533),
.A2(n_6279),
.B(n_6297),
.Y(n_6757)
);

INVx2_ASAP7_75t_L g6758 ( 
.A(n_6616),
.Y(n_6758)
);

AOI21xp5_ASAP7_75t_L g6759 ( 
.A1(n_6474),
.A2(n_6330),
.B(n_6246),
.Y(n_6759)
);

NAND2xp5_ASAP7_75t_L g6760 ( 
.A(n_6471),
.B(n_6421),
.Y(n_6760)
);

AO21x2_ASAP7_75t_L g6761 ( 
.A1(n_6652),
.A2(n_6251),
.B(n_6293),
.Y(n_6761)
);

A2O1A1Ixp33_ASAP7_75t_L g6762 ( 
.A1(n_6528),
.A2(n_6330),
.B(n_6409),
.C(n_6421),
.Y(n_6762)
);

AO31x2_ASAP7_75t_L g6763 ( 
.A1(n_6685),
.A2(n_6196),
.A3(n_6359),
.B(n_6296),
.Y(n_6763)
);

OAI21xp5_ASAP7_75t_L g6764 ( 
.A1(n_6435),
.A2(n_6308),
.B(n_6409),
.Y(n_6764)
);

NAND2xp5_ASAP7_75t_L g6765 ( 
.A(n_6479),
.B(n_6225),
.Y(n_6765)
);

AO31x2_ASAP7_75t_L g6766 ( 
.A1(n_6630),
.A2(n_6359),
.A3(n_6361),
.B(n_6296),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6653),
.B(n_6217),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6616),
.Y(n_6768)
);

NAND2xp5_ASAP7_75t_L g6769 ( 
.A(n_6493),
.B(n_6249),
.Y(n_6769)
);

NOR2xp67_ASAP7_75t_L g6770 ( 
.A(n_6491),
.B(n_6238),
.Y(n_6770)
);

OAI21x1_ASAP7_75t_L g6771 ( 
.A1(n_6476),
.A2(n_6355),
.B(n_6354),
.Y(n_6771)
);

INVx3_ASAP7_75t_L g6772 ( 
.A(n_6565),
.Y(n_6772)
);

INVx2_ASAP7_75t_SL g6773 ( 
.A(n_6481),
.Y(n_6773)
);

AOI21xp5_ASAP7_75t_L g6774 ( 
.A1(n_6510),
.A2(n_6210),
.B(n_6315),
.Y(n_6774)
);

AO31x2_ASAP7_75t_L g6775 ( 
.A1(n_6680),
.A2(n_6361),
.A3(n_6207),
.B(n_6221),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6556),
.Y(n_6776)
);

OAI21x1_ASAP7_75t_L g6777 ( 
.A1(n_6515),
.A2(n_6419),
.B(n_6412),
.Y(n_6777)
);

INVx2_ASAP7_75t_L g6778 ( 
.A(n_6616),
.Y(n_6778)
);

AO31x2_ASAP7_75t_L g6779 ( 
.A1(n_6496),
.A2(n_6221),
.A3(n_6216),
.B(n_6244),
.Y(n_6779)
);

A2O1A1Ixp33_ASAP7_75t_L g6780 ( 
.A1(n_6692),
.A2(n_6238),
.B(n_6199),
.C(n_6407),
.Y(n_6780)
);

NOR2xp33_ASAP7_75t_L g6781 ( 
.A(n_6543),
.B(n_6248),
.Y(n_6781)
);

AOI21x1_ASAP7_75t_L g6782 ( 
.A1(n_6632),
.A2(n_6411),
.B(n_6293),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6566),
.Y(n_6783)
);

OAI21x1_ASAP7_75t_L g6784 ( 
.A1(n_6453),
.A2(n_6419),
.B(n_6382),
.Y(n_6784)
);

INVx2_ASAP7_75t_L g6785 ( 
.A(n_6636),
.Y(n_6785)
);

OR2x2_ASAP7_75t_L g6786 ( 
.A(n_6580),
.B(n_6313),
.Y(n_6786)
);

AO21x2_ASAP7_75t_L g6787 ( 
.A1(n_6645),
.A2(n_6210),
.B(n_6399),
.Y(n_6787)
);

A2O1A1Ixp33_ASAP7_75t_L g6788 ( 
.A1(n_6628),
.A2(n_6238),
.B(n_6407),
.C(n_6294),
.Y(n_6788)
);

OAI21x1_ASAP7_75t_L g6789 ( 
.A1(n_6460),
.A2(n_6382),
.B(n_6357),
.Y(n_6789)
);

OAI21xp5_ASAP7_75t_L g6790 ( 
.A1(n_6504),
.A2(n_6315),
.B(n_6263),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6577),
.Y(n_6791)
);

OR2x2_ASAP7_75t_L g6792 ( 
.A(n_6573),
.B(n_6313),
.Y(n_6792)
);

AOI21xp5_ASAP7_75t_L g6793 ( 
.A1(n_6503),
.A2(n_6411),
.B(n_6263),
.Y(n_6793)
);

OA21x2_ASAP7_75t_L g6794 ( 
.A1(n_6439),
.A2(n_6343),
.B(n_6428),
.Y(n_6794)
);

AOI21xp5_ASAP7_75t_L g6795 ( 
.A1(n_6529),
.A2(n_6411),
.B(n_6294),
.Y(n_6795)
);

INVx2_ASAP7_75t_L g6796 ( 
.A(n_6636),
.Y(n_6796)
);

AOI21xp5_ASAP7_75t_L g6797 ( 
.A1(n_6457),
.A2(n_6331),
.B(n_6208),
.Y(n_6797)
);

NAND2x1p5_ASAP7_75t_L g6798 ( 
.A(n_6583),
.B(n_6259),
.Y(n_6798)
);

NAND2xp5_ASAP7_75t_L g6799 ( 
.A(n_6472),
.B(n_6271),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6555),
.Y(n_6800)
);

AOI221xp5_ASAP7_75t_SL g6801 ( 
.A1(n_6647),
.A2(n_6221),
.B1(n_6216),
.B2(n_6405),
.C(n_6310),
.Y(n_6801)
);

AO21x2_ASAP7_75t_L g6802 ( 
.A1(n_6475),
.A2(n_6331),
.B(n_6291),
.Y(n_6802)
);

NAND2xp5_ASAP7_75t_L g6803 ( 
.A(n_6445),
.B(n_6358),
.Y(n_6803)
);

NAND2xp5_ASAP7_75t_L g6804 ( 
.A(n_6445),
.B(n_6216),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_L g6805 ( 
.A(n_6574),
.B(n_6337),
.Y(n_6805)
);

OA21x2_ASAP7_75t_L g6806 ( 
.A1(n_6441),
.A2(n_6367),
.B(n_6366),
.Y(n_6806)
);

OA21x2_ASAP7_75t_L g6807 ( 
.A1(n_6644),
.A2(n_6388),
.B(n_6365),
.Y(n_6807)
);

INVx3_ASAP7_75t_L g6808 ( 
.A(n_6565),
.Y(n_6808)
);

BUFx6f_ASAP7_75t_L g6809 ( 
.A(n_6437),
.Y(n_6809)
);

AND2x4_ASAP7_75t_L g6810 ( 
.A(n_6658),
.B(n_6410),
.Y(n_6810)
);

OR2x2_ASAP7_75t_L g6811 ( 
.A(n_6552),
.B(n_6291),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6561),
.Y(n_6812)
);

OAI21x1_ASAP7_75t_L g6813 ( 
.A1(n_6590),
.A2(n_6373),
.B(n_6370),
.Y(n_6813)
);

NAND2xp5_ASAP7_75t_L g6814 ( 
.A(n_6617),
.B(n_6356),
.Y(n_6814)
);

AND2x4_ASAP7_75t_L g6815 ( 
.A(n_6658),
.B(n_6375),
.Y(n_6815)
);

AOI21xp5_ASAP7_75t_L g6816 ( 
.A1(n_6633),
.A2(n_6370),
.B(n_6285),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6570),
.B(n_6380),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_6579),
.Y(n_6818)
);

BUFx3_ASAP7_75t_L g6819 ( 
.A(n_6502),
.Y(n_6819)
);

INVx2_ASAP7_75t_L g6820 ( 
.A(n_6636),
.Y(n_6820)
);

AOI21xp5_ASAP7_75t_L g6821 ( 
.A1(n_6484),
.A2(n_6285),
.B(n_6280),
.Y(n_6821)
);

INVx1_ASAP7_75t_L g6822 ( 
.A(n_6582),
.Y(n_6822)
);

AO31x2_ASAP7_75t_L g6823 ( 
.A1(n_6496),
.A2(n_6310),
.A3(n_6312),
.B(n_6244),
.Y(n_6823)
);

NAND2xp5_ASAP7_75t_SL g6824 ( 
.A(n_6475),
.B(n_6324),
.Y(n_6824)
);

INVx2_ASAP7_75t_SL g6825 ( 
.A(n_6481),
.Y(n_6825)
);

OR2x2_ASAP7_75t_L g6826 ( 
.A(n_6671),
.B(n_6381),
.Y(n_6826)
);

AND2x2_ASAP7_75t_L g6827 ( 
.A(n_6446),
.B(n_6381),
.Y(n_6827)
);

AOI21x1_ASAP7_75t_L g6828 ( 
.A1(n_6632),
.A2(n_6324),
.B(n_6310),
.Y(n_6828)
);

OR2x2_ASAP7_75t_L g6829 ( 
.A(n_6516),
.B(n_6381),
.Y(n_6829)
);

INVx3_ASAP7_75t_L g6830 ( 
.A(n_6437),
.Y(n_6830)
);

AND2x2_ASAP7_75t_L g6831 ( 
.A(n_6602),
.B(n_6244),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6585),
.Y(n_6832)
);

OAI21xp5_ASAP7_75t_L g6833 ( 
.A1(n_6690),
.A2(n_6324),
.B(n_6416),
.Y(n_6833)
);

OA21x2_ASAP7_75t_L g6834 ( 
.A1(n_6483),
.A2(n_6324),
.B(n_6312),
.Y(n_6834)
);

OAI21xp5_ASAP7_75t_L g6835 ( 
.A1(n_6639),
.A2(n_6324),
.B(n_6312),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_L g6836 ( 
.A(n_6576),
.B(n_6349),
.Y(n_6836)
);

HB1xp67_ASAP7_75t_L g6837 ( 
.A(n_6480),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6681),
.B(n_6349),
.Y(n_6838)
);

NAND2xp5_ASAP7_75t_L g6839 ( 
.A(n_6682),
.B(n_6586),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_6522),
.Y(n_6840)
);

AND2x4_ASAP7_75t_L g6841 ( 
.A(n_6544),
.B(n_6349),
.Y(n_6841)
);

NAND2x1p5_ASAP7_75t_L g6842 ( 
.A(n_6583),
.B(n_6280),
.Y(n_6842)
);

NAND2xp5_ASAP7_75t_L g6843 ( 
.A(n_6618),
.B(n_6591),
.Y(n_6843)
);

OA21x2_ASAP7_75t_L g6844 ( 
.A1(n_6508),
.A2(n_6377),
.B(n_6384),
.Y(n_6844)
);

AOI21xp5_ASAP7_75t_L g6845 ( 
.A1(n_6499),
.A2(n_6377),
.B(n_6298),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_6606),
.Y(n_6846)
);

A2O1A1Ixp33_ASAP7_75t_L g6847 ( 
.A1(n_6651),
.A2(n_170),
.B(n_167),
.C(n_169),
.Y(n_6847)
);

AOI21xp5_ASAP7_75t_L g6848 ( 
.A1(n_6588),
.A2(n_6298),
.B(n_6384),
.Y(n_6848)
);

OR2x2_ASAP7_75t_L g6849 ( 
.A(n_6581),
.B(n_170),
.Y(n_6849)
);

INVx1_ASAP7_75t_L g6850 ( 
.A(n_6606),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_6619),
.Y(n_6851)
);

AOI21xp5_ASAP7_75t_L g6852 ( 
.A1(n_6643),
.A2(n_171),
.B(n_173),
.Y(n_6852)
);

NAND2xp5_ASAP7_75t_L g6853 ( 
.A(n_6596),
.B(n_175),
.Y(n_6853)
);

NAND2x1p5_ASAP7_75t_L g6854 ( 
.A(n_6598),
.B(n_2745),
.Y(n_6854)
);

HB1xp67_ASAP7_75t_L g6855 ( 
.A(n_6662),
.Y(n_6855)
);

INVx6_ASAP7_75t_L g6856 ( 
.A(n_6482),
.Y(n_6856)
);

OAI21x1_ASAP7_75t_SL g6857 ( 
.A1(n_6603),
.A2(n_176),
.B(n_177),
.Y(n_6857)
);

AOI21xp5_ASAP7_75t_L g6858 ( 
.A1(n_6646),
.A2(n_178),
.B(n_179),
.Y(n_6858)
);

INVx2_ASAP7_75t_L g6859 ( 
.A(n_6654),
.Y(n_6859)
);

NAND2xp5_ASAP7_75t_L g6860 ( 
.A(n_6605),
.B(n_6620),
.Y(n_6860)
);

NOR2xp33_ASAP7_75t_L g6861 ( 
.A(n_6455),
.B(n_178),
.Y(n_6861)
);

OAI21x1_ASAP7_75t_L g6862 ( 
.A1(n_6600),
.A2(n_6608),
.B(n_6673),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_L g6863 ( 
.A(n_6627),
.B(n_179),
.Y(n_6863)
);

NOR2xp33_ASAP7_75t_L g6864 ( 
.A(n_6455),
.B(n_6511),
.Y(n_6864)
);

A2O1A1Ixp33_ASAP7_75t_L g6865 ( 
.A1(n_6597),
.A2(n_183),
.B(n_180),
.C(n_182),
.Y(n_6865)
);

AO31x2_ASAP7_75t_L g6866 ( 
.A1(n_6456),
.A2(n_186),
.A3(n_182),
.B(n_185),
.Y(n_6866)
);

NAND2xp5_ASAP7_75t_L g6867 ( 
.A(n_6635),
.B(n_188),
.Y(n_6867)
);

NAND2xp5_ASAP7_75t_L g6868 ( 
.A(n_6670),
.B(n_188),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_L g6869 ( 
.A(n_6668),
.B(n_189),
.Y(n_6869)
);

OAI21x1_ASAP7_75t_L g6870 ( 
.A1(n_6513),
.A2(n_6572),
.B(n_6568),
.Y(n_6870)
);

AOI21xp5_ASAP7_75t_L g6871 ( 
.A1(n_6527),
.A2(n_190),
.B(n_191),
.Y(n_6871)
);

AND2x2_ASAP7_75t_L g6872 ( 
.A(n_6544),
.B(n_190),
.Y(n_6872)
);

INVx2_ASAP7_75t_L g6873 ( 
.A(n_6654),
.Y(n_6873)
);

OR2x2_ASAP7_75t_L g6874 ( 
.A(n_6545),
.B(n_193),
.Y(n_6874)
);

NAND2xp5_ASAP7_75t_SL g6875 ( 
.A(n_6599),
.B(n_2408),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_6619),
.Y(n_6876)
);

OAI21x1_ASAP7_75t_L g6877 ( 
.A1(n_6509),
.A2(n_194),
.B(n_195),
.Y(n_6877)
);

CKINVDCx8_ASAP7_75t_R g6878 ( 
.A(n_6592),
.Y(n_6878)
);

NAND2xp5_ASAP7_75t_L g6879 ( 
.A(n_6642),
.B(n_194),
.Y(n_6879)
);

OAI21xp5_ASAP7_75t_L g6880 ( 
.A1(n_6462),
.A2(n_196),
.B(n_197),
.Y(n_6880)
);

NAND2x1p5_ASAP7_75t_L g6881 ( 
.A(n_6598),
.B(n_6648),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6464),
.Y(n_6882)
);

NAND2xp5_ASAP7_75t_L g6883 ( 
.A(n_6521),
.B(n_197),
.Y(n_6883)
);

NAND2x1p5_ASAP7_75t_L g6884 ( 
.A(n_6648),
.B(n_2745),
.Y(n_6884)
);

BUFx6f_ASAP7_75t_L g6885 ( 
.A(n_6437),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6500),
.B(n_199),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_L g6887 ( 
.A(n_6655),
.B(n_200),
.Y(n_6887)
);

OAI21x1_ASAP7_75t_L g6888 ( 
.A1(n_6542),
.A2(n_200),
.B(n_201),
.Y(n_6888)
);

HB1xp67_ASAP7_75t_L g6889 ( 
.A(n_6485),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6498),
.Y(n_6890)
);

INVx4_ASAP7_75t_L g6891 ( 
.A(n_6482),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6519),
.Y(n_6892)
);

AOI21x1_ASAP7_75t_L g6893 ( 
.A1(n_6655),
.A2(n_201),
.B(n_205),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6531),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_6547),
.Y(n_6895)
);

OA21x2_ASAP7_75t_L g6896 ( 
.A1(n_6684),
.A2(n_205),
.B(n_206),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_L g6897 ( 
.A(n_6686),
.B(n_206),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6575),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6654),
.Y(n_6899)
);

AND2x4_ASAP7_75t_L g6900 ( 
.A(n_6664),
.B(n_207),
.Y(n_6900)
);

OA21x2_ASAP7_75t_L g6901 ( 
.A1(n_6691),
.A2(n_208),
.B(n_209),
.Y(n_6901)
);

AND2x4_ASAP7_75t_L g6902 ( 
.A(n_6664),
.B(n_6500),
.Y(n_6902)
);

AO31x2_ASAP7_75t_L g6903 ( 
.A1(n_6675),
.A2(n_212),
.A3(n_210),
.B(n_211),
.Y(n_6903)
);

OA21x2_ASAP7_75t_L g6904 ( 
.A1(n_6626),
.A2(n_211),
.B(n_214),
.Y(n_6904)
);

AOI21xp5_ASAP7_75t_L g6905 ( 
.A1(n_6497),
.A2(n_214),
.B(n_216),
.Y(n_6905)
);

AO31x2_ASAP7_75t_L g6906 ( 
.A1(n_6637),
.A2(n_219),
.A3(n_217),
.B(n_218),
.Y(n_6906)
);

AOI21xp33_ASAP7_75t_SL g6907 ( 
.A1(n_6468),
.A2(n_219),
.B(n_220),
.Y(n_6907)
);

NAND2xp5_ASAP7_75t_L g6908 ( 
.A(n_6672),
.B(n_221),
.Y(n_6908)
);

AOI22xp33_ASAP7_75t_L g6909 ( 
.A1(n_6551),
.A2(n_2413),
.B1(n_2408),
.B2(n_2343),
.Y(n_6909)
);

OA21x2_ASAP7_75t_L g6910 ( 
.A1(n_6678),
.A2(n_221),
.B(n_222),
.Y(n_6910)
);

INVx2_ASAP7_75t_L g6911 ( 
.A(n_6672),
.Y(n_6911)
);

INVx8_ASAP7_75t_L g6912 ( 
.A(n_6599),
.Y(n_6912)
);

AND2x4_ASAP7_75t_L g6913 ( 
.A(n_6518),
.B(n_222),
.Y(n_6913)
);

OAI21x1_ASAP7_75t_L g6914 ( 
.A1(n_6487),
.A2(n_223),
.B(n_224),
.Y(n_6914)
);

NAND2xp5_ASAP7_75t_L g6915 ( 
.A(n_6672),
.B(n_223),
.Y(n_6915)
);

AND2x2_ASAP7_75t_L g6916 ( 
.A(n_6518),
.B(n_6478),
.Y(n_6916)
);

OAI21x1_ASAP7_75t_L g6917 ( 
.A1(n_6467),
.A2(n_225),
.B(n_227),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6575),
.Y(n_6918)
);

INVx2_ASAP7_75t_L g6919 ( 
.A(n_6478),
.Y(n_6919)
);

BUFx2_ASAP7_75t_L g6920 ( 
.A(n_6440),
.Y(n_6920)
);

INVx1_ASAP7_75t_L g6921 ( 
.A(n_6575),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6613),
.Y(n_6922)
);

OAI21xp5_ASAP7_75t_L g6923 ( 
.A1(n_6659),
.A2(n_227),
.B(n_228),
.Y(n_6923)
);

AO21x2_ASAP7_75t_L g6924 ( 
.A1(n_6603),
.A2(n_229),
.B(n_230),
.Y(n_6924)
);

OR2x6_ASAP7_75t_L g6925 ( 
.A(n_6599),
.B(n_6478),
.Y(n_6925)
);

INVx2_ASAP7_75t_L g6926 ( 
.A(n_6550),
.Y(n_6926)
);

AOI21xp33_ASAP7_75t_SL g6927 ( 
.A1(n_6683),
.A2(n_230),
.B(n_231),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6613),
.Y(n_6928)
);

BUFx3_ASAP7_75t_L g6929 ( 
.A(n_6558),
.Y(n_6929)
);

NAND2x1_ASAP7_75t_L g6930 ( 
.A(n_6440),
.B(n_3948),
.Y(n_6930)
);

AOI21xp5_ASAP7_75t_L g6931 ( 
.A1(n_6557),
.A2(n_231),
.B(n_232),
.Y(n_6931)
);

AO21x2_ASAP7_75t_L g6932 ( 
.A1(n_6666),
.A2(n_232),
.B(n_235),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6613),
.Y(n_6933)
);

NAND2xp5_ASAP7_75t_L g6934 ( 
.A(n_6548),
.B(n_6525),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_6550),
.Y(n_6935)
);

INVx2_ASAP7_75t_L g6936 ( 
.A(n_6550),
.Y(n_6936)
);

AOI21xp5_ASAP7_75t_L g6937 ( 
.A1(n_6541),
.A2(n_236),
.B(n_237),
.Y(n_6937)
);

OA21x2_ASAP7_75t_L g6938 ( 
.A1(n_6534),
.A2(n_237),
.B(n_238),
.Y(n_6938)
);

AO21x2_ASAP7_75t_L g6939 ( 
.A1(n_6666),
.A2(n_238),
.B(n_239),
.Y(n_6939)
);

NAND2xp5_ASAP7_75t_L g6940 ( 
.A(n_6548),
.B(n_239),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6615),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_6694),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6699),
.Y(n_6943)
);

INVx2_ASAP7_75t_L g6944 ( 
.A(n_6779),
.Y(n_6944)
);

INVx2_ASAP7_75t_L g6945 ( 
.A(n_6779),
.Y(n_6945)
);

INVx3_ASAP7_75t_L g6946 ( 
.A(n_6696),
.Y(n_6946)
);

NAND2xp5_ASAP7_75t_L g6947 ( 
.A(n_6922),
.B(n_6615),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_L g6948 ( 
.A(n_6928),
.B(n_6615),
.Y(n_6948)
);

OAI21x1_ASAP7_75t_L g6949 ( 
.A1(n_6733),
.A2(n_6687),
.B(n_6661),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6703),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6706),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_6779),
.Y(n_6952)
);

OA21x2_ASAP7_75t_L g6953 ( 
.A1(n_6747),
.A2(n_6571),
.B(n_6567),
.Y(n_6953)
);

AO31x2_ASAP7_75t_L g6954 ( 
.A1(n_6747),
.A2(n_6578),
.A3(n_6621),
.B(n_6610),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6720),
.Y(n_6955)
);

BUFx3_ASAP7_75t_L g6956 ( 
.A(n_6738),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6721),
.Y(n_6957)
);

HB1xp67_ASAP7_75t_L g6958 ( 
.A(n_6855),
.Y(n_6958)
);

AOI22xp33_ASAP7_75t_SL g6959 ( 
.A1(n_6713),
.A2(n_6569),
.B1(n_6649),
.B2(n_6563),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6726),
.Y(n_6960)
);

NAND2xp5_ASAP7_75t_L g6961 ( 
.A(n_6933),
.B(n_6941),
.Y(n_6961)
);

OR2x2_ASAP7_75t_L g6962 ( 
.A(n_6843),
.B(n_6525),
.Y(n_6962)
);

INVx2_ASAP7_75t_L g6963 ( 
.A(n_6823),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_6823),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6727),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6730),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6739),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6740),
.Y(n_6968)
);

BUFx3_ASAP7_75t_L g6969 ( 
.A(n_6752),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6776),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6783),
.Y(n_6971)
);

OAI21x1_ASAP7_75t_L g6972 ( 
.A1(n_6733),
.A2(n_6708),
.B(n_6704),
.Y(n_6972)
);

OAI21x1_ASAP7_75t_L g6973 ( 
.A1(n_6723),
.A2(n_6734),
.B(n_6702),
.Y(n_6973)
);

NAND2xp5_ASAP7_75t_L g6974 ( 
.A(n_6846),
.B(n_6621),
.Y(n_6974)
);

INVx2_ASAP7_75t_L g6975 ( 
.A(n_6753),
.Y(n_6975)
);

OR2x2_ASAP7_75t_L g6976 ( 
.A(n_6711),
.B(n_6525),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6818),
.Y(n_6977)
);

BUFx3_ASAP7_75t_L g6978 ( 
.A(n_6929),
.Y(n_6978)
);

AND2x4_ASAP7_75t_L g6979 ( 
.A(n_6724),
.B(n_6549),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6822),
.Y(n_6980)
);

BUFx2_ASAP7_75t_L g6981 ( 
.A(n_6925),
.Y(n_6981)
);

INVx2_ASAP7_75t_L g6982 ( 
.A(n_6823),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_6832),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6809),
.Y(n_6984)
);

OAI21x1_ASAP7_75t_L g6985 ( 
.A1(n_6824),
.A2(n_6589),
.B(n_6524),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6791),
.Y(n_6986)
);

OAI21x1_ASAP7_75t_L g6987 ( 
.A1(n_6724),
.A2(n_6524),
.B(n_6562),
.Y(n_6987)
);

OR2x2_ASAP7_75t_L g6988 ( 
.A(n_6874),
.B(n_6548),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6837),
.Y(n_6989)
);

HB1xp67_ASAP7_75t_L g6990 ( 
.A(n_6761),
.Y(n_6990)
);

AOI21xp5_ASAP7_75t_L g6991 ( 
.A1(n_6710),
.A2(n_6774),
.B(n_6714),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6896),
.Y(n_6992)
);

OAI22xp5_ASAP7_75t_L g6993 ( 
.A1(n_6732),
.A2(n_6473),
.B1(n_6459),
.B2(n_6625),
.Y(n_6993)
);

BUFx3_ASAP7_75t_L g6994 ( 
.A(n_6819),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6896),
.Y(n_6995)
);

INVx2_ASAP7_75t_L g6996 ( 
.A(n_6705),
.Y(n_6996)
);

INVx2_ASAP7_75t_L g6997 ( 
.A(n_6705),
.Y(n_6997)
);

BUFx2_ASAP7_75t_L g6998 ( 
.A(n_6925),
.Y(n_6998)
);

INVx2_ASAP7_75t_L g6999 ( 
.A(n_6809),
.Y(n_6999)
);

INVx3_ASAP7_75t_L g7000 ( 
.A(n_6912),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6901),
.Y(n_7001)
);

OAI22xp5_ASAP7_75t_L g7002 ( 
.A1(n_6741),
.A2(n_6459),
.B1(n_6539),
.B2(n_6665),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_L g7003 ( 
.A(n_6850),
.B(n_6621),
.Y(n_7003)
);

INVx1_ASAP7_75t_SL g7004 ( 
.A(n_6718),
.Y(n_7004)
);

INVx2_ASAP7_75t_L g7005 ( 
.A(n_6885),
.Y(n_7005)
);

OR2x2_ASAP7_75t_L g7006 ( 
.A(n_6839),
.B(n_6728),
.Y(n_7006)
);

AO21x2_ASAP7_75t_L g7007 ( 
.A1(n_6851),
.A2(n_6638),
.B(n_6631),
.Y(n_7007)
);

OAI21x1_ASAP7_75t_L g7008 ( 
.A1(n_6862),
.A2(n_6640),
.B(n_6587),
.Y(n_7008)
);

OA21x2_ASAP7_75t_L g7009 ( 
.A1(n_6698),
.A2(n_6669),
.B(n_6663),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6901),
.Y(n_7010)
);

NAND2x1p5_ASAP7_75t_L g7011 ( 
.A(n_6770),
.B(n_6938),
.Y(n_7011)
);

INVx3_ASAP7_75t_L g7012 ( 
.A(n_6912),
.Y(n_7012)
);

BUFx6f_ASAP7_75t_L g7013 ( 
.A(n_6735),
.Y(n_7013)
);

INVx2_ASAP7_75t_L g7014 ( 
.A(n_6885),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_6881),
.Y(n_7015)
);

OA21x2_ASAP7_75t_L g7016 ( 
.A1(n_6876),
.A2(n_6676),
.B(n_6624),
.Y(n_7016)
);

INVx2_ASAP7_75t_L g7017 ( 
.A(n_6798),
.Y(n_7017)
);

AND2x2_ASAP7_75t_L g7018 ( 
.A(n_6831),
.B(n_6535),
.Y(n_7018)
);

OAI22xp5_ASAP7_75t_L g7019 ( 
.A1(n_6701),
.A2(n_6760),
.B1(n_6709),
.B2(n_6847),
.Y(n_7019)
);

INVx2_ASAP7_75t_L g7020 ( 
.A(n_6751),
.Y(n_7020)
);

INVx2_ASAP7_75t_L g7021 ( 
.A(n_6830),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6746),
.Y(n_7022)
);

HB1xp67_ASAP7_75t_L g7023 ( 
.A(n_6938),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6800),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6812),
.Y(n_7025)
);

OAI21xp33_ASAP7_75t_SL g7026 ( 
.A1(n_6790),
.A2(n_6623),
.B(n_6650),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6860),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6840),
.Y(n_7028)
);

INVx2_ASAP7_75t_L g7029 ( 
.A(n_6772),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6898),
.Y(n_7030)
);

INVx2_ASAP7_75t_L g7031 ( 
.A(n_6808),
.Y(n_7031)
);

HB1xp67_ASAP7_75t_SL g7032 ( 
.A(n_6878),
.Y(n_7032)
);

INVx1_ASAP7_75t_L g7033 ( 
.A(n_6918),
.Y(n_7033)
);

INVx2_ASAP7_75t_L g7034 ( 
.A(n_6920),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6921),
.Y(n_7035)
);

AOI21x1_ASAP7_75t_L g7036 ( 
.A1(n_6883),
.A2(n_6539),
.B(n_6535),
.Y(n_7036)
);

INVx2_ASAP7_75t_L g7037 ( 
.A(n_6913),
.Y(n_7037)
);

AND2x4_ASAP7_75t_L g7038 ( 
.A(n_6913),
.B(n_6549),
.Y(n_7038)
);

INVx1_ASAP7_75t_L g7039 ( 
.A(n_6882),
.Y(n_7039)
);

BUFx2_ASAP7_75t_L g7040 ( 
.A(n_6773),
.Y(n_7040)
);

AOI22xp5_ASAP7_75t_L g7041 ( 
.A1(n_6905),
.A2(n_6560),
.B1(n_6559),
.B2(n_6629),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6920),
.Y(n_7042)
);

CKINVDCx20_ASAP7_75t_R g7043 ( 
.A(n_6717),
.Y(n_7043)
);

AOI22xp33_ASAP7_75t_SL g7044 ( 
.A1(n_6764),
.A2(n_6641),
.B1(n_6486),
.B2(n_6517),
.Y(n_7044)
);

INVx2_ASAP7_75t_L g7045 ( 
.A(n_6775),
.Y(n_7045)
);

INVx2_ASAP7_75t_L g7046 ( 
.A(n_6775),
.Y(n_7046)
);

INVx2_ASAP7_75t_L g7047 ( 
.A(n_6722),
.Y(n_7047)
);

AND2x2_ASAP7_75t_L g7048 ( 
.A(n_6916),
.B(n_6486),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6890),
.Y(n_7049)
);

AND2x2_ASAP7_75t_L g7050 ( 
.A(n_6841),
.B(n_6815),
.Y(n_7050)
);

AND2x2_ASAP7_75t_L g7051 ( 
.A(n_6841),
.B(n_6486),
.Y(n_7051)
);

OA21x2_ASAP7_75t_L g7052 ( 
.A1(n_6801),
.A2(n_6517),
.B(n_240),
.Y(n_7052)
);

OR2x2_ASAP7_75t_L g7053 ( 
.A(n_6934),
.B(n_242),
.Y(n_7053)
);

INVx1_ASAP7_75t_L g7054 ( 
.A(n_6892),
.Y(n_7054)
);

INVx2_ASAP7_75t_L g7055 ( 
.A(n_6763),
.Y(n_7055)
);

INVx2_ASAP7_75t_SL g7056 ( 
.A(n_6735),
.Y(n_7056)
);

INVxp33_ASAP7_75t_L g7057 ( 
.A(n_6697),
.Y(n_7057)
);

INVx1_ASAP7_75t_L g7058 ( 
.A(n_6894),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_6895),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6889),
.Y(n_7060)
);

NAND2xp5_ASAP7_75t_L g7061 ( 
.A(n_6712),
.B(n_242),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_6940),
.Y(n_7062)
);

INVx2_ASAP7_75t_L g7063 ( 
.A(n_6763),
.Y(n_7063)
);

BUFx3_ASAP7_75t_L g7064 ( 
.A(n_6856),
.Y(n_7064)
);

OAI21x1_ASAP7_75t_L g7065 ( 
.A1(n_6748),
.A2(n_245),
.B(n_247),
.Y(n_7065)
);

AOI21xp5_ASAP7_75t_L g7066 ( 
.A1(n_6780),
.A2(n_245),
.B(n_248),
.Y(n_7066)
);

HB1xp67_ASAP7_75t_L g7067 ( 
.A(n_6910),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6919),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6926),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6935),
.Y(n_7070)
);

INVx2_ASAP7_75t_L g7071 ( 
.A(n_6763),
.Y(n_7071)
);

CKINVDCx6p67_ASAP7_75t_R g7072 ( 
.A(n_6716),
.Y(n_7072)
);

AND2x2_ASAP7_75t_L g7073 ( 
.A(n_6815),
.B(n_6827),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6936),
.Y(n_7074)
);

AND2x2_ASAP7_75t_L g7075 ( 
.A(n_6810),
.B(n_249),
.Y(n_7075)
);

INVx1_ASAP7_75t_L g7076 ( 
.A(n_6886),
.Y(n_7076)
);

AO21x2_ASAP7_75t_L g7077 ( 
.A1(n_6868),
.A2(n_250),
.B(n_251),
.Y(n_7077)
);

INVx2_ASAP7_75t_L g7078 ( 
.A(n_6825),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6749),
.Y(n_7079)
);

INVx2_ASAP7_75t_L g7080 ( 
.A(n_6754),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_6758),
.Y(n_7081)
);

INVx2_ASAP7_75t_L g7082 ( 
.A(n_6768),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_6829),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6778),
.Y(n_7084)
);

HB1xp67_ASAP7_75t_L g7085 ( 
.A(n_6910),
.Y(n_7085)
);

INVx3_ASAP7_75t_L g7086 ( 
.A(n_6891),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6785),
.Y(n_7087)
);

INVx2_ASAP7_75t_L g7088 ( 
.A(n_6842),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_6796),
.B(n_250),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6820),
.Y(n_7090)
);

INVx2_ASAP7_75t_L g7091 ( 
.A(n_6859),
.Y(n_7091)
);

AO21x2_ASAP7_75t_L g7092 ( 
.A1(n_6700),
.A2(n_252),
.B(n_253),
.Y(n_7092)
);

AND2x2_ASAP7_75t_L g7093 ( 
.A(n_6810),
.B(n_6873),
.Y(n_7093)
);

INVx2_ASAP7_75t_L g7094 ( 
.A(n_6899),
.Y(n_7094)
);

INVx5_ASAP7_75t_SL g7095 ( 
.A(n_6924),
.Y(n_7095)
);

OAI21x1_ASAP7_75t_L g7096 ( 
.A1(n_6870),
.A2(n_252),
.B(n_253),
.Y(n_7096)
);

NAND2x1p5_ASAP7_75t_L g7097 ( 
.A(n_6828),
.B(n_6743),
.Y(n_7097)
);

INVxp67_ASAP7_75t_L g7098 ( 
.A(n_6742),
.Y(n_7098)
);

AOI22xp33_ASAP7_75t_L g7099 ( 
.A1(n_6744),
.A2(n_2247),
.B1(n_2278),
.B2(n_2166),
.Y(n_7099)
);

OR2x2_ASAP7_75t_L g7100 ( 
.A(n_6826),
.B(n_254),
.Y(n_7100)
);

OA21x2_ASAP7_75t_L g7101 ( 
.A1(n_6750),
.A2(n_254),
.B(n_255),
.Y(n_7101)
);

CKINVDCx5p33_ASAP7_75t_R g7102 ( 
.A(n_6856),
.Y(n_7102)
);

INVx2_ASAP7_75t_L g7103 ( 
.A(n_6911),
.Y(n_7103)
);

INVx2_ASAP7_75t_L g7104 ( 
.A(n_6854),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6853),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6863),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_6867),
.Y(n_7107)
);

INVx1_ASAP7_75t_SL g7108 ( 
.A(n_6804),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6849),
.Y(n_7109)
);

INVx2_ASAP7_75t_L g7110 ( 
.A(n_6719),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_6745),
.B(n_255),
.Y(n_7111)
);

AND2x2_ASAP7_75t_L g7112 ( 
.A(n_6731),
.B(n_257),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_6932),
.Y(n_7113)
);

AO21x2_ASAP7_75t_L g7114 ( 
.A1(n_6797),
.A2(n_258),
.B(n_260),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_6939),
.Y(n_7115)
);

INVx2_ASAP7_75t_SL g7116 ( 
.A(n_6872),
.Y(n_7116)
);

INVx2_ASAP7_75t_SL g7117 ( 
.A(n_6731),
.Y(n_7117)
);

OA21x2_ASAP7_75t_L g7118 ( 
.A1(n_6765),
.A2(n_261),
.B(n_262),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6805),
.Y(n_7119)
);

OAI21x1_ASAP7_75t_L g7120 ( 
.A1(n_6729),
.A2(n_261),
.B(n_265),
.Y(n_7120)
);

BUFx2_ASAP7_75t_L g7121 ( 
.A(n_6833),
.Y(n_7121)
);

INVx1_ASAP7_75t_L g7122 ( 
.A(n_6904),
.Y(n_7122)
);

INVx1_ASAP7_75t_L g7123 ( 
.A(n_6904),
.Y(n_7123)
);

INVx2_ASAP7_75t_L g7124 ( 
.A(n_6884),
.Y(n_7124)
);

INVx2_ASAP7_75t_L g7125 ( 
.A(n_6902),
.Y(n_7125)
);

AND2x2_ASAP7_75t_L g7126 ( 
.A(n_6803),
.B(n_265),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6917),
.Y(n_7127)
);

OR2x2_ASAP7_75t_L g7128 ( 
.A(n_6869),
.B(n_266),
.Y(n_7128)
);

AND2x2_ASAP7_75t_L g7129 ( 
.A(n_6756),
.B(n_266),
.Y(n_7129)
);

BUFx3_ASAP7_75t_L g7130 ( 
.A(n_6864),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_6893),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6893),
.Y(n_7132)
);

BUFx3_ASAP7_75t_L g7133 ( 
.A(n_6857),
.Y(n_7133)
);

AOI21xp33_ASAP7_75t_SL g7134 ( 
.A1(n_6880),
.A2(n_6762),
.B(n_6781),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6838),
.Y(n_7135)
);

BUFx2_ASAP7_75t_SL g7136 ( 
.A(n_6900),
.Y(n_7136)
);

CKINVDCx20_ASAP7_75t_R g7137 ( 
.A(n_6897),
.Y(n_7137)
);

HB1xp67_ASAP7_75t_L g7138 ( 
.A(n_6695),
.Y(n_7138)
);

INVx2_ASAP7_75t_L g7139 ( 
.A(n_6902),
.Y(n_7139)
);

INVx2_ASAP7_75t_SL g7140 ( 
.A(n_6766),
.Y(n_7140)
);

OAI22xp5_ASAP7_75t_L g7141 ( 
.A1(n_6788),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_7141)
);

INVx2_ASAP7_75t_SL g7142 ( 
.A(n_6766),
.Y(n_7142)
);

INVx2_ASAP7_75t_L g7143 ( 
.A(n_6813),
.Y(n_7143)
);

AND2x2_ASAP7_75t_L g7144 ( 
.A(n_6766),
.B(n_6795),
.Y(n_7144)
);

NAND2xp33_ASAP7_75t_L g7145 ( 
.A(n_6865),
.B(n_3948),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6877),
.Y(n_7146)
);

AND2x2_ASAP7_75t_L g7147 ( 
.A(n_6759),
.B(n_267),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6914),
.Y(n_7148)
);

INVx3_ASAP7_75t_L g7149 ( 
.A(n_6719),
.Y(n_7149)
);

INVxp67_ASAP7_75t_L g7150 ( 
.A(n_6857),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6836),
.Y(n_7151)
);

INVx1_ASAP7_75t_L g7152 ( 
.A(n_6737),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6737),
.Y(n_7153)
);

AO21x2_ASAP7_75t_L g7154 ( 
.A1(n_6725),
.A2(n_6828),
.B(n_6845),
.Y(n_7154)
);

AND2x4_ASAP7_75t_L g7155 ( 
.A(n_6737),
.B(n_269),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6888),
.Y(n_7156)
);

INVx2_ASAP7_75t_L g7157 ( 
.A(n_6784),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_6908),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_6900),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_6806),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6915),
.Y(n_7161)
);

BUFx3_ASAP7_75t_L g7162 ( 
.A(n_6866),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_6792),
.Y(n_7163)
);

CKINVDCx20_ASAP7_75t_R g7164 ( 
.A(n_6879),
.Y(n_7164)
);

HB1xp67_ASAP7_75t_L g7165 ( 
.A(n_6736),
.Y(n_7165)
);

INVx3_ASAP7_75t_L g7166 ( 
.A(n_6834),
.Y(n_7166)
);

AND2x2_ASAP7_75t_L g7167 ( 
.A(n_6793),
.B(n_270),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6767),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6799),
.Y(n_7169)
);

AND2x2_ASAP7_75t_L g7170 ( 
.A(n_6769),
.B(n_271),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_6725),
.Y(n_7171)
);

HB1xp67_ASAP7_75t_L g7172 ( 
.A(n_6736),
.Y(n_7172)
);

AND2x2_ASAP7_75t_L g7173 ( 
.A(n_7050),
.B(n_6861),
.Y(n_7173)
);

AOI22xp33_ASAP7_75t_L g7174 ( 
.A1(n_7019),
.A2(n_6937),
.B1(n_6871),
.B2(n_6816),
.Y(n_7174)
);

AOI22xp33_ASAP7_75t_SL g7175 ( 
.A1(n_7019),
.A2(n_6835),
.B1(n_6923),
.B2(n_6852),
.Y(n_7175)
);

OAI22xp5_ASAP7_75t_L g7176 ( 
.A1(n_6991),
.A2(n_6909),
.B1(n_6821),
.B2(n_6848),
.Y(n_7176)
);

A2O1A1Ixp33_ASAP7_75t_L g7177 ( 
.A1(n_6991),
.A2(n_6927),
.B(n_6858),
.C(n_6907),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6958),
.Y(n_7178)
);

OAI221xp5_ASAP7_75t_L g7179 ( 
.A1(n_7026),
.A2(n_6887),
.B1(n_6817),
.B2(n_6814),
.C(n_6786),
.Y(n_7179)
);

AOI22xp33_ASAP7_75t_L g7180 ( 
.A1(n_7057),
.A2(n_6787),
.B1(n_6693),
.B2(n_6802),
.Y(n_7180)
);

OAI22xp5_ASAP7_75t_L g7181 ( 
.A1(n_7095),
.A2(n_6782),
.B1(n_6930),
.B2(n_6693),
.Y(n_7181)
);

OAI22xp33_ASAP7_75t_L g7182 ( 
.A1(n_7004),
.A2(n_6782),
.B1(n_6930),
.B2(n_6834),
.Y(n_7182)
);

OAI221xp5_ASAP7_75t_L g7183 ( 
.A1(n_7026),
.A2(n_6811),
.B1(n_6931),
.B2(n_6875),
.C(n_6757),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6958),
.Y(n_7184)
);

OAI21xp33_ASAP7_75t_L g7185 ( 
.A1(n_7057),
.A2(n_6777),
.B(n_6755),
.Y(n_7185)
);

OAI22xp5_ASAP7_75t_L g7186 ( 
.A1(n_7095),
.A2(n_6707),
.B1(n_6757),
.B2(n_6844),
.Y(n_7186)
);

AND2x2_ASAP7_75t_L g7187 ( 
.A(n_7040),
.B(n_6736),
.Y(n_7187)
);

OR2x2_ASAP7_75t_L g7188 ( 
.A(n_7108),
.B(n_6866),
.Y(n_7188)
);

AOI22xp33_ASAP7_75t_SL g7189 ( 
.A1(n_7095),
.A2(n_6707),
.B1(n_6806),
.B2(n_6771),
.Y(n_7189)
);

AOI22xp33_ASAP7_75t_L g7190 ( 
.A1(n_6993),
.A2(n_6715),
.B1(n_6794),
.B2(n_6807),
.Y(n_7190)
);

AOI22xp33_ASAP7_75t_L g7191 ( 
.A1(n_6993),
.A2(n_6715),
.B1(n_6794),
.B2(n_6807),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_7030),
.Y(n_7192)
);

INVx2_ASAP7_75t_L g7193 ( 
.A(n_6978),
.Y(n_7193)
);

AND2x4_ASAP7_75t_L g7194 ( 
.A(n_7064),
.B(n_6789),
.Y(n_7194)
);

AOI222xp33_ASAP7_75t_L g7195 ( 
.A1(n_7062),
.A2(n_6903),
.B1(n_6906),
.B2(n_273),
.C1(n_275),
.C2(n_271),
.Y(n_7195)
);

OAI21xp33_ASAP7_75t_SL g7196 ( 
.A1(n_7004),
.A2(n_6903),
.B(n_6906),
.Y(n_7196)
);

AND2x2_ASAP7_75t_L g7197 ( 
.A(n_7073),
.B(n_6844),
.Y(n_7197)
);

OAI22xp5_ASAP7_75t_L g7198 ( 
.A1(n_6959),
.A2(n_275),
.B1(n_272),
.B2(n_274),
.Y(n_7198)
);

AND2x2_ASAP7_75t_L g7199 ( 
.A(n_7086),
.B(n_272),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_7033),
.Y(n_7200)
);

AOI22xp33_ASAP7_75t_L g7201 ( 
.A1(n_7044),
.A2(n_2413),
.B1(n_2343),
.B2(n_2344),
.Y(n_7201)
);

AOI221xp5_ASAP7_75t_L g7202 ( 
.A1(n_7141),
.A2(n_277),
.B1(n_274),
.B2(n_276),
.C(n_278),
.Y(n_7202)
);

AND2x2_ASAP7_75t_L g7203 ( 
.A(n_7086),
.B(n_7072),
.Y(n_7203)
);

AOI21xp5_ASAP7_75t_L g7204 ( 
.A1(n_7066),
.A2(n_277),
.B(n_278),
.Y(n_7204)
);

INVx1_ASAP7_75t_L g7205 ( 
.A(n_7035),
.Y(n_7205)
);

OAI22xp5_ASAP7_75t_L g7206 ( 
.A1(n_6959),
.A2(n_282),
.B1(n_279),
.B2(n_280),
.Y(n_7206)
);

AOI21xp5_ASAP7_75t_L g7207 ( 
.A1(n_7066),
.A2(n_279),
.B(n_282),
.Y(n_7207)
);

AOI21xp5_ASAP7_75t_L g7208 ( 
.A1(n_7141),
.A2(n_284),
.B(n_285),
.Y(n_7208)
);

INVx2_ASAP7_75t_L g7209 ( 
.A(n_6978),
.Y(n_7209)
);

A2O1A1Ixp33_ASAP7_75t_L g7210 ( 
.A1(n_7134),
.A2(n_7162),
.B(n_7133),
.C(n_7150),
.Y(n_7210)
);

OR2x2_ASAP7_75t_L g7211 ( 
.A(n_7108),
.B(n_285),
.Y(n_7211)
);

AOI221xp5_ASAP7_75t_L g7212 ( 
.A1(n_7002),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.C(n_291),
.Y(n_7212)
);

HB1xp67_ASAP7_75t_L g7213 ( 
.A(n_6990),
.Y(n_7213)
);

OAI22xp5_ASAP7_75t_L g7214 ( 
.A1(n_7044),
.A2(n_296),
.B1(n_292),
.B2(n_293),
.Y(n_7214)
);

NAND3xp33_ASAP7_75t_L g7215 ( 
.A(n_7023),
.B(n_293),
.C(n_299),
.Y(n_7215)
);

AND2x4_ASAP7_75t_L g7216 ( 
.A(n_7064),
.B(n_299),
.Y(n_7216)
);

AND2x2_ASAP7_75t_L g7217 ( 
.A(n_7093),
.B(n_300),
.Y(n_7217)
);

OAI22xp33_ASAP7_75t_L g7218 ( 
.A1(n_7041),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_7218)
);

INVx1_ASAP7_75t_L g7219 ( 
.A(n_6961),
.Y(n_7219)
);

AOI22xp33_ASAP7_75t_SL g7220 ( 
.A1(n_7162),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_7220)
);

AOI22xp33_ASAP7_75t_L g7221 ( 
.A1(n_7009),
.A2(n_2343),
.B1(n_2344),
.B2(n_2332),
.Y(n_7221)
);

BUFx4f_ASAP7_75t_SL g7222 ( 
.A(n_6969),
.Y(n_7222)
);

OAI221xp5_ASAP7_75t_L g7223 ( 
.A1(n_7002),
.A2(n_307),
.B1(n_303),
.B2(n_306),
.C(n_309),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_6981),
.B(n_306),
.Y(n_7224)
);

NAND2xp5_ASAP7_75t_L g7225 ( 
.A(n_7150),
.B(n_309),
.Y(n_7225)
);

NOR2x1_ASAP7_75t_L g7226 ( 
.A(n_7092),
.B(n_310),
.Y(n_7226)
);

OR2x6_ASAP7_75t_L g7227 ( 
.A(n_7130),
.B(n_310),
.Y(n_7227)
);

AOI22xp33_ASAP7_75t_L g7228 ( 
.A1(n_7009),
.A2(n_2343),
.B1(n_2344),
.B2(n_2332),
.Y(n_7228)
);

AND2x2_ASAP7_75t_L g7229 ( 
.A(n_6998),
.B(n_311),
.Y(n_7229)
);

AOI22xp33_ASAP7_75t_L g7230 ( 
.A1(n_7130),
.A2(n_2343),
.B1(n_2344),
.B2(n_2332),
.Y(n_7230)
);

OAI22xp5_ASAP7_75t_L g7231 ( 
.A1(n_7041),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_7231)
);

AOI22xp5_ASAP7_75t_L g7232 ( 
.A1(n_7092),
.A2(n_4070),
.B1(n_4049),
.B2(n_4003),
.Y(n_7232)
);

AOI22xp33_ASAP7_75t_L g7233 ( 
.A1(n_7121),
.A2(n_2344),
.B1(n_2345),
.B2(n_2332),
.Y(n_7233)
);

INVx2_ASAP7_75t_L g7234 ( 
.A(n_7013),
.Y(n_7234)
);

OAI21x1_ASAP7_75t_L g7235 ( 
.A1(n_6972),
.A2(n_313),
.B(n_314),
.Y(n_7235)
);

AOI21xp5_ASAP7_75t_L g7236 ( 
.A1(n_7155),
.A2(n_314),
.B(n_315),
.Y(n_7236)
);

BUFx3_ASAP7_75t_L g7237 ( 
.A(n_6969),
.Y(n_7237)
);

AO21x2_ASAP7_75t_L g7238 ( 
.A1(n_7138),
.A2(n_316),
.B(n_317),
.Y(n_7238)
);

AOI221xp5_ASAP7_75t_L g7239 ( 
.A1(n_6990),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.C(n_319),
.Y(n_7239)
);

OAI21xp33_ASAP7_75t_L g7240 ( 
.A1(n_6989),
.A2(n_318),
.B(n_319),
.Y(n_7240)
);

AOI221xp5_ASAP7_75t_L g7241 ( 
.A1(n_7023),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C(n_326),
.Y(n_7241)
);

INVx3_ASAP7_75t_L g7242 ( 
.A(n_7013),
.Y(n_7242)
);

INVx2_ASAP7_75t_L g7243 ( 
.A(n_7013),
.Y(n_7243)
);

NAND3xp33_ASAP7_75t_SL g7244 ( 
.A(n_7144),
.B(n_326),
.C(n_327),
.Y(n_7244)
);

INVx4_ASAP7_75t_L g7245 ( 
.A(n_7102),
.Y(n_7245)
);

OAI22xp5_ASAP7_75t_L g7246 ( 
.A1(n_7052),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_7246)
);

AOI22xp33_ASAP7_75t_L g7247 ( 
.A1(n_7168),
.A2(n_2345),
.B1(n_2357),
.B2(n_2332),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_6961),
.Y(n_7248)
);

AOI22xp33_ASAP7_75t_L g7249 ( 
.A1(n_7015),
.A2(n_2357),
.B1(n_2366),
.B2(n_2345),
.Y(n_7249)
);

AOI21xp5_ASAP7_75t_L g7250 ( 
.A1(n_7155),
.A2(n_7115),
.B(n_7113),
.Y(n_7250)
);

AOI22xp33_ASAP7_75t_L g7251 ( 
.A1(n_7169),
.A2(n_2357),
.B1(n_2366),
.B2(n_2345),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6942),
.Y(n_7252)
);

AND2x4_ASAP7_75t_L g7253 ( 
.A(n_7078),
.B(n_329),
.Y(n_7253)
);

OAI221xp5_ASAP7_75t_L g7254 ( 
.A1(n_7133),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_7254)
);

OAI22xp5_ASAP7_75t_L g7255 ( 
.A1(n_7052),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_7255)
);

NOR2xp33_ASAP7_75t_L g7256 ( 
.A(n_7032),
.B(n_334),
.Y(n_7256)
);

AOI22xp33_ASAP7_75t_L g7257 ( 
.A1(n_7151),
.A2(n_2357),
.B1(n_2366),
.B2(n_2345),
.Y(n_7257)
);

NOR2xp33_ASAP7_75t_L g7258 ( 
.A(n_7032),
.B(n_335),
.Y(n_7258)
);

AOI22xp33_ASAP7_75t_L g7259 ( 
.A1(n_7119),
.A2(n_2366),
.B1(n_2371),
.B2(n_2357),
.Y(n_7259)
);

INVx1_ASAP7_75t_L g7260 ( 
.A(n_6943),
.Y(n_7260)
);

OAI22xp5_ASAP7_75t_L g7261 ( 
.A1(n_7067),
.A2(n_339),
.B1(n_335),
.B2(n_338),
.Y(n_7261)
);

INVx2_ASAP7_75t_L g7262 ( 
.A(n_6994),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_6950),
.Y(n_7263)
);

INVx1_ASAP7_75t_L g7264 ( 
.A(n_6951),
.Y(n_7264)
);

AOI22xp33_ASAP7_75t_L g7265 ( 
.A1(n_7017),
.A2(n_2371),
.B1(n_2387),
.B2(n_2366),
.Y(n_7265)
);

INVx1_ASAP7_75t_SL g7266 ( 
.A(n_7043),
.Y(n_7266)
);

AOI22xp33_ASAP7_75t_SL g7267 ( 
.A1(n_7067),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_7267)
);

AND2x2_ASAP7_75t_L g7268 ( 
.A(n_7136),
.B(n_341),
.Y(n_7268)
);

OAI211xp5_ASAP7_75t_L g7269 ( 
.A1(n_7085),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_7269)
);

AOI22xp33_ASAP7_75t_L g7270 ( 
.A1(n_7047),
.A2(n_2387),
.B1(n_2393),
.B2(n_2371),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_6994),
.Y(n_7271)
);

OR2x2_ASAP7_75t_L g7272 ( 
.A(n_7109),
.B(n_343),
.Y(n_7272)
);

INVx2_ASAP7_75t_L g7273 ( 
.A(n_7056),
.Y(n_7273)
);

AOI221xp5_ASAP7_75t_L g7274 ( 
.A1(n_7098),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.C(n_347),
.Y(n_7274)
);

NAND2xp5_ASAP7_75t_L g7275 ( 
.A(n_7037),
.B(n_344),
.Y(n_7275)
);

OAI22xp5_ASAP7_75t_L g7276 ( 
.A1(n_7085),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_7276)
);

AOI221xp5_ASAP7_75t_L g7277 ( 
.A1(n_7098),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.C(n_352),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_6955),
.Y(n_7278)
);

AOI22xp33_ASAP7_75t_L g7279 ( 
.A1(n_7020),
.A2(n_2387),
.B1(n_2393),
.B2(n_2371),
.Y(n_7279)
);

OAI22xp33_ASAP7_75t_L g7280 ( 
.A1(n_6992),
.A2(n_353),
.B1(n_350),
.B2(n_352),
.Y(n_7280)
);

OAI22xp5_ASAP7_75t_L g7281 ( 
.A1(n_7011),
.A2(n_357),
.B1(n_354),
.B2(n_356),
.Y(n_7281)
);

OAI22xp33_ASAP7_75t_L g7282 ( 
.A1(n_6995),
.A2(n_359),
.B1(n_354),
.B2(n_356),
.Y(n_7282)
);

AOI22xp33_ASAP7_75t_L g7283 ( 
.A1(n_7135),
.A2(n_6946),
.B1(n_7018),
.B2(n_7114),
.Y(n_7283)
);

INVx2_ASAP7_75t_L g7284 ( 
.A(n_7000),
.Y(n_7284)
);

BUFx3_ASAP7_75t_L g7285 ( 
.A(n_7043),
.Y(n_7285)
);

AOI211xp5_ASAP7_75t_L g7286 ( 
.A1(n_7001),
.A2(n_365),
.B(n_361),
.C(n_362),
.Y(n_7286)
);

AOI222xp33_ASAP7_75t_L g7287 ( 
.A1(n_7129),
.A2(n_368),
.B1(n_370),
.B2(n_366),
.C1(n_367),
.C2(n_369),
.Y(n_7287)
);

HB1xp67_ASAP7_75t_L g7288 ( 
.A(n_7034),
.Y(n_7288)
);

OAI222xp33_ASAP7_75t_L g7289 ( 
.A1(n_7011),
.A2(n_371),
.B1(n_373),
.B2(n_369),
.C1(n_370),
.C2(n_372),
.Y(n_7289)
);

AOI22xp33_ASAP7_75t_SL g7290 ( 
.A1(n_7114),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_7290)
);

INVx1_ASAP7_75t_L g7291 ( 
.A(n_6957),
.Y(n_7291)
);

AOI33xp33_ASAP7_75t_L g7292 ( 
.A1(n_7010),
.A2(n_7122),
.A3(n_7123),
.B1(n_7152),
.B2(n_7153),
.B3(n_6975),
.Y(n_7292)
);

AOI22xp33_ASAP7_75t_L g7293 ( 
.A1(n_6946),
.A2(n_7154),
.B1(n_7117),
.B2(n_7139),
.Y(n_7293)
);

OAI221xp5_ASAP7_75t_L g7294 ( 
.A1(n_7171),
.A2(n_377),
.B1(n_374),
.B2(n_376),
.C(n_378),
.Y(n_7294)
);

OAI22xp33_ASAP7_75t_L g7295 ( 
.A1(n_6975),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_7295)
);

AOI22xp33_ASAP7_75t_L g7296 ( 
.A1(n_7154),
.A2(n_2387),
.B1(n_2393),
.B2(n_2371),
.Y(n_7296)
);

INVx2_ASAP7_75t_L g7297 ( 
.A(n_7000),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6960),
.Y(n_7298)
);

OAI21xp5_ASAP7_75t_L g7299 ( 
.A1(n_7120),
.A2(n_7138),
.B(n_6987),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_6965),
.Y(n_7300)
);

A2O1A1Ixp33_ASAP7_75t_L g7301 ( 
.A1(n_7167),
.A2(n_7145),
.B(n_6988),
.C(n_7147),
.Y(n_7301)
);

AOI22xp33_ASAP7_75t_L g7302 ( 
.A1(n_7125),
.A2(n_2393),
.B1(n_2401),
.B2(n_2387),
.Y(n_7302)
);

AND2x4_ASAP7_75t_L g7303 ( 
.A(n_7012),
.B(n_380),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6966),
.Y(n_7304)
);

AOI22xp33_ASAP7_75t_L g7305 ( 
.A1(n_7116),
.A2(n_2401),
.B1(n_2411),
.B2(n_2393),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6967),
.Y(n_7306)
);

NAND3xp33_ASAP7_75t_L g7307 ( 
.A(n_6976),
.B(n_381),
.C(n_382),
.Y(n_7307)
);

OAI22xp33_ASAP7_75t_L g7308 ( 
.A1(n_7165),
.A2(n_388),
.B1(n_382),
.B2(n_386),
.Y(n_7308)
);

OAI22xp5_ASAP7_75t_L g7309 ( 
.A1(n_7164),
.A2(n_389),
.B1(n_386),
.B2(n_388),
.Y(n_7309)
);

INVx2_ASAP7_75t_L g7310 ( 
.A(n_7012),
.Y(n_7310)
);

AOI22xp33_ASAP7_75t_L g7311 ( 
.A1(n_7105),
.A2(n_7107),
.B1(n_7106),
.B2(n_7029),
.Y(n_7311)
);

OAI22xp5_ASAP7_75t_L g7312 ( 
.A1(n_7164),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_7312)
);

CKINVDCx8_ASAP7_75t_R g7313 ( 
.A(n_7102),
.Y(n_7313)
);

OAI22xp5_ASAP7_75t_L g7314 ( 
.A1(n_7159),
.A2(n_395),
.B1(n_391),
.B2(n_393),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_6968),
.Y(n_7315)
);

OAI22xp5_ASAP7_75t_L g7316 ( 
.A1(n_7037),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_7316)
);

AOI22xp33_ASAP7_75t_L g7317 ( 
.A1(n_7022),
.A2(n_2411),
.B1(n_2412),
.B2(n_2401),
.Y(n_7317)
);

INVx1_ASAP7_75t_L g7318 ( 
.A(n_6970),
.Y(n_7318)
);

OAI22xp5_ASAP7_75t_L g7319 ( 
.A1(n_7118),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_7076),
.B(n_399),
.Y(n_7320)
);

OAI22xp5_ASAP7_75t_L g7321 ( 
.A1(n_7118),
.A2(n_7137),
.B1(n_7031),
.B2(n_7021),
.Y(n_7321)
);

AND2x4_ASAP7_75t_L g7322 ( 
.A(n_7042),
.B(n_400),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_6971),
.Y(n_7323)
);

AOI22xp33_ASAP7_75t_SL g7324 ( 
.A1(n_7111),
.A2(n_403),
.B1(n_400),
.B2(n_402),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_6977),
.Y(n_7325)
);

OAI22xp5_ASAP7_75t_L g7326 ( 
.A1(n_7137),
.A2(n_405),
.B1(n_402),
.B2(n_404),
.Y(n_7326)
);

AOI21xp33_ASAP7_75t_L g7327 ( 
.A1(n_6962),
.A2(n_406),
.B(n_407),
.Y(n_7327)
);

AOI22xp33_ASAP7_75t_L g7328 ( 
.A1(n_7145),
.A2(n_2411),
.B1(n_2412),
.B2(n_2401),
.Y(n_7328)
);

AOI22xp33_ASAP7_75t_L g7329 ( 
.A1(n_7158),
.A2(n_2411),
.B1(n_2412),
.B2(n_2401),
.Y(n_7329)
);

AOI22xp33_ASAP7_75t_L g7330 ( 
.A1(n_7161),
.A2(n_2412),
.B1(n_2415),
.B2(n_2411),
.Y(n_7330)
);

OR2x6_ASAP7_75t_L g7331 ( 
.A(n_6956),
.B(n_7100),
.Y(n_7331)
);

BUFx4f_ASAP7_75t_SL g7332 ( 
.A(n_6956),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6980),
.Y(n_7333)
);

AOI221xp5_ASAP7_75t_L g7334 ( 
.A1(n_6974),
.A2(n_7003),
.B1(n_7131),
.B2(n_7132),
.C(n_7028),
.Y(n_7334)
);

HB1xp67_ASAP7_75t_L g7335 ( 
.A(n_6953),
.Y(n_7335)
);

OAI22xp33_ASAP7_75t_L g7336 ( 
.A1(n_7165),
.A2(n_410),
.B1(n_406),
.B2(n_409),
.Y(n_7336)
);

NAND2xp5_ASAP7_75t_L g7337 ( 
.A(n_7156),
.B(n_410),
.Y(n_7337)
);

AOI22xp5_ASAP7_75t_L g7338 ( 
.A1(n_7038),
.A2(n_4070),
.B1(n_4049),
.B2(n_4003),
.Y(n_7338)
);

AOI22xp33_ASAP7_75t_SL g7339 ( 
.A1(n_7172),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_7339)
);

NOR2x1_ASAP7_75t_L g7340 ( 
.A(n_7101),
.B(n_412),
.Y(n_7340)
);

NAND3xp33_ASAP7_75t_SL g7341 ( 
.A(n_7097),
.B(n_413),
.C(n_415),
.Y(n_7341)
);

AOI22xp33_ASAP7_75t_L g7342 ( 
.A1(n_7038),
.A2(n_2415),
.B1(n_2412),
.B2(n_2247),
.Y(n_7342)
);

OAI21x1_ASAP7_75t_L g7343 ( 
.A1(n_7097),
.A2(n_6973),
.B(n_6985),
.Y(n_7343)
);

AOI22xp33_ASAP7_75t_L g7344 ( 
.A1(n_7027),
.A2(n_2415),
.B1(n_2247),
.B2(n_2278),
.Y(n_7344)
);

NOR2x1p5_ASAP7_75t_L g7345 ( 
.A(n_6984),
.B(n_417),
.Y(n_7345)
);

OAI21xp33_ASAP7_75t_L g7346 ( 
.A1(n_7060),
.A2(n_7003),
.B(n_6974),
.Y(n_7346)
);

A2O1A1Ixp33_ASAP7_75t_L g7347 ( 
.A1(n_7127),
.A2(n_419),
.B(n_417),
.C(n_418),
.Y(n_7347)
);

HB1xp67_ASAP7_75t_L g7348 ( 
.A(n_6953),
.Y(n_7348)
);

AOI22xp33_ASAP7_75t_L g7349 ( 
.A1(n_7007),
.A2(n_2415),
.B1(n_2278),
.B2(n_2326),
.Y(n_7349)
);

AOI21xp5_ASAP7_75t_L g7350 ( 
.A1(n_7101),
.A2(n_420),
.B(n_422),
.Y(n_7350)
);

AOI22xp5_ASAP7_75t_L g7351 ( 
.A1(n_6999),
.A2(n_4070),
.B1(n_4049),
.B2(n_4003),
.Y(n_7351)
);

OAI221xp5_ASAP7_75t_L g7352 ( 
.A1(n_7006),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.C(n_425),
.Y(n_7352)
);

NAND2x1p5_ASAP7_75t_L g7353 ( 
.A(n_7096),
.B(n_423),
.Y(n_7353)
);

AO31x2_ASAP7_75t_L g7354 ( 
.A1(n_6947),
.A2(n_428),
.A3(n_424),
.B(n_426),
.Y(n_7354)
);

BUFx2_ASAP7_75t_L g7355 ( 
.A(n_7016),
.Y(n_7355)
);

INVx4_ASAP7_75t_L g7356 ( 
.A(n_7112),
.Y(n_7356)
);

INVxp67_ASAP7_75t_L g7357 ( 
.A(n_7077),
.Y(n_7357)
);

AND2x2_ASAP7_75t_L g7358 ( 
.A(n_7203),
.B(n_7005),
.Y(n_7358)
);

OR2x2_ASAP7_75t_L g7359 ( 
.A(n_7288),
.B(n_7321),
.Y(n_7359)
);

BUFx3_ASAP7_75t_L g7360 ( 
.A(n_7313),
.Y(n_7360)
);

BUFx3_ASAP7_75t_L g7361 ( 
.A(n_7285),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_7213),
.Y(n_7362)
);

AND2x2_ASAP7_75t_L g7363 ( 
.A(n_7266),
.B(n_7014),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_7178),
.Y(n_7364)
);

OR2x2_ASAP7_75t_L g7365 ( 
.A(n_7193),
.B(n_7083),
.Y(n_7365)
);

AND2x4_ASAP7_75t_L g7366 ( 
.A(n_7237),
.B(n_7080),
.Y(n_7366)
);

BUFx3_ASAP7_75t_L g7367 ( 
.A(n_7222),
.Y(n_7367)
);

AND2x4_ASAP7_75t_L g7368 ( 
.A(n_7242),
.B(n_7245),
.Y(n_7368)
);

BUFx2_ASAP7_75t_L g7369 ( 
.A(n_7245),
.Y(n_7369)
);

INVx2_ASAP7_75t_L g7370 ( 
.A(n_7238),
.Y(n_7370)
);

AND2x2_ASAP7_75t_L g7371 ( 
.A(n_7209),
.B(n_7051),
.Y(n_7371)
);

INVx1_ASAP7_75t_L g7372 ( 
.A(n_7184),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_7238),
.Y(n_7373)
);

OR2x2_ASAP7_75t_L g7374 ( 
.A(n_7331),
.B(n_7083),
.Y(n_7374)
);

INVx1_ASAP7_75t_SL g7375 ( 
.A(n_7332),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_7292),
.Y(n_7376)
);

BUFx3_ASAP7_75t_L g7377 ( 
.A(n_7242),
.Y(n_7377)
);

OR2x2_ASAP7_75t_L g7378 ( 
.A(n_7331),
.B(n_7068),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_7192),
.Y(n_7379)
);

AND2x4_ASAP7_75t_L g7380 ( 
.A(n_7262),
.B(n_7081),
.Y(n_7380)
);

AND2x2_ASAP7_75t_L g7381 ( 
.A(n_7271),
.B(n_7082),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_7173),
.B(n_7091),
.Y(n_7382)
);

AND2x2_ASAP7_75t_L g7383 ( 
.A(n_7273),
.B(n_7094),
.Y(n_7383)
);

AND2x2_ASAP7_75t_L g7384 ( 
.A(n_7356),
.B(n_7103),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_7200),
.Y(n_7385)
);

INVx1_ASAP7_75t_SL g7386 ( 
.A(n_7268),
.Y(n_7386)
);

OR2x2_ASAP7_75t_L g7387 ( 
.A(n_7214),
.B(n_7069),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_7205),
.Y(n_7388)
);

INVx3_ASAP7_75t_L g7389 ( 
.A(n_7356),
.Y(n_7389)
);

NAND2xp5_ASAP7_75t_L g7390 ( 
.A(n_7340),
.B(n_7357),
.Y(n_7390)
);

AND2x2_ASAP7_75t_L g7391 ( 
.A(n_7284),
.B(n_7048),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_7355),
.Y(n_7392)
);

AND2x2_ASAP7_75t_L g7393 ( 
.A(n_7297),
.B(n_7070),
.Y(n_7393)
);

INVx2_ASAP7_75t_L g7394 ( 
.A(n_7226),
.Y(n_7394)
);

HB1xp67_ASAP7_75t_L g7395 ( 
.A(n_7335),
.Y(n_7395)
);

INVx2_ASAP7_75t_SL g7396 ( 
.A(n_7303),
.Y(n_7396)
);

HB1xp67_ASAP7_75t_L g7397 ( 
.A(n_7348),
.Y(n_7397)
);

INVx3_ASAP7_75t_L g7398 ( 
.A(n_7303),
.Y(n_7398)
);

BUFx3_ASAP7_75t_L g7399 ( 
.A(n_7216),
.Y(n_7399)
);

NAND2x1_ASAP7_75t_L g7400 ( 
.A(n_7194),
.B(n_6979),
.Y(n_7400)
);

AND2x2_ASAP7_75t_L g7401 ( 
.A(n_7310),
.B(n_7074),
.Y(n_7401)
);

AND2x2_ASAP7_75t_L g7402 ( 
.A(n_7234),
.B(n_7079),
.Y(n_7402)
);

AND2x4_ASAP7_75t_SL g7403 ( 
.A(n_7243),
.B(n_7075),
.Y(n_7403)
);

AND2x2_ASAP7_75t_L g7404 ( 
.A(n_7224),
.B(n_7084),
.Y(n_7404)
);

INVx2_ASAP7_75t_L g7405 ( 
.A(n_7253),
.Y(n_7405)
);

AND2x2_ASAP7_75t_L g7406 ( 
.A(n_7229),
.B(n_7087),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_7272),
.Y(n_7407)
);

AND2x2_ASAP7_75t_L g7408 ( 
.A(n_7217),
.B(n_7090),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_7227),
.Y(n_7409)
);

INVx1_ASAP7_75t_L g7410 ( 
.A(n_7252),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_7260),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_7263),
.Y(n_7412)
);

AND2x2_ASAP7_75t_L g7413 ( 
.A(n_7187),
.B(n_7126),
.Y(n_7413)
);

INVx2_ASAP7_75t_L g7414 ( 
.A(n_7227),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_7264),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_7278),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7291),
.Y(n_7417)
);

BUFx3_ASAP7_75t_L g7418 ( 
.A(n_7216),
.Y(n_7418)
);

AOI21xp33_ASAP7_75t_L g7419 ( 
.A1(n_7198),
.A2(n_7053),
.B(n_7172),
.Y(n_7419)
);

AND2x4_ASAP7_75t_L g7420 ( 
.A(n_7322),
.B(n_6979),
.Y(n_7420)
);

INVx2_ASAP7_75t_L g7421 ( 
.A(n_7253),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_7298),
.Y(n_7422)
);

OR2x2_ASAP7_75t_L g7423 ( 
.A(n_7188),
.B(n_7007),
.Y(n_7423)
);

BUFx3_ASAP7_75t_L g7424 ( 
.A(n_7322),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_7300),
.Y(n_7425)
);

AND2x2_ASAP7_75t_L g7426 ( 
.A(n_7256),
.B(n_7146),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_7304),
.Y(n_7427)
);

INVx2_ASAP7_75t_L g7428 ( 
.A(n_7227),
.Y(n_7428)
);

BUFx2_ASAP7_75t_L g7429 ( 
.A(n_7211),
.Y(n_7429)
);

INVx2_ASAP7_75t_L g7430 ( 
.A(n_7235),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_7306),
.Y(n_7431)
);

INVx3_ASAP7_75t_L g7432 ( 
.A(n_7194),
.Y(n_7432)
);

HB1xp67_ASAP7_75t_L g7433 ( 
.A(n_7206),
.Y(n_7433)
);

AND2x2_ASAP7_75t_L g7434 ( 
.A(n_7258),
.B(n_7016),
.Y(n_7434)
);

BUFx2_ASAP7_75t_L g7435 ( 
.A(n_7196),
.Y(n_7435)
);

INVx3_ASAP7_75t_L g7436 ( 
.A(n_7199),
.Y(n_7436)
);

AND2x2_ASAP7_75t_L g7437 ( 
.A(n_7345),
.B(n_7104),
.Y(n_7437)
);

INVx1_ASAP7_75t_L g7438 ( 
.A(n_7315),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_7318),
.Y(n_7439)
);

INVx2_ASAP7_75t_L g7440 ( 
.A(n_7354),
.Y(n_7440)
);

INVx2_ASAP7_75t_SL g7441 ( 
.A(n_7353),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_7323),
.Y(n_7442)
);

INVx2_ASAP7_75t_L g7443 ( 
.A(n_7354),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_7325),
.Y(n_7444)
);

INVx2_ASAP7_75t_L g7445 ( 
.A(n_7354),
.Y(n_7445)
);

INVx2_ASAP7_75t_L g7446 ( 
.A(n_7343),
.Y(n_7446)
);

INVx2_ASAP7_75t_SL g7447 ( 
.A(n_7225),
.Y(n_7447)
);

HB1xp67_ASAP7_75t_L g7448 ( 
.A(n_7246),
.Y(n_7448)
);

OR2x2_ASAP7_75t_L g7449 ( 
.A(n_7231),
.B(n_7148),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_7333),
.Y(n_7450)
);

AND2x4_ASAP7_75t_L g7451 ( 
.A(n_7250),
.B(n_7140),
.Y(n_7451)
);

INVx3_ASAP7_75t_L g7452 ( 
.A(n_7197),
.Y(n_7452)
);

AND2x2_ASAP7_75t_L g7453 ( 
.A(n_7311),
.B(n_7124),
.Y(n_7453)
);

AND2x4_ASAP7_75t_L g7454 ( 
.A(n_7210),
.B(n_7142),
.Y(n_7454)
);

INVx2_ASAP7_75t_L g7455 ( 
.A(n_7275),
.Y(n_7455)
);

AND2x2_ASAP7_75t_L g7456 ( 
.A(n_7301),
.B(n_7170),
.Y(n_7456)
);

NAND2xp5_ASAP7_75t_L g7457 ( 
.A(n_7334),
.B(n_6983),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_L g7458 ( 
.A(n_7218),
.B(n_6986),
.Y(n_7458)
);

INVx2_ASAP7_75t_L g7459 ( 
.A(n_7219),
.Y(n_7459)
);

OR2x6_ASAP7_75t_L g7460 ( 
.A(n_7204),
.B(n_7061),
.Y(n_7460)
);

AND2x2_ASAP7_75t_L g7461 ( 
.A(n_7293),
.B(n_7036),
.Y(n_7461)
);

AND2x4_ASAP7_75t_L g7462 ( 
.A(n_7299),
.B(n_7045),
.Y(n_7462)
);

AND2x2_ASAP7_75t_L g7463 ( 
.A(n_7175),
.B(n_7065),
.Y(n_7463)
);

INVx1_ASAP7_75t_L g7464 ( 
.A(n_7320),
.Y(n_7464)
);

INVx1_ASAP7_75t_L g7465 ( 
.A(n_7248),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_7212),
.B(n_7077),
.Y(n_7466)
);

INVx2_ASAP7_75t_SL g7467 ( 
.A(n_7337),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_7215),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_7319),
.Y(n_7469)
);

INVx2_ASAP7_75t_L g7470 ( 
.A(n_7181),
.Y(n_7470)
);

AND2x2_ASAP7_75t_L g7471 ( 
.A(n_7283),
.B(n_7177),
.Y(n_7471)
);

BUFx2_ASAP7_75t_L g7472 ( 
.A(n_7307),
.Y(n_7472)
);

OR2x2_ASAP7_75t_L g7473 ( 
.A(n_7244),
.B(n_7061),
.Y(n_7473)
);

OR2x2_ASAP7_75t_L g7474 ( 
.A(n_7341),
.B(n_7255),
.Y(n_7474)
);

INVx2_ASAP7_75t_L g7475 ( 
.A(n_7186),
.Y(n_7475)
);

AND2x2_ASAP7_75t_L g7476 ( 
.A(n_7174),
.B(n_7039),
.Y(n_7476)
);

OR2x2_ASAP7_75t_L g7477 ( 
.A(n_7223),
.B(n_7089),
.Y(n_7477)
);

OR2x2_ASAP7_75t_L g7478 ( 
.A(n_7350),
.B(n_7089),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_7346),
.Y(n_7479)
);

AND2x2_ASAP7_75t_L g7480 ( 
.A(n_7236),
.B(n_7049),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_L g7481 ( 
.A(n_7195),
.B(n_7024),
.Y(n_7481)
);

AND2x2_ASAP7_75t_L g7482 ( 
.A(n_7281),
.B(n_7054),
.Y(n_7482)
);

INVxp67_ASAP7_75t_SL g7483 ( 
.A(n_7207),
.Y(n_7483)
);

AND2x2_ASAP7_75t_L g7484 ( 
.A(n_7327),
.B(n_7058),
.Y(n_7484)
);

AO31x2_ASAP7_75t_L g7485 ( 
.A1(n_7176),
.A2(n_7046),
.A3(n_7063),
.B(n_7055),
.Y(n_7485)
);

NAND2x1p5_ASAP7_75t_L g7486 ( 
.A(n_7208),
.B(n_6949),
.Y(n_7486)
);

AND2x2_ASAP7_75t_L g7487 ( 
.A(n_7324),
.B(n_7059),
.Y(n_7487)
);

AND2x2_ASAP7_75t_L g7488 ( 
.A(n_7180),
.B(n_7025),
.Y(n_7488)
);

INVx2_ASAP7_75t_L g7489 ( 
.A(n_7183),
.Y(n_7489)
);

AND2x2_ASAP7_75t_L g7490 ( 
.A(n_7201),
.B(n_7088),
.Y(n_7490)
);

NAND2xp5_ASAP7_75t_L g7491 ( 
.A(n_7274),
.B(n_6947),
.Y(n_7491)
);

INVx2_ASAP7_75t_L g7492 ( 
.A(n_7179),
.Y(n_7492)
);

HB1xp67_ASAP7_75t_L g7493 ( 
.A(n_7289),
.Y(n_7493)
);

HB1xp67_ASAP7_75t_L g7494 ( 
.A(n_7261),
.Y(n_7494)
);

AND2x2_ASAP7_75t_L g7495 ( 
.A(n_7240),
.B(n_7088),
.Y(n_7495)
);

INVxp67_ASAP7_75t_SL g7496 ( 
.A(n_7308),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7276),
.Y(n_7497)
);

BUFx2_ASAP7_75t_L g7498 ( 
.A(n_7232),
.Y(n_7498)
);

AND2x2_ASAP7_75t_L g7499 ( 
.A(n_7185),
.B(n_7008),
.Y(n_7499)
);

AND2x2_ASAP7_75t_L g7500 ( 
.A(n_7287),
.B(n_7128),
.Y(n_7500)
);

INVx1_ASAP7_75t_SL g7501 ( 
.A(n_7290),
.Y(n_7501)
);

AND2x2_ASAP7_75t_L g7502 ( 
.A(n_7375),
.B(n_7071),
.Y(n_7502)
);

AND2x2_ASAP7_75t_L g7503 ( 
.A(n_7375),
.B(n_6948),
.Y(n_7503)
);

INVx2_ASAP7_75t_L g7504 ( 
.A(n_7367),
.Y(n_7504)
);

OR2x2_ASAP7_75t_L g7505 ( 
.A(n_7386),
.B(n_7309),
.Y(n_7505)
);

INVx1_ASAP7_75t_L g7506 ( 
.A(n_7395),
.Y(n_7506)
);

OR2x2_ASAP7_75t_L g7507 ( 
.A(n_7386),
.B(n_7312),
.Y(n_7507)
);

INVx1_ASAP7_75t_L g7508 ( 
.A(n_7395),
.Y(n_7508)
);

NAND2xp5_ASAP7_75t_L g7509 ( 
.A(n_7493),
.B(n_6948),
.Y(n_7509)
);

INVx1_ASAP7_75t_SL g7510 ( 
.A(n_7435),
.Y(n_7510)
);

INVx4_ASAP7_75t_L g7511 ( 
.A(n_7367),
.Y(n_7511)
);

AND2x2_ASAP7_75t_L g7512 ( 
.A(n_7360),
.B(n_7157),
.Y(n_7512)
);

AND2x2_ASAP7_75t_L g7513 ( 
.A(n_7360),
.B(n_7163),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7397),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7397),
.Y(n_7515)
);

AND2x2_ASAP7_75t_L g7516 ( 
.A(n_7371),
.B(n_7143),
.Y(n_7516)
);

AND2x2_ASAP7_75t_L g7517 ( 
.A(n_7391),
.B(n_7286),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7392),
.Y(n_7518)
);

AND2x4_ASAP7_75t_L g7519 ( 
.A(n_7420),
.B(n_7166),
.Y(n_7519)
);

OR2x2_ASAP7_75t_L g7520 ( 
.A(n_7359),
.B(n_7326),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7392),
.Y(n_7521)
);

AND2x2_ASAP7_75t_L g7522 ( 
.A(n_7361),
.B(n_7358),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7362),
.Y(n_7523)
);

BUFx2_ASAP7_75t_L g7524 ( 
.A(n_7424),
.Y(n_7524)
);

BUFx2_ASAP7_75t_L g7525 ( 
.A(n_7424),
.Y(n_7525)
);

HB1xp67_ASAP7_75t_L g7526 ( 
.A(n_7399),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7394),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7394),
.Y(n_7528)
);

AND2x2_ASAP7_75t_L g7529 ( 
.A(n_7361),
.B(n_7369),
.Y(n_7529)
);

NOR2x1_ASAP7_75t_L g7530 ( 
.A(n_7370),
.B(n_7373),
.Y(n_7530)
);

HB1xp67_ASAP7_75t_L g7531 ( 
.A(n_7399),
.Y(n_7531)
);

AND2x4_ASAP7_75t_L g7532 ( 
.A(n_7420),
.B(n_7418),
.Y(n_7532)
);

AND2x2_ASAP7_75t_L g7533 ( 
.A(n_7363),
.B(n_7166),
.Y(n_7533)
);

NAND2xp5_ASAP7_75t_L g7534 ( 
.A(n_7493),
.B(n_7269),
.Y(n_7534)
);

AND2x2_ASAP7_75t_L g7535 ( 
.A(n_7437),
.B(n_7403),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7429),
.Y(n_7536)
);

INVx2_ASAP7_75t_L g7537 ( 
.A(n_7400),
.Y(n_7537)
);

INVx2_ASAP7_75t_L g7538 ( 
.A(n_7432),
.Y(n_7538)
);

NAND2xp5_ASAP7_75t_L g7539 ( 
.A(n_7501),
.B(n_7277),
.Y(n_7539)
);

BUFx3_ASAP7_75t_L g7540 ( 
.A(n_7418),
.Y(n_7540)
);

INVx2_ASAP7_75t_L g7541 ( 
.A(n_7432),
.Y(n_7541)
);

HB1xp67_ASAP7_75t_L g7542 ( 
.A(n_7398),
.Y(n_7542)
);

OR2x2_ASAP7_75t_L g7543 ( 
.A(n_7473),
.B(n_7347),
.Y(n_7543)
);

INVx2_ASAP7_75t_L g7544 ( 
.A(n_7398),
.Y(n_7544)
);

AND2x2_ASAP7_75t_L g7545 ( 
.A(n_7403),
.B(n_7267),
.Y(n_7545)
);

NAND3xp33_ASAP7_75t_L g7546 ( 
.A(n_7390),
.B(n_7239),
.C(n_7241),
.Y(n_7546)
);

NAND2xp5_ASAP7_75t_L g7547 ( 
.A(n_7501),
.B(n_7336),
.Y(n_7547)
);

INVx2_ASAP7_75t_L g7548 ( 
.A(n_7377),
.Y(n_7548)
);

AND2x2_ASAP7_75t_L g7549 ( 
.A(n_7368),
.B(n_7110),
.Y(n_7549)
);

OAI222xp33_ASAP7_75t_L g7550 ( 
.A1(n_7466),
.A2(n_7491),
.B1(n_7486),
.B2(n_7472),
.C1(n_7474),
.C2(n_7461),
.Y(n_7550)
);

INVxp67_ASAP7_75t_L g7551 ( 
.A(n_7390),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7365),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_7377),
.Y(n_7553)
);

AND2x4_ASAP7_75t_SL g7554 ( 
.A(n_7368),
.B(n_7338),
.Y(n_7554)
);

INVx4_ASAP7_75t_L g7555 ( 
.A(n_7389),
.Y(n_7555)
);

AND2x2_ASAP7_75t_L g7556 ( 
.A(n_7396),
.B(n_7110),
.Y(n_7556)
);

INVxp67_ASAP7_75t_SL g7557 ( 
.A(n_7452),
.Y(n_7557)
);

INVx2_ASAP7_75t_L g7558 ( 
.A(n_7389),
.Y(n_7558)
);

INVx1_ASAP7_75t_L g7559 ( 
.A(n_7370),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7374),
.Y(n_7560)
);

NOR2x1_ASAP7_75t_SL g7561 ( 
.A(n_7441),
.B(n_6996),
.Y(n_7561)
);

NAND2xp5_ASAP7_75t_L g7562 ( 
.A(n_7433),
.B(n_7339),
.Y(n_7562)
);

NOR2xp33_ASAP7_75t_L g7563 ( 
.A(n_7436),
.B(n_7352),
.Y(n_7563)
);

INVx2_ASAP7_75t_L g7564 ( 
.A(n_7366),
.Y(n_7564)
);

INVx1_ASAP7_75t_L g7565 ( 
.A(n_7373),
.Y(n_7565)
);

INVx1_ASAP7_75t_L g7566 ( 
.A(n_7407),
.Y(n_7566)
);

NAND2xp5_ASAP7_75t_L g7567 ( 
.A(n_7433),
.B(n_7280),
.Y(n_7567)
);

AND2x2_ASAP7_75t_L g7568 ( 
.A(n_7366),
.B(n_7382),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_7364),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_7372),
.Y(n_7570)
);

NAND2xp5_ASAP7_75t_L g7571 ( 
.A(n_7496),
.B(n_7448),
.Y(n_7571)
);

AND2x2_ASAP7_75t_L g7572 ( 
.A(n_7436),
.B(n_6954),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7405),
.Y(n_7573)
);

AND2x2_ASAP7_75t_L g7574 ( 
.A(n_7404),
.B(n_6954),
.Y(n_7574)
);

HB1xp67_ASAP7_75t_L g7575 ( 
.A(n_7451),
.Y(n_7575)
);

AND2x2_ASAP7_75t_L g7576 ( 
.A(n_7406),
.B(n_6954),
.Y(n_7576)
);

AND2x2_ASAP7_75t_L g7577 ( 
.A(n_7413),
.B(n_7149),
.Y(n_7577)
);

AND2x2_ASAP7_75t_L g7578 ( 
.A(n_7421),
.B(n_7149),
.Y(n_7578)
);

OAI22xp5_ASAP7_75t_L g7579 ( 
.A1(n_7466),
.A2(n_7220),
.B1(n_7202),
.B2(n_7254),
.Y(n_7579)
);

AND2x2_ASAP7_75t_L g7580 ( 
.A(n_7408),
.B(n_6944),
.Y(n_7580)
);

NAND2xp5_ASAP7_75t_L g7581 ( 
.A(n_7496),
.B(n_7282),
.Y(n_7581)
);

INVx1_ASAP7_75t_L g7582 ( 
.A(n_7409),
.Y(n_7582)
);

AOI22xp33_ASAP7_75t_L g7583 ( 
.A1(n_7471),
.A2(n_7190),
.B1(n_7191),
.B2(n_7189),
.Y(n_7583)
);

AND2x2_ASAP7_75t_L g7584 ( 
.A(n_7426),
.B(n_6945),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_7409),
.Y(n_7585)
);

NAND2xp5_ASAP7_75t_L g7586 ( 
.A(n_7448),
.B(n_7295),
.Y(n_7586)
);

BUFx6f_ASAP7_75t_L g7587 ( 
.A(n_7414),
.Y(n_7587)
);

INVx1_ASAP7_75t_L g7588 ( 
.A(n_7414),
.Y(n_7588)
);

OR2x2_ASAP7_75t_L g7589 ( 
.A(n_7387),
.B(n_7316),
.Y(n_7589)
);

AND2x4_ASAP7_75t_L g7590 ( 
.A(n_7428),
.B(n_6952),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7428),
.Y(n_7591)
);

AOI22xp33_ASAP7_75t_SL g7592 ( 
.A1(n_7463),
.A2(n_7294),
.B1(n_7314),
.B2(n_6997),
.Y(n_7592)
);

AND2x2_ASAP7_75t_L g7593 ( 
.A(n_7383),
.B(n_7381),
.Y(n_7593)
);

NAND4xp25_ASAP7_75t_L g7594 ( 
.A(n_7376),
.B(n_7221),
.C(n_7228),
.D(n_7296),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_7440),
.Y(n_7595)
);

INVx1_ASAP7_75t_SL g7596 ( 
.A(n_7434),
.Y(n_7596)
);

BUFx2_ASAP7_75t_L g7597 ( 
.A(n_7451),
.Y(n_7597)
);

NAND2xp5_ASAP7_75t_L g7598 ( 
.A(n_7483),
.B(n_7182),
.Y(n_7598)
);

AOI221xp5_ASAP7_75t_L g7599 ( 
.A1(n_7419),
.A2(n_7160),
.B1(n_6997),
.B2(n_6996),
.C(n_7233),
.Y(n_7599)
);

NAND2xp5_ASAP7_75t_L g7600 ( 
.A(n_7483),
.B(n_7160),
.Y(n_7600)
);

OAI22xp5_ASAP7_75t_L g7601 ( 
.A1(n_7494),
.A2(n_7328),
.B1(n_7349),
.B2(n_6964),
.Y(n_7601)
);

BUFx2_ASAP7_75t_L g7602 ( 
.A(n_7380),
.Y(n_7602)
);

INVx4_ASAP7_75t_SL g7603 ( 
.A(n_7384),
.Y(n_7603)
);

AND2x2_ASAP7_75t_L g7604 ( 
.A(n_7453),
.B(n_6963),
.Y(n_7604)
);

INVx2_ASAP7_75t_L g7605 ( 
.A(n_7378),
.Y(n_7605)
);

INVx1_ASAP7_75t_L g7606 ( 
.A(n_7440),
.Y(n_7606)
);

INVx2_ASAP7_75t_L g7607 ( 
.A(n_7380),
.Y(n_7607)
);

NAND2xp5_ASAP7_75t_L g7608 ( 
.A(n_7494),
.B(n_7500),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_7443),
.Y(n_7609)
);

OR2x2_ASAP7_75t_L g7610 ( 
.A(n_7478),
.B(n_7469),
.Y(n_7610)
);

INVx2_ASAP7_75t_L g7611 ( 
.A(n_7452),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_7443),
.Y(n_7612)
);

INVx2_ASAP7_75t_L g7613 ( 
.A(n_7402),
.Y(n_7613)
);

AND2x2_ASAP7_75t_L g7614 ( 
.A(n_7495),
.B(n_6982),
.Y(n_7614)
);

AND2x4_ASAP7_75t_L g7615 ( 
.A(n_7393),
.B(n_7305),
.Y(n_7615)
);

HB1xp67_ASAP7_75t_L g7616 ( 
.A(n_7430),
.Y(n_7616)
);

AND2x4_ASAP7_75t_L g7617 ( 
.A(n_7401),
.B(n_7265),
.Y(n_7617)
);

NOR2xp67_ASAP7_75t_L g7618 ( 
.A(n_7430),
.B(n_7423),
.Y(n_7618)
);

AND2x2_ASAP7_75t_L g7619 ( 
.A(n_7482),
.B(n_7249),
.Y(n_7619)
);

INVx1_ASAP7_75t_L g7620 ( 
.A(n_7445),
.Y(n_7620)
);

INVx2_ASAP7_75t_L g7621 ( 
.A(n_7454),
.Y(n_7621)
);

NAND2xp5_ASAP7_75t_L g7622 ( 
.A(n_7491),
.B(n_7251),
.Y(n_7622)
);

AND2x2_ASAP7_75t_L g7623 ( 
.A(n_7487),
.B(n_7302),
.Y(n_7623)
);

AOI22xp33_ASAP7_75t_L g7624 ( 
.A1(n_7489),
.A2(n_7257),
.B1(n_7259),
.B2(n_7247),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7445),
.Y(n_7625)
);

INVx1_ASAP7_75t_L g7626 ( 
.A(n_7459),
.Y(n_7626)
);

AND2x2_ASAP7_75t_L g7627 ( 
.A(n_7456),
.B(n_7317),
.Y(n_7627)
);

INVx3_ASAP7_75t_L g7628 ( 
.A(n_7454),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7459),
.Y(n_7629)
);

AND2x2_ASAP7_75t_L g7630 ( 
.A(n_7447),
.B(n_7279),
.Y(n_7630)
);

AOI22xp33_ASAP7_75t_L g7631 ( 
.A1(n_7489),
.A2(n_7329),
.B1(n_7330),
.B2(n_7270),
.Y(n_7631)
);

INVx2_ASAP7_75t_L g7632 ( 
.A(n_7446),
.Y(n_7632)
);

INVx1_ASAP7_75t_L g7633 ( 
.A(n_7379),
.Y(n_7633)
);

AND2x2_ASAP7_75t_L g7634 ( 
.A(n_7476),
.B(n_7351),
.Y(n_7634)
);

CKINVDCx5p33_ASAP7_75t_R g7635 ( 
.A(n_7460),
.Y(n_7635)
);

HB1xp67_ASAP7_75t_L g7636 ( 
.A(n_7460),
.Y(n_7636)
);

INVx2_ASAP7_75t_L g7637 ( 
.A(n_7446),
.Y(n_7637)
);

AOI22xp33_ASAP7_75t_L g7638 ( 
.A1(n_7492),
.A2(n_7230),
.B1(n_7342),
.B2(n_7344),
.Y(n_7638)
);

AND2x2_ASAP7_75t_L g7639 ( 
.A(n_7455),
.B(n_7099),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_7385),
.Y(n_7640)
);

AND2x2_ASAP7_75t_L g7641 ( 
.A(n_7522),
.B(n_7468),
.Y(n_7641)
);

INVx2_ASAP7_75t_L g7642 ( 
.A(n_7561),
.Y(n_7642)
);

AND2x2_ASAP7_75t_L g7643 ( 
.A(n_7535),
.B(n_7497),
.Y(n_7643)
);

AND2x2_ASAP7_75t_L g7644 ( 
.A(n_7511),
.B(n_7484),
.Y(n_7644)
);

INVxp67_ASAP7_75t_SL g7645 ( 
.A(n_7575),
.Y(n_7645)
);

INVx2_ASAP7_75t_L g7646 ( 
.A(n_7602),
.Y(n_7646)
);

NAND2xp5_ASAP7_75t_L g7647 ( 
.A(n_7510),
.B(n_7479),
.Y(n_7647)
);

AND2x2_ASAP7_75t_L g7648 ( 
.A(n_7511),
.B(n_7480),
.Y(n_7648)
);

NAND2xp5_ASAP7_75t_L g7649 ( 
.A(n_7510),
.B(n_7457),
.Y(n_7649)
);

AND2x4_ASAP7_75t_L g7650 ( 
.A(n_7603),
.B(n_7467),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_7542),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_L g7652 ( 
.A(n_7534),
.B(n_7457),
.Y(n_7652)
);

OR2x2_ASAP7_75t_L g7653 ( 
.A(n_7571),
.B(n_7449),
.Y(n_7653)
);

NAND2xp5_ASAP7_75t_L g7654 ( 
.A(n_7534),
.B(n_7481),
.Y(n_7654)
);

BUFx2_ASAP7_75t_L g7655 ( 
.A(n_7597),
.Y(n_7655)
);

INVx2_ASAP7_75t_L g7656 ( 
.A(n_7603),
.Y(n_7656)
);

NAND2xp5_ASAP7_75t_L g7657 ( 
.A(n_7526),
.B(n_7481),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7531),
.Y(n_7658)
);

AND2x4_ASAP7_75t_L g7659 ( 
.A(n_7532),
.B(n_7388),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7506),
.Y(n_7660)
);

NAND4xp75_ASAP7_75t_L g7661 ( 
.A(n_7530),
.B(n_7419),
.C(n_7475),
.D(n_7470),
.Y(n_7661)
);

INVx1_ASAP7_75t_L g7662 ( 
.A(n_7508),
.Y(n_7662)
);

AND2x2_ASAP7_75t_L g7663 ( 
.A(n_7529),
.B(n_7455),
.Y(n_7663)
);

NAND2xp5_ASAP7_75t_SL g7664 ( 
.A(n_7635),
.B(n_7486),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7514),
.Y(n_7665)
);

INVx2_ASAP7_75t_L g7666 ( 
.A(n_7532),
.Y(n_7666)
);

INVx1_ASAP7_75t_L g7667 ( 
.A(n_7515),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_7524),
.Y(n_7668)
);

AND2x2_ASAP7_75t_L g7669 ( 
.A(n_7568),
.B(n_7464),
.Y(n_7669)
);

OR2x6_ASAP7_75t_SL g7670 ( 
.A(n_7571),
.B(n_7477),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_7525),
.Y(n_7671)
);

NAND2xp5_ASAP7_75t_L g7672 ( 
.A(n_7579),
.B(n_7492),
.Y(n_7672)
);

OR2x2_ASAP7_75t_L g7673 ( 
.A(n_7610),
.B(n_7458),
.Y(n_7673)
);

HB1xp67_ASAP7_75t_L g7674 ( 
.A(n_7519),
.Y(n_7674)
);

OR2x2_ASAP7_75t_L g7675 ( 
.A(n_7505),
.B(n_7458),
.Y(n_7675)
);

NAND2xp5_ASAP7_75t_L g7676 ( 
.A(n_7579),
.B(n_7410),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7557),
.Y(n_7677)
);

NAND2xp5_ASAP7_75t_L g7678 ( 
.A(n_7587),
.B(n_7411),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_7587),
.Y(n_7679)
);

OR2x2_ASAP7_75t_L g7680 ( 
.A(n_7507),
.B(n_7460),
.Y(n_7680)
);

BUFx2_ASAP7_75t_L g7681 ( 
.A(n_7519),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_7587),
.Y(n_7682)
);

NAND2xp5_ASAP7_75t_L g7683 ( 
.A(n_7608),
.B(n_7412),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_7616),
.Y(n_7684)
);

AND2x2_ASAP7_75t_L g7685 ( 
.A(n_7504),
.B(n_7470),
.Y(n_7685)
);

INVx1_ASAP7_75t_L g7686 ( 
.A(n_7518),
.Y(n_7686)
);

INVxp67_ASAP7_75t_L g7687 ( 
.A(n_7636),
.Y(n_7687)
);

AND2x4_ASAP7_75t_L g7688 ( 
.A(n_7537),
.B(n_7415),
.Y(n_7688)
);

AND2x2_ASAP7_75t_L g7689 ( 
.A(n_7545),
.B(n_7498),
.Y(n_7689)
);

INVx2_ASAP7_75t_L g7690 ( 
.A(n_7540),
.Y(n_7690)
);

INVx3_ASAP7_75t_L g7691 ( 
.A(n_7555),
.Y(n_7691)
);

AND2x2_ASAP7_75t_L g7692 ( 
.A(n_7560),
.B(n_7475),
.Y(n_7692)
);

HB1xp67_ASAP7_75t_L g7693 ( 
.A(n_7628),
.Y(n_7693)
);

OR2x2_ASAP7_75t_L g7694 ( 
.A(n_7544),
.B(n_7488),
.Y(n_7694)
);

AND2x2_ASAP7_75t_L g7695 ( 
.A(n_7593),
.B(n_7462),
.Y(n_7695)
);

NOR2xp33_ASAP7_75t_L g7696 ( 
.A(n_7550),
.B(n_7416),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7521),
.Y(n_7697)
);

AND2x2_ASAP7_75t_L g7698 ( 
.A(n_7564),
.B(n_7462),
.Y(n_7698)
);

BUFx2_ASAP7_75t_L g7699 ( 
.A(n_7555),
.Y(n_7699)
);

AND2x4_ASAP7_75t_L g7700 ( 
.A(n_7538),
.B(n_7417),
.Y(n_7700)
);

NOR2x1p5_ASAP7_75t_L g7701 ( 
.A(n_7628),
.B(n_7422),
.Y(n_7701)
);

OR2x2_ASAP7_75t_L g7702 ( 
.A(n_7586),
.B(n_7465),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7595),
.Y(n_7703)
);

NAND2xp5_ASAP7_75t_L g7704 ( 
.A(n_7608),
.B(n_7425),
.Y(n_7704)
);

AND2x2_ASAP7_75t_L g7705 ( 
.A(n_7533),
.B(n_7605),
.Y(n_7705)
);

AND2x4_ASAP7_75t_L g7706 ( 
.A(n_7541),
.B(n_7427),
.Y(n_7706)
);

INVx2_ASAP7_75t_L g7707 ( 
.A(n_7611),
.Y(n_7707)
);

INVx2_ASAP7_75t_L g7708 ( 
.A(n_7548),
.Y(n_7708)
);

AND2x2_ASAP7_75t_L g7709 ( 
.A(n_7553),
.B(n_7431),
.Y(n_7709)
);

INVx1_ASAP7_75t_SL g7710 ( 
.A(n_7596),
.Y(n_7710)
);

INVx2_ASAP7_75t_L g7711 ( 
.A(n_7607),
.Y(n_7711)
);

INVx2_ASAP7_75t_L g7712 ( 
.A(n_7558),
.Y(n_7712)
);

INVxp67_ASAP7_75t_L g7713 ( 
.A(n_7517),
.Y(n_7713)
);

HB1xp67_ASAP7_75t_L g7714 ( 
.A(n_7618),
.Y(n_7714)
);

AND2x4_ASAP7_75t_L g7715 ( 
.A(n_7536),
.B(n_7438),
.Y(n_7715)
);

AND2x2_ASAP7_75t_L g7716 ( 
.A(n_7513),
.B(n_7439),
.Y(n_7716)
);

BUFx3_ASAP7_75t_L g7717 ( 
.A(n_7502),
.Y(n_7717)
);

INVx1_ASAP7_75t_SL g7718 ( 
.A(n_7596),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_7606),
.Y(n_7719)
);

NAND2xp5_ASAP7_75t_L g7720 ( 
.A(n_7539),
.B(n_7442),
.Y(n_7720)
);

INVx2_ASAP7_75t_L g7721 ( 
.A(n_7577),
.Y(n_7721)
);

INVx2_ASAP7_75t_L g7722 ( 
.A(n_7590),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_SL g7723 ( 
.A(n_7592),
.B(n_7499),
.Y(n_7723)
);

INVx2_ASAP7_75t_SL g7724 ( 
.A(n_7578),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_L g7725 ( 
.A(n_7539),
.B(n_7444),
.Y(n_7725)
);

INVx1_ASAP7_75t_L g7726 ( 
.A(n_7609),
.Y(n_7726)
);

INVx6_ASAP7_75t_L g7727 ( 
.A(n_7590),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_7612),
.Y(n_7728)
);

AND2x2_ASAP7_75t_L g7729 ( 
.A(n_7512),
.B(n_7503),
.Y(n_7729)
);

INVx5_ASAP7_75t_L g7730 ( 
.A(n_7549),
.Y(n_7730)
);

INVx1_ASAP7_75t_L g7731 ( 
.A(n_7620),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7625),
.Y(n_7732)
);

INVx2_ASAP7_75t_L g7733 ( 
.A(n_7556),
.Y(n_7733)
);

INVx1_ASAP7_75t_L g7734 ( 
.A(n_7559),
.Y(n_7734)
);

BUFx3_ASAP7_75t_L g7735 ( 
.A(n_7613),
.Y(n_7735)
);

OR2x2_ASAP7_75t_L g7736 ( 
.A(n_7586),
.B(n_7450),
.Y(n_7736)
);

NAND2xp5_ASAP7_75t_L g7737 ( 
.A(n_7618),
.B(n_7485),
.Y(n_7737)
);

HB1xp67_ASAP7_75t_L g7738 ( 
.A(n_7621),
.Y(n_7738)
);

BUFx3_ASAP7_75t_L g7739 ( 
.A(n_7552),
.Y(n_7739)
);

OR2x2_ASAP7_75t_L g7740 ( 
.A(n_7543),
.B(n_7485),
.Y(n_7740)
);

NAND2xp5_ASAP7_75t_L g7741 ( 
.A(n_7546),
.B(n_7485),
.Y(n_7741)
);

INVx2_ASAP7_75t_L g7742 ( 
.A(n_7582),
.Y(n_7742)
);

INVx2_ASAP7_75t_L g7743 ( 
.A(n_7585),
.Y(n_7743)
);

AND2x2_ASAP7_75t_L g7744 ( 
.A(n_7614),
.B(n_7490),
.Y(n_7744)
);

AND2x2_ASAP7_75t_L g7745 ( 
.A(n_7516),
.B(n_7485),
.Y(n_7745)
);

AND2x4_ASAP7_75t_L g7746 ( 
.A(n_7527),
.B(n_426),
.Y(n_7746)
);

INVx1_ASAP7_75t_SL g7747 ( 
.A(n_7520),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_7565),
.Y(n_7748)
);

AND2x2_ASAP7_75t_L g7749 ( 
.A(n_7604),
.B(n_7099),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7588),
.Y(n_7750)
);

INVx2_ASAP7_75t_L g7751 ( 
.A(n_7591),
.Y(n_7751)
);

HB1xp67_ASAP7_75t_L g7752 ( 
.A(n_7572),
.Y(n_7752)
);

AOI211xp5_ASAP7_75t_SL g7753 ( 
.A1(n_7550),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_7753)
);

AND2x2_ASAP7_75t_L g7754 ( 
.A(n_7573),
.B(n_429),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7528),
.Y(n_7755)
);

INVx2_ASAP7_75t_L g7756 ( 
.A(n_7580),
.Y(n_7756)
);

OR2x2_ASAP7_75t_L g7757 ( 
.A(n_7509),
.B(n_430),
.Y(n_7757)
);

INVxp67_ASAP7_75t_SL g7758 ( 
.A(n_7600),
.Y(n_7758)
);

INVx2_ASAP7_75t_L g7759 ( 
.A(n_7632),
.Y(n_7759)
);

AND2x4_ASAP7_75t_L g7760 ( 
.A(n_7681),
.B(n_7523),
.Y(n_7760)
);

HB1xp67_ASAP7_75t_L g7761 ( 
.A(n_7655),
.Y(n_7761)
);

HB1xp67_ASAP7_75t_L g7762 ( 
.A(n_7693),
.Y(n_7762)
);

INVx3_ASAP7_75t_L g7763 ( 
.A(n_7727),
.Y(n_7763)
);

OR2x2_ASAP7_75t_L g7764 ( 
.A(n_7710),
.B(n_7509),
.Y(n_7764)
);

AND2x2_ASAP7_75t_L g7765 ( 
.A(n_7666),
.B(n_7634),
.Y(n_7765)
);

NAND2xp5_ASAP7_75t_L g7766 ( 
.A(n_7753),
.B(n_7546),
.Y(n_7766)
);

HB1xp67_ASAP7_75t_L g7767 ( 
.A(n_7714),
.Y(n_7767)
);

HB1xp67_ASAP7_75t_L g7768 ( 
.A(n_7674),
.Y(n_7768)
);

INVx2_ASAP7_75t_L g7769 ( 
.A(n_7727),
.Y(n_7769)
);

INVx2_ASAP7_75t_L g7770 ( 
.A(n_7650),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7645),
.Y(n_7771)
);

OR2x2_ASAP7_75t_L g7772 ( 
.A(n_7710),
.B(n_7581),
.Y(n_7772)
);

INVx2_ASAP7_75t_L g7773 ( 
.A(n_7650),
.Y(n_7773)
);

NAND2xp5_ASAP7_75t_L g7774 ( 
.A(n_7753),
.B(n_7562),
.Y(n_7774)
);

NOR2xp33_ASAP7_75t_L g7775 ( 
.A(n_7747),
.B(n_7589),
.Y(n_7775)
);

AND2x2_ASAP7_75t_L g7776 ( 
.A(n_7695),
.B(n_7554),
.Y(n_7776)
);

AND2x2_ASAP7_75t_L g7777 ( 
.A(n_7643),
.B(n_7551),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7738),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7722),
.Y(n_7779)
);

AND2x2_ASAP7_75t_L g7780 ( 
.A(n_7729),
.B(n_7563),
.Y(n_7780)
);

AOI222xp33_ASAP7_75t_L g7781 ( 
.A1(n_7723),
.A2(n_7562),
.B1(n_7547),
.B2(n_7581),
.C1(n_7598),
.C2(n_7567),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7718),
.Y(n_7782)
);

AO21x2_ASAP7_75t_L g7783 ( 
.A1(n_7741),
.A2(n_7598),
.B(n_7600),
.Y(n_7783)
);

AOI31xp33_ASAP7_75t_L g7784 ( 
.A1(n_7696),
.A2(n_7567),
.A3(n_7547),
.B(n_7592),
.Y(n_7784)
);

INVx3_ASAP7_75t_L g7785 ( 
.A(n_7691),
.Y(n_7785)
);

AOI22xp33_ASAP7_75t_L g7786 ( 
.A1(n_7654),
.A2(n_7583),
.B1(n_7652),
.B2(n_7672),
.Y(n_7786)
);

INVx2_ASAP7_75t_L g7787 ( 
.A(n_7691),
.Y(n_7787)
);

AND2x2_ASAP7_75t_L g7788 ( 
.A(n_7744),
.B(n_7584),
.Y(n_7788)
);

AND2x2_ASAP7_75t_L g7789 ( 
.A(n_7692),
.B(n_7705),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_7718),
.Y(n_7790)
);

NAND2xp5_ASAP7_75t_L g7791 ( 
.A(n_7670),
.B(n_7637),
.Y(n_7791)
);

AND2x2_ASAP7_75t_L g7792 ( 
.A(n_7641),
.B(n_7566),
.Y(n_7792)
);

HB1xp67_ASAP7_75t_L g7793 ( 
.A(n_7730),
.Y(n_7793)
);

AND2x2_ASAP7_75t_L g7794 ( 
.A(n_7685),
.B(n_7619),
.Y(n_7794)
);

BUFx2_ASAP7_75t_L g7795 ( 
.A(n_7699),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7646),
.Y(n_7796)
);

AND2x2_ASAP7_75t_L g7797 ( 
.A(n_7644),
.B(n_7630),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_7651),
.Y(n_7798)
);

AND2x4_ASAP7_75t_L g7799 ( 
.A(n_7730),
.B(n_7701),
.Y(n_7799)
);

INVxp67_ASAP7_75t_L g7800 ( 
.A(n_7648),
.Y(n_7800)
);

INVx2_ASAP7_75t_L g7801 ( 
.A(n_7730),
.Y(n_7801)
);

OR2x2_ASAP7_75t_L g7802 ( 
.A(n_7747),
.B(n_7569),
.Y(n_7802)
);

INVx2_ASAP7_75t_L g7803 ( 
.A(n_7642),
.Y(n_7803)
);

AND2x2_ASAP7_75t_L g7804 ( 
.A(n_7689),
.B(n_7717),
.Y(n_7804)
);

BUFx8_ASAP7_75t_L g7805 ( 
.A(n_7656),
.Y(n_7805)
);

OAI22xp33_ASAP7_75t_L g7806 ( 
.A1(n_7652),
.A2(n_7622),
.B1(n_7594),
.B2(n_7601),
.Y(n_7806)
);

AND2x2_ASAP7_75t_L g7807 ( 
.A(n_7698),
.B(n_7623),
.Y(n_7807)
);

NAND3xp33_ASAP7_75t_L g7808 ( 
.A(n_7741),
.B(n_7599),
.C(n_7626),
.Y(n_7808)
);

INVx1_ASAP7_75t_L g7809 ( 
.A(n_7668),
.Y(n_7809)
);

AND2x2_ASAP7_75t_L g7810 ( 
.A(n_7690),
.B(n_7663),
.Y(n_7810)
);

AND2x2_ASAP7_75t_L g7811 ( 
.A(n_7671),
.B(n_7574),
.Y(n_7811)
);

OA21x2_ASAP7_75t_L g7812 ( 
.A1(n_7661),
.A2(n_7599),
.B(n_7629),
.Y(n_7812)
);

INVx1_ASAP7_75t_L g7813 ( 
.A(n_7678),
.Y(n_7813)
);

AND2x2_ASAP7_75t_L g7814 ( 
.A(n_7669),
.B(n_7576),
.Y(n_7814)
);

NOR2xp33_ASAP7_75t_L g7815 ( 
.A(n_7687),
.B(n_7622),
.Y(n_7815)
);

OAI22xp5_ASAP7_75t_SL g7816 ( 
.A1(n_7654),
.A2(n_7570),
.B1(n_7640),
.B2(n_7633),
.Y(n_7816)
);

INVx1_ASAP7_75t_L g7817 ( 
.A(n_7678),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7658),
.Y(n_7818)
);

INVx5_ASAP7_75t_L g7819 ( 
.A(n_7746),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_7752),
.Y(n_7820)
);

AND2x2_ASAP7_75t_L g7821 ( 
.A(n_7721),
.B(n_7724),
.Y(n_7821)
);

INVx5_ASAP7_75t_SL g7822 ( 
.A(n_7746),
.Y(n_7822)
);

HB1xp67_ASAP7_75t_L g7823 ( 
.A(n_7659),
.Y(n_7823)
);

AND2x4_ASAP7_75t_L g7824 ( 
.A(n_7659),
.B(n_7617),
.Y(n_7824)
);

INVx1_ASAP7_75t_L g7825 ( 
.A(n_7679),
.Y(n_7825)
);

NOR2xp33_ASAP7_75t_R g7826 ( 
.A(n_7680),
.B(n_7627),
.Y(n_7826)
);

AND2x2_ASAP7_75t_L g7827 ( 
.A(n_7756),
.B(n_7639),
.Y(n_7827)
);

INVx2_ASAP7_75t_L g7828 ( 
.A(n_7739),
.Y(n_7828)
);

INVx2_ASAP7_75t_SL g7829 ( 
.A(n_7688),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7682),
.Y(n_7830)
);

BUFx3_ASAP7_75t_L g7831 ( 
.A(n_7735),
.Y(n_7831)
);

NAND2xp5_ASAP7_75t_L g7832 ( 
.A(n_7677),
.B(n_7615),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7737),
.Y(n_7833)
);

AOI22xp5_ASAP7_75t_L g7834 ( 
.A1(n_7672),
.A2(n_7594),
.B1(n_7601),
.B2(n_7617),
.Y(n_7834)
);

AO21x2_ASAP7_75t_L g7835 ( 
.A1(n_7737),
.A2(n_7649),
.B(n_7757),
.Y(n_7835)
);

NAND2xp5_ASAP7_75t_SL g7836 ( 
.A(n_7649),
.B(n_7615),
.Y(n_7836)
);

OAI21xp5_ASAP7_75t_L g7837 ( 
.A1(n_7676),
.A2(n_7631),
.B(n_7624),
.Y(n_7837)
);

INVx2_ASAP7_75t_SL g7838 ( 
.A(n_7688),
.Y(n_7838)
);

OAI22xp5_ASAP7_75t_L g7839 ( 
.A1(n_7653),
.A2(n_7638),
.B1(n_434),
.B2(n_432),
.Y(n_7839)
);

AND2x4_ASAP7_75t_L g7840 ( 
.A(n_7684),
.B(n_433),
.Y(n_7840)
);

AND2x2_ASAP7_75t_L g7841 ( 
.A(n_7708),
.B(n_433),
.Y(n_7841)
);

NOR3xp33_ASAP7_75t_L g7842 ( 
.A(n_7657),
.B(n_7676),
.C(n_7758),
.Y(n_7842)
);

INVx2_ASAP7_75t_L g7843 ( 
.A(n_7733),
.Y(n_7843)
);

OR2x2_ASAP7_75t_L g7844 ( 
.A(n_7657),
.B(n_7675),
.Y(n_7844)
);

INVx1_ASAP7_75t_L g7845 ( 
.A(n_7716),
.Y(n_7845)
);

AND2x2_ASAP7_75t_L g7846 ( 
.A(n_7713),
.B(n_434),
.Y(n_7846)
);

AND2x2_ASAP7_75t_L g7847 ( 
.A(n_7711),
.B(n_435),
.Y(n_7847)
);

OR2x2_ASAP7_75t_L g7848 ( 
.A(n_7823),
.B(n_7647),
.Y(n_7848)
);

NAND2xp5_ASAP7_75t_L g7849 ( 
.A(n_7822),
.B(n_7700),
.Y(n_7849)
);

AND2x4_ASAP7_75t_L g7850 ( 
.A(n_7799),
.B(n_7700),
.Y(n_7850)
);

AND2x2_ASAP7_75t_L g7851 ( 
.A(n_7804),
.B(n_7712),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7783),
.Y(n_7852)
);

AND2x4_ASAP7_75t_L g7853 ( 
.A(n_7799),
.B(n_7706),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_L g7854 ( 
.A(n_7822),
.B(n_7706),
.Y(n_7854)
);

OR2x2_ASAP7_75t_L g7855 ( 
.A(n_7764),
.B(n_7822),
.Y(n_7855)
);

NOR2xp67_ASAP7_75t_L g7856 ( 
.A(n_7819),
.B(n_7829),
.Y(n_7856)
);

INVx1_ASAP7_75t_L g7857 ( 
.A(n_7793),
.Y(n_7857)
);

AND2x2_ASAP7_75t_L g7858 ( 
.A(n_7776),
.B(n_7707),
.Y(n_7858)
);

AND2x2_ASAP7_75t_L g7859 ( 
.A(n_7789),
.B(n_7709),
.Y(n_7859)
);

AND2x4_ASAP7_75t_L g7860 ( 
.A(n_7824),
.B(n_7819),
.Y(n_7860)
);

OR2x2_ASAP7_75t_L g7861 ( 
.A(n_7772),
.B(n_7647),
.Y(n_7861)
);

AND2x2_ASAP7_75t_L g7862 ( 
.A(n_7780),
.B(n_7807),
.Y(n_7862)
);

OR2x2_ASAP7_75t_L g7863 ( 
.A(n_7768),
.B(n_7673),
.Y(n_7863)
);

AND2x2_ASAP7_75t_L g7864 ( 
.A(n_7788),
.B(n_7694),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_7767),
.Y(n_7865)
);

NAND2xp5_ASAP7_75t_L g7866 ( 
.A(n_7770),
.B(n_7773),
.Y(n_7866)
);

AND2x2_ASAP7_75t_L g7867 ( 
.A(n_7794),
.B(n_7715),
.Y(n_7867)
);

NAND2x1_ASAP7_75t_SL g7868 ( 
.A(n_7761),
.B(n_7745),
.Y(n_7868)
);

AND2x2_ASAP7_75t_L g7869 ( 
.A(n_7797),
.B(n_7715),
.Y(n_7869)
);

NAND2xp5_ASAP7_75t_L g7870 ( 
.A(n_7824),
.B(n_7754),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7767),
.Y(n_7871)
);

INVx2_ASAP7_75t_L g7872 ( 
.A(n_7819),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_7762),
.Y(n_7873)
);

NAND2x1p5_ASAP7_75t_L g7874 ( 
.A(n_7831),
.B(n_7664),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7795),
.Y(n_7875)
);

INVx1_ASAP7_75t_L g7876 ( 
.A(n_7838),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_7760),
.Y(n_7877)
);

OR2x2_ASAP7_75t_L g7878 ( 
.A(n_7774),
.B(n_7791),
.Y(n_7878)
);

INVx2_ASAP7_75t_L g7879 ( 
.A(n_7785),
.Y(n_7879)
);

NAND2xp5_ASAP7_75t_L g7880 ( 
.A(n_7805),
.B(n_7750),
.Y(n_7880)
);

NAND2xp5_ASAP7_75t_L g7881 ( 
.A(n_7805),
.B(n_7660),
.Y(n_7881)
);

NAND2xp5_ASAP7_75t_SL g7882 ( 
.A(n_7784),
.B(n_7683),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_7760),
.Y(n_7883)
);

INVx2_ASAP7_75t_L g7884 ( 
.A(n_7785),
.Y(n_7884)
);

AND2x4_ASAP7_75t_L g7885 ( 
.A(n_7763),
.B(n_7742),
.Y(n_7885)
);

INVx1_ASAP7_75t_L g7886 ( 
.A(n_7783),
.Y(n_7886)
);

OR2x2_ASAP7_75t_L g7887 ( 
.A(n_7774),
.B(n_7683),
.Y(n_7887)
);

OR2x2_ASAP7_75t_L g7888 ( 
.A(n_7791),
.B(n_7704),
.Y(n_7888)
);

OAI21xp5_ASAP7_75t_L g7889 ( 
.A1(n_7784),
.A2(n_7725),
.B(n_7720),
.Y(n_7889)
);

AND2x2_ASAP7_75t_L g7890 ( 
.A(n_7765),
.B(n_7777),
.Y(n_7890)
);

AND2x2_ASAP7_75t_L g7891 ( 
.A(n_7810),
.B(n_7743),
.Y(n_7891)
);

NAND2xp5_ASAP7_75t_L g7892 ( 
.A(n_7763),
.B(n_7781),
.Y(n_7892)
);

INVx2_ASAP7_75t_L g7893 ( 
.A(n_7801),
.Y(n_7893)
);

HB1xp67_ASAP7_75t_L g7894 ( 
.A(n_7835),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_L g7895 ( 
.A(n_7781),
.B(n_7662),
.Y(n_7895)
);

INVx1_ASAP7_75t_L g7896 ( 
.A(n_7792),
.Y(n_7896)
);

OR2x2_ASAP7_75t_L g7897 ( 
.A(n_7766),
.B(n_7704),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_7771),
.Y(n_7898)
);

NAND2xp5_ASAP7_75t_L g7899 ( 
.A(n_7775),
.B(n_7665),
.Y(n_7899)
);

INVx1_ASAP7_75t_L g7900 ( 
.A(n_7832),
.Y(n_7900)
);

AND2x2_ASAP7_75t_L g7901 ( 
.A(n_7821),
.B(n_7751),
.Y(n_7901)
);

AND2x2_ASAP7_75t_L g7902 ( 
.A(n_7769),
.B(n_7828),
.Y(n_7902)
);

INVx1_ASAP7_75t_SL g7903 ( 
.A(n_7844),
.Y(n_7903)
);

INVx2_ASAP7_75t_L g7904 ( 
.A(n_7787),
.Y(n_7904)
);

INVx1_ASAP7_75t_L g7905 ( 
.A(n_7812),
.Y(n_7905)
);

AND2x2_ASAP7_75t_L g7906 ( 
.A(n_7814),
.B(n_7667),
.Y(n_7906)
);

NAND2x1p5_ASAP7_75t_L g7907 ( 
.A(n_7782),
.B(n_7759),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7812),
.Y(n_7908)
);

AND2x2_ASAP7_75t_L g7909 ( 
.A(n_7790),
.B(n_7702),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7835),
.Y(n_7910)
);

NAND2xp5_ASAP7_75t_L g7911 ( 
.A(n_7800),
.B(n_7686),
.Y(n_7911)
);

AND2x2_ASAP7_75t_L g7912 ( 
.A(n_7845),
.B(n_7736),
.Y(n_7912)
);

INVx1_ASAP7_75t_L g7913 ( 
.A(n_7808),
.Y(n_7913)
);

INVx1_ASAP7_75t_L g7914 ( 
.A(n_7808),
.Y(n_7914)
);

INVx1_ASAP7_75t_L g7915 ( 
.A(n_7802),
.Y(n_7915)
);

NAND2xp5_ASAP7_75t_L g7916 ( 
.A(n_7800),
.B(n_7697),
.Y(n_7916)
);

NAND2xp5_ASAP7_75t_L g7917 ( 
.A(n_7803),
.B(n_7786),
.Y(n_7917)
);

OR2x2_ASAP7_75t_L g7918 ( 
.A(n_7766),
.B(n_7720),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7811),
.Y(n_7919)
);

NOR2xp33_ASAP7_75t_L g7920 ( 
.A(n_7836),
.B(n_7832),
.Y(n_7920)
);

OR2x2_ASAP7_75t_L g7921 ( 
.A(n_7778),
.B(n_7725),
.Y(n_7921)
);

AND2x2_ASAP7_75t_L g7922 ( 
.A(n_7827),
.B(n_7755),
.Y(n_7922)
);

AND2x2_ASAP7_75t_L g7923 ( 
.A(n_7796),
.B(n_7843),
.Y(n_7923)
);

NAND2xp5_ASAP7_75t_L g7924 ( 
.A(n_7820),
.B(n_7740),
.Y(n_7924)
);

AND2x2_ASAP7_75t_L g7925 ( 
.A(n_7862),
.B(n_7779),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_7894),
.Y(n_7926)
);

AND2x2_ASAP7_75t_L g7927 ( 
.A(n_7869),
.B(n_7809),
.Y(n_7927)
);

INVx2_ASAP7_75t_L g7928 ( 
.A(n_7860),
.Y(n_7928)
);

INVx1_ASAP7_75t_L g7929 ( 
.A(n_7852),
.Y(n_7929)
);

AND2x2_ASAP7_75t_L g7930 ( 
.A(n_7867),
.B(n_7846),
.Y(n_7930)
);

AND2x2_ASAP7_75t_L g7931 ( 
.A(n_7864),
.B(n_7815),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7860),
.Y(n_7932)
);

INVx1_ASAP7_75t_L g7933 ( 
.A(n_7856),
.Y(n_7933)
);

HB1xp67_ASAP7_75t_L g7934 ( 
.A(n_7905),
.Y(n_7934)
);

OR2x6_ASAP7_75t_L g7935 ( 
.A(n_7849),
.B(n_7854),
.Y(n_7935)
);

NOR2xp33_ASAP7_75t_L g7936 ( 
.A(n_7861),
.B(n_7818),
.Y(n_7936)
);

INVx1_ASAP7_75t_L g7937 ( 
.A(n_7848),
.Y(n_7937)
);

BUFx3_ASAP7_75t_L g7938 ( 
.A(n_7850),
.Y(n_7938)
);

INVx2_ASAP7_75t_L g7939 ( 
.A(n_7850),
.Y(n_7939)
);

INVx1_ASAP7_75t_L g7940 ( 
.A(n_7852),
.Y(n_7940)
);

INVx2_ASAP7_75t_SL g7941 ( 
.A(n_7853),
.Y(n_7941)
);

NAND2xp5_ASAP7_75t_L g7942 ( 
.A(n_7853),
.B(n_7842),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7886),
.Y(n_7943)
);

NAND2x1_ASAP7_75t_L g7944 ( 
.A(n_7872),
.B(n_7840),
.Y(n_7944)
);

INVx2_ASAP7_75t_L g7945 ( 
.A(n_7855),
.Y(n_7945)
);

NAND2x1_ASAP7_75t_L g7946 ( 
.A(n_7877),
.B(n_7883),
.Y(n_7946)
);

NAND2xp5_ASAP7_75t_L g7947 ( 
.A(n_7859),
.B(n_7842),
.Y(n_7947)
);

INVx1_ASAP7_75t_L g7948 ( 
.A(n_7886),
.Y(n_7948)
);

HB1xp67_ASAP7_75t_L g7949 ( 
.A(n_7905),
.Y(n_7949)
);

AND2x2_ASAP7_75t_L g7950 ( 
.A(n_7890),
.B(n_7847),
.Y(n_7950)
);

OR2x2_ASAP7_75t_L g7951 ( 
.A(n_7863),
.B(n_7813),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7910),
.Y(n_7952)
);

INVx1_ASAP7_75t_L g7953 ( 
.A(n_7910),
.Y(n_7953)
);

AND2x2_ASAP7_75t_L g7954 ( 
.A(n_7858),
.B(n_7841),
.Y(n_7954)
);

INVx2_ASAP7_75t_L g7955 ( 
.A(n_7868),
.Y(n_7955)
);

INVx4_ASAP7_75t_L g7956 ( 
.A(n_7885),
.Y(n_7956)
);

INVx1_ASAP7_75t_L g7957 ( 
.A(n_7866),
.Y(n_7957)
);

AND2x2_ASAP7_75t_L g7958 ( 
.A(n_7851),
.B(n_7798),
.Y(n_7958)
);

NOR2x1_ASAP7_75t_L g7959 ( 
.A(n_7908),
.B(n_7840),
.Y(n_7959)
);

INVx1_ASAP7_75t_L g7960 ( 
.A(n_7870),
.Y(n_7960)
);

INVx1_ASAP7_75t_L g7961 ( 
.A(n_7865),
.Y(n_7961)
);

AND2x2_ASAP7_75t_L g7962 ( 
.A(n_7919),
.B(n_7826),
.Y(n_7962)
);

NAND2xp5_ASAP7_75t_L g7963 ( 
.A(n_7885),
.B(n_7834),
.Y(n_7963)
);

INVx1_ASAP7_75t_SL g7964 ( 
.A(n_7903),
.Y(n_7964)
);

NAND2x1p5_ASAP7_75t_L g7965 ( 
.A(n_7875),
.B(n_7817),
.Y(n_7965)
);

OR2x2_ASAP7_75t_L g7966 ( 
.A(n_7878),
.B(n_7825),
.Y(n_7966)
);

OR2x2_ASAP7_75t_L g7967 ( 
.A(n_7892),
.B(n_7830),
.Y(n_7967)
);

INVx1_ASAP7_75t_L g7968 ( 
.A(n_7871),
.Y(n_7968)
);

NAND2xp5_ASAP7_75t_L g7969 ( 
.A(n_7879),
.B(n_7834),
.Y(n_7969)
);

INVx1_ASAP7_75t_L g7970 ( 
.A(n_7908),
.Y(n_7970)
);

OR2x6_ASAP7_75t_L g7971 ( 
.A(n_7907),
.B(n_7816),
.Y(n_7971)
);

INVx2_ASAP7_75t_L g7972 ( 
.A(n_7884),
.Y(n_7972)
);

INVxp67_ASAP7_75t_L g7973 ( 
.A(n_7920),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_7906),
.Y(n_7974)
);

OR2x2_ASAP7_75t_L g7975 ( 
.A(n_7887),
.B(n_7839),
.Y(n_7975)
);

INVx1_ASAP7_75t_L g7976 ( 
.A(n_7857),
.Y(n_7976)
);

INVx1_ASAP7_75t_L g7977 ( 
.A(n_7876),
.Y(n_7977)
);

INVx1_ASAP7_75t_L g7978 ( 
.A(n_7881),
.Y(n_7978)
);

INVx3_ASAP7_75t_R g7979 ( 
.A(n_7921),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_7909),
.Y(n_7980)
);

BUFx2_ASAP7_75t_L g7981 ( 
.A(n_7913),
.Y(n_7981)
);

AND2x2_ASAP7_75t_L g7982 ( 
.A(n_7891),
.B(n_7837),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_L g7983 ( 
.A(n_7913),
.B(n_7806),
.Y(n_7983)
);

AO221x1_ASAP7_75t_L g7984 ( 
.A1(n_7914),
.A2(n_7839),
.B1(n_7816),
.B2(n_7726),
.C(n_7728),
.Y(n_7984)
);

INVx1_ASAP7_75t_L g7985 ( 
.A(n_7901),
.Y(n_7985)
);

AO22x1_ASAP7_75t_L g7986 ( 
.A1(n_7914),
.A2(n_7889),
.B1(n_7895),
.B2(n_7915),
.Y(n_7986)
);

NAND2xp5_ASAP7_75t_L g7987 ( 
.A(n_7915),
.B(n_7703),
.Y(n_7987)
);

OR2x2_ASAP7_75t_L g7988 ( 
.A(n_7897),
.B(n_7918),
.Y(n_7988)
);

INVx1_ASAP7_75t_L g7989 ( 
.A(n_7934),
.Y(n_7989)
);

NOR2x1p5_ASAP7_75t_L g7990 ( 
.A(n_7946),
.B(n_7899),
.Y(n_7990)
);

OAI21xp33_ASAP7_75t_L g7991 ( 
.A1(n_7964),
.A2(n_7917),
.B(n_7880),
.Y(n_7991)
);

NAND2xp33_ASAP7_75t_R g7992 ( 
.A(n_7971),
.B(n_7912),
.Y(n_7992)
);

INVx1_ASAP7_75t_L g7993 ( 
.A(n_7949),
.Y(n_7993)
);

OR2x2_ASAP7_75t_L g7994 ( 
.A(n_7941),
.B(n_7882),
.Y(n_7994)
);

INVx1_ASAP7_75t_L g7995 ( 
.A(n_7959),
.Y(n_7995)
);

NAND2xp5_ASAP7_75t_SL g7996 ( 
.A(n_7956),
.B(n_7873),
.Y(n_7996)
);

INVx1_ASAP7_75t_SL g7997 ( 
.A(n_7938),
.Y(n_7997)
);

OR2x2_ASAP7_75t_L g7998 ( 
.A(n_7956),
.B(n_7888),
.Y(n_7998)
);

INVx1_ASAP7_75t_L g7999 ( 
.A(n_7970),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_7970),
.Y(n_8000)
);

INVx1_ASAP7_75t_L g8001 ( 
.A(n_7932),
.Y(n_8001)
);

INVx1_ASAP7_75t_L g8002 ( 
.A(n_7928),
.Y(n_8002)
);

INVx1_ASAP7_75t_L g8003 ( 
.A(n_7925),
.Y(n_8003)
);

INVxp67_ASAP7_75t_L g8004 ( 
.A(n_7971),
.Y(n_8004)
);

AND2x2_ASAP7_75t_L g8005 ( 
.A(n_7939),
.B(n_7902),
.Y(n_8005)
);

NOR2x1_ASAP7_75t_L g8006 ( 
.A(n_7981),
.B(n_7924),
.Y(n_8006)
);

AND2x2_ASAP7_75t_L g8007 ( 
.A(n_7930),
.B(n_7922),
.Y(n_8007)
);

NAND4xp75_ASAP7_75t_L g8008 ( 
.A(n_7931),
.B(n_7923),
.C(n_7900),
.D(n_7898),
.Y(n_8008)
);

AND2x2_ASAP7_75t_L g8009 ( 
.A(n_7927),
.B(n_7874),
.Y(n_8009)
);

OR2x2_ASAP7_75t_L g8010 ( 
.A(n_7944),
.B(n_7893),
.Y(n_8010)
);

INVx1_ASAP7_75t_L g8011 ( 
.A(n_7986),
.Y(n_8011)
);

NAND2xp5_ASAP7_75t_SL g8012 ( 
.A(n_7955),
.B(n_7896),
.Y(n_8012)
);

INVx2_ASAP7_75t_L g8013 ( 
.A(n_7935),
.Y(n_8013)
);

HB1xp67_ASAP7_75t_L g8014 ( 
.A(n_7979),
.Y(n_8014)
);

INVx1_ASAP7_75t_L g8015 ( 
.A(n_7950),
.Y(n_8015)
);

OR2x2_ASAP7_75t_L g8016 ( 
.A(n_7963),
.B(n_7942),
.Y(n_8016)
);

INVx1_ASAP7_75t_L g8017 ( 
.A(n_7954),
.Y(n_8017)
);

AOI221xp5_ASAP7_75t_L g8018 ( 
.A1(n_7986),
.A2(n_7837),
.B1(n_7904),
.B2(n_7916),
.C(n_7911),
.Y(n_8018)
);

OR2x6_ASAP7_75t_L g8019 ( 
.A(n_7965),
.B(n_7734),
.Y(n_8019)
);

INVx1_ASAP7_75t_L g8020 ( 
.A(n_7966),
.Y(n_8020)
);

INVx1_ASAP7_75t_SL g8021 ( 
.A(n_7951),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7958),
.Y(n_8022)
);

NAND2xp5_ASAP7_75t_L g8023 ( 
.A(n_7933),
.B(n_7719),
.Y(n_8023)
);

OR2x2_ASAP7_75t_L g8024 ( 
.A(n_7975),
.B(n_7748),
.Y(n_8024)
);

NAND2xp5_ASAP7_75t_L g8025 ( 
.A(n_7962),
.B(n_7731),
.Y(n_8025)
);

INVx2_ASAP7_75t_L g8026 ( 
.A(n_7935),
.Y(n_8026)
);

BUFx12f_ASAP7_75t_L g8027 ( 
.A(n_7988),
.Y(n_8027)
);

OR2x2_ASAP7_75t_L g8028 ( 
.A(n_7947),
.B(n_7732),
.Y(n_8028)
);

OR2x2_ASAP7_75t_L g8029 ( 
.A(n_7969),
.B(n_7974),
.Y(n_8029)
);

AND2x4_ASAP7_75t_L g8030 ( 
.A(n_7937),
.B(n_7833),
.Y(n_8030)
);

NAND2xp5_ASAP7_75t_L g8031 ( 
.A(n_7982),
.B(n_7980),
.Y(n_8031)
);

NAND2xp5_ASAP7_75t_L g8032 ( 
.A(n_7984),
.B(n_7749),
.Y(n_8032)
);

INVx1_ASAP7_75t_L g8033 ( 
.A(n_7945),
.Y(n_8033)
);

OR2x2_ASAP7_75t_L g8034 ( 
.A(n_7985),
.B(n_435),
.Y(n_8034)
);

INVx2_ASAP7_75t_SL g8035 ( 
.A(n_7972),
.Y(n_8035)
);

INVx2_ASAP7_75t_L g8036 ( 
.A(n_7977),
.Y(n_8036)
);

OR2x2_ASAP7_75t_L g8037 ( 
.A(n_7983),
.B(n_436),
.Y(n_8037)
);

CKINVDCx14_ASAP7_75t_R g8038 ( 
.A(n_8009),
.Y(n_8038)
);

AOI32xp33_ASAP7_75t_L g8039 ( 
.A1(n_8011),
.A2(n_7978),
.A3(n_7976),
.B1(n_7936),
.B2(n_7957),
.Y(n_8039)
);

INVx1_ASAP7_75t_L g8040 ( 
.A(n_8010),
.Y(n_8040)
);

AND2x2_ASAP7_75t_L g8041 ( 
.A(n_8007),
.B(n_7973),
.Y(n_8041)
);

NOR2x1_ASAP7_75t_L g8042 ( 
.A(n_8019),
.B(n_7987),
.Y(n_8042)
);

INVx1_ASAP7_75t_L g8043 ( 
.A(n_8019),
.Y(n_8043)
);

AOI21xp5_ASAP7_75t_L g8044 ( 
.A1(n_7996),
.A2(n_7926),
.B(n_7960),
.Y(n_8044)
);

HB1xp67_ASAP7_75t_L g8045 ( 
.A(n_7992),
.Y(n_8045)
);

INVx2_ASAP7_75t_SL g8046 ( 
.A(n_7998),
.Y(n_8046)
);

NAND2x2_ASAP7_75t_L g8047 ( 
.A(n_7990),
.B(n_7967),
.Y(n_8047)
);

INVx1_ASAP7_75t_SL g8048 ( 
.A(n_8027),
.Y(n_8048)
);

NAND2xp5_ASAP7_75t_L g8049 ( 
.A(n_7997),
.B(n_7961),
.Y(n_8049)
);

INVx1_ASAP7_75t_SL g8050 ( 
.A(n_7994),
.Y(n_8050)
);

INVx1_ASAP7_75t_L g8051 ( 
.A(n_8005),
.Y(n_8051)
);

INVx1_ASAP7_75t_L g8052 ( 
.A(n_8014),
.Y(n_8052)
);

OAI31xp33_ASAP7_75t_L g8053 ( 
.A1(n_8011),
.A2(n_8021),
.A3(n_7995),
.B(n_7993),
.Y(n_8053)
);

NOR2x1_ASAP7_75t_L g8054 ( 
.A(n_8006),
.B(n_7926),
.Y(n_8054)
);

OR2x2_ASAP7_75t_L g8055 ( 
.A(n_8002),
.B(n_7968),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_7989),
.Y(n_8056)
);

INVx1_ASAP7_75t_L g8057 ( 
.A(n_7989),
.Y(n_8057)
);

AOI33xp33_ASAP7_75t_L g8058 ( 
.A1(n_8001),
.A2(n_7953),
.A3(n_7952),
.B1(n_7943),
.B2(n_7940),
.B3(n_7948),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_8013),
.Y(n_8059)
);

OAI21xp5_ASAP7_75t_L g8060 ( 
.A1(n_8004),
.A2(n_7948),
.B(n_7929),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_8015),
.Y(n_8061)
);

INVx1_ASAP7_75t_L g8062 ( 
.A(n_8034),
.Y(n_8062)
);

NOR2xp33_ASAP7_75t_L g8063 ( 
.A(n_8003),
.B(n_7929),
.Y(n_8063)
);

AND2x4_ASAP7_75t_L g8064 ( 
.A(n_8030),
.B(n_437),
.Y(n_8064)
);

AND2x4_ASAP7_75t_L g8065 ( 
.A(n_8030),
.B(n_8026),
.Y(n_8065)
);

INVx1_ASAP7_75t_L g8066 ( 
.A(n_8024),
.Y(n_8066)
);

OR2x2_ASAP7_75t_L g8067 ( 
.A(n_8017),
.B(n_8031),
.Y(n_8067)
);

INVx1_ASAP7_75t_L g8068 ( 
.A(n_8016),
.Y(n_8068)
);

XNOR2x1_ASAP7_75t_L g8069 ( 
.A(n_8008),
.B(n_438),
.Y(n_8069)
);

AND2x2_ASAP7_75t_L g8070 ( 
.A(n_8022),
.B(n_438),
.Y(n_8070)
);

NAND3xp33_ASAP7_75t_L g8071 ( 
.A(n_8053),
.B(n_8018),
.C(n_8042),
.Y(n_8071)
);

NAND2x1p5_ASAP7_75t_L g8072 ( 
.A(n_8046),
.B(n_8020),
.Y(n_8072)
);

AOI21xp33_ASAP7_75t_L g8073 ( 
.A1(n_8045),
.A2(n_7991),
.B(n_8033),
.Y(n_8073)
);

AOI22xp5_ASAP7_75t_L g8074 ( 
.A1(n_8038),
.A2(n_8035),
.B1(n_8012),
.B2(n_8032),
.Y(n_8074)
);

INVx2_ASAP7_75t_SL g8075 ( 
.A(n_8065),
.Y(n_8075)
);

INVx1_ASAP7_75t_SL g8076 ( 
.A(n_8048),
.Y(n_8076)
);

AOI21xp33_ASAP7_75t_L g8077 ( 
.A1(n_8054),
.A2(n_8029),
.B(n_8028),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_8064),
.Y(n_8078)
);

INVx1_ASAP7_75t_SL g8079 ( 
.A(n_8065),
.Y(n_8079)
);

INVx2_ASAP7_75t_L g8080 ( 
.A(n_8064),
.Y(n_8080)
);

NAND2xp5_ASAP7_75t_L g8081 ( 
.A(n_8050),
.B(n_8036),
.Y(n_8081)
);

AOI21xp33_ASAP7_75t_L g8082 ( 
.A1(n_8043),
.A2(n_8025),
.B(n_8023),
.Y(n_8082)
);

AND2x2_ASAP7_75t_L g8083 ( 
.A(n_8041),
.B(n_8037),
.Y(n_8083)
);

AND2x2_ASAP7_75t_L g8084 ( 
.A(n_8051),
.B(n_7999),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_8070),
.Y(n_8085)
);

NAND2xp5_ASAP7_75t_L g8086 ( 
.A(n_8040),
.B(n_8000),
.Y(n_8086)
);

OR2x2_ASAP7_75t_L g8087 ( 
.A(n_8055),
.B(n_439),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_8069),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_8058),
.Y(n_8089)
);

INVx1_ASAP7_75t_L g8090 ( 
.A(n_8047),
.Y(n_8090)
);

INVxp67_ASAP7_75t_L g8091 ( 
.A(n_8063),
.Y(n_8091)
);

NAND2xp5_ASAP7_75t_L g8092 ( 
.A(n_8052),
.B(n_440),
.Y(n_8092)
);

OR2x2_ASAP7_75t_L g8093 ( 
.A(n_8067),
.B(n_441),
.Y(n_8093)
);

NOR3xp33_ASAP7_75t_L g8094 ( 
.A(n_8068),
.B(n_441),
.C(n_442),
.Y(n_8094)
);

INVx1_ASAP7_75t_L g8095 ( 
.A(n_8049),
.Y(n_8095)
);

AND2x2_ASAP7_75t_L g8096 ( 
.A(n_8059),
.B(n_444),
.Y(n_8096)
);

NAND2xp5_ASAP7_75t_L g8097 ( 
.A(n_8056),
.B(n_445),
.Y(n_8097)
);

AOI22xp5_ASAP7_75t_L g8098 ( 
.A1(n_8061),
.A2(n_4003),
.B1(n_3948),
.B2(n_4049),
.Y(n_8098)
);

INVx1_ASAP7_75t_L g8099 ( 
.A(n_8057),
.Y(n_8099)
);

INVx2_ASAP7_75t_L g8100 ( 
.A(n_8066),
.Y(n_8100)
);

AOI21xp5_ASAP7_75t_L g8101 ( 
.A1(n_8044),
.A2(n_446),
.B(n_447),
.Y(n_8101)
);

O2A1O1Ixp33_ASAP7_75t_L g8102 ( 
.A1(n_8060),
.A2(n_449),
.B(n_447),
.C(n_448),
.Y(n_8102)
);

AND2x2_ASAP7_75t_L g8103 ( 
.A(n_8079),
.B(n_8062),
.Y(n_8103)
);

OAI22xp5_ASAP7_75t_L g8104 ( 
.A1(n_8074),
.A2(n_8039),
.B1(n_452),
.B2(n_448),
.Y(n_8104)
);

INVx1_ASAP7_75t_L g8105 ( 
.A(n_8075),
.Y(n_8105)
);

NAND2xp33_ASAP7_75t_SL g8106 ( 
.A(n_8080),
.B(n_450),
.Y(n_8106)
);

INVxp67_ASAP7_75t_L g8107 ( 
.A(n_8096),
.Y(n_8107)
);

NAND3xp33_ASAP7_75t_L g8108 ( 
.A(n_8071),
.B(n_453),
.C(n_454),
.Y(n_8108)
);

INVx1_ASAP7_75t_L g8109 ( 
.A(n_8072),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_8087),
.Y(n_8110)
);

XNOR2xp5_ASAP7_75t_L g8111 ( 
.A(n_8076),
.B(n_453),
.Y(n_8111)
);

INVx3_ASAP7_75t_L g8112 ( 
.A(n_8078),
.Y(n_8112)
);

AOI32xp33_ASAP7_75t_L g8113 ( 
.A1(n_8089),
.A2(n_457),
.A3(n_455),
.B1(n_456),
.B2(n_458),
.Y(n_8113)
);

AOI22xp5_ASAP7_75t_L g8114 ( 
.A1(n_8090),
.A2(n_4003),
.B1(n_3948),
.B2(n_4049),
.Y(n_8114)
);

AOI22xp5_ASAP7_75t_L g8115 ( 
.A1(n_8090),
.A2(n_3948),
.B1(n_4070),
.B2(n_2278),
.Y(n_8115)
);

OAI22xp5_ASAP7_75t_L g8116 ( 
.A1(n_8091),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_8116)
);

AOI22xp5_ASAP7_75t_L g8117 ( 
.A1(n_8100),
.A2(n_4070),
.B1(n_2278),
.B2(n_2326),
.Y(n_8117)
);

OAI21xp5_ASAP7_75t_L g8118 ( 
.A1(n_8073),
.A2(n_460),
.B(n_462),
.Y(n_8118)
);

OAI22xp5_ASAP7_75t_L g8119 ( 
.A1(n_8081),
.A2(n_464),
.B1(n_460),
.B2(n_462),
.Y(n_8119)
);

AOI22xp33_ASAP7_75t_L g8120 ( 
.A1(n_8095),
.A2(n_2278),
.B1(n_2326),
.B2(n_2166),
.Y(n_8120)
);

NAND5xp2_ASAP7_75t_L g8121 ( 
.A(n_8088),
.B(n_465),
.C(n_466),
.D(n_468),
.E(n_469),
.Y(n_8121)
);

OAI22xp5_ASAP7_75t_L g8122 ( 
.A1(n_8086),
.A2(n_8092),
.B1(n_8093),
.B2(n_8085),
.Y(n_8122)
);

NAND2xp5_ASAP7_75t_SL g8123 ( 
.A(n_8077),
.B(n_465),
.Y(n_8123)
);

OAI21xp33_ASAP7_75t_SL g8124 ( 
.A1(n_8082),
.A2(n_466),
.B(n_468),
.Y(n_8124)
);

INVxp67_ASAP7_75t_SL g8125 ( 
.A(n_8102),
.Y(n_8125)
);

OR2x2_ASAP7_75t_L g8126 ( 
.A(n_8097),
.B(n_8099),
.Y(n_8126)
);

OR2x2_ASAP7_75t_L g8127 ( 
.A(n_8084),
.B(n_470),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_8083),
.Y(n_8128)
);

NAND2xp5_ASAP7_75t_L g8129 ( 
.A(n_8101),
.B(n_8094),
.Y(n_8129)
);

NOR2xp33_ASAP7_75t_L g8130 ( 
.A(n_8098),
.B(n_470),
.Y(n_8130)
);

INVx2_ASAP7_75t_L g8131 ( 
.A(n_8075),
.Y(n_8131)
);

A2O1A1Ixp33_ASAP7_75t_L g8132 ( 
.A1(n_8071),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_8132)
);

NAND2xp5_ASAP7_75t_L g8133 ( 
.A(n_8075),
.B(n_474),
.Y(n_8133)
);

OAI221xp5_ASAP7_75t_L g8134 ( 
.A1(n_8074),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.C(n_480),
.Y(n_8134)
);

OAI21xp33_ASAP7_75t_L g8135 ( 
.A1(n_8074),
.A2(n_477),
.B(n_481),
.Y(n_8135)
);

AOI21xp5_ASAP7_75t_L g8136 ( 
.A1(n_8077),
.A2(n_482),
.B(n_485),
.Y(n_8136)
);

NAND2xp5_ASAP7_75t_SL g8137 ( 
.A(n_8075),
.B(n_482),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_8075),
.Y(n_8138)
);

INVx1_ASAP7_75t_L g8139 ( 
.A(n_8111),
.Y(n_8139)
);

AOI22xp5_ASAP7_75t_L g8140 ( 
.A1(n_8109),
.A2(n_2326),
.B1(n_2166),
.B2(n_488),
.Y(n_8140)
);

AOI22xp5_ASAP7_75t_L g8141 ( 
.A1(n_8105),
.A2(n_2326),
.B1(n_2166),
.B2(n_488),
.Y(n_8141)
);

NOR2xp33_ASAP7_75t_L g8142 ( 
.A(n_8121),
.B(n_485),
.Y(n_8142)
);

OAI22xp5_ASAP7_75t_L g8143 ( 
.A1(n_8138),
.A2(n_490),
.B1(n_486),
.B2(n_489),
.Y(n_8143)
);

INVxp67_ASAP7_75t_L g8144 ( 
.A(n_8127),
.Y(n_8144)
);

NAND2xp5_ASAP7_75t_L g8145 ( 
.A(n_8112),
.B(n_486),
.Y(n_8145)
);

NOR2xp33_ASAP7_75t_L g8146 ( 
.A(n_8112),
.B(n_490),
.Y(n_8146)
);

AOI322xp5_ASAP7_75t_L g8147 ( 
.A1(n_8135),
.A2(n_492),
.A3(n_494),
.B1(n_495),
.B2(n_496),
.C1(n_497),
.C2(n_499),
.Y(n_8147)
);

INVx1_ASAP7_75t_L g8148 ( 
.A(n_8103),
.Y(n_8148)
);

OAI221xp5_ASAP7_75t_L g8149 ( 
.A1(n_8113),
.A2(n_494),
.B1(n_497),
.B2(n_500),
.C(n_501),
.Y(n_8149)
);

INVx1_ASAP7_75t_L g8150 ( 
.A(n_8133),
.Y(n_8150)
);

NAND2xp5_ASAP7_75t_L g8151 ( 
.A(n_8131),
.B(n_501),
.Y(n_8151)
);

INVx1_ASAP7_75t_L g8152 ( 
.A(n_8128),
.Y(n_8152)
);

INVx1_ASAP7_75t_SL g8153 ( 
.A(n_8106),
.Y(n_8153)
);

INVx1_ASAP7_75t_L g8154 ( 
.A(n_8137),
.Y(n_8154)
);

OAI311xp33_ASAP7_75t_L g8155 ( 
.A1(n_8108),
.A2(n_502),
.A3(n_503),
.B1(n_504),
.C1(n_507),
.Y(n_8155)
);

INVxp67_ASAP7_75t_L g8156 ( 
.A(n_8123),
.Y(n_8156)
);

NOR2xp33_ASAP7_75t_L g8157 ( 
.A(n_8134),
.B(n_503),
.Y(n_8157)
);

AOI22xp5_ASAP7_75t_L g8158 ( 
.A1(n_8104),
.A2(n_2326),
.B1(n_509),
.B2(n_504),
.Y(n_8158)
);

OAI211xp5_ASAP7_75t_L g8159 ( 
.A1(n_8124),
.A2(n_512),
.B(n_508),
.C(n_511),
.Y(n_8159)
);

AND2x4_ASAP7_75t_L g8160 ( 
.A(n_8110),
.B(n_508),
.Y(n_8160)
);

AOI22xp33_ASAP7_75t_L g8161 ( 
.A1(n_8125),
.A2(n_514),
.B1(n_511),
.B2(n_512),
.Y(n_8161)
);

OR2x2_ASAP7_75t_L g8162 ( 
.A(n_8132),
.B(n_514),
.Y(n_8162)
);

AOI222xp33_ASAP7_75t_L g8163 ( 
.A1(n_8107),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.C1(n_518),
.C2(n_519),
.Y(n_8163)
);

NAND2xp5_ASAP7_75t_L g8164 ( 
.A(n_8136),
.B(n_517),
.Y(n_8164)
);

O2A1O1Ixp33_ASAP7_75t_L g8165 ( 
.A1(n_8118),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_8165)
);

NOR2xp33_ASAP7_75t_L g8166 ( 
.A(n_8129),
.B(n_520),
.Y(n_8166)
);

OAI221xp5_ASAP7_75t_L g8167 ( 
.A1(n_8122),
.A2(n_522),
.B1(n_523),
.B2(n_524),
.C(n_526),
.Y(n_8167)
);

AND2x2_ASAP7_75t_L g8168 ( 
.A(n_8126),
.B(n_522),
.Y(n_8168)
);

NOR2xp33_ASAP7_75t_L g8169 ( 
.A(n_8119),
.B(n_526),
.Y(n_8169)
);

INVx1_ASAP7_75t_L g8170 ( 
.A(n_8116),
.Y(n_8170)
);

NAND2xp5_ASAP7_75t_L g8171 ( 
.A(n_8130),
.B(n_527),
.Y(n_8171)
);

INVx1_ASAP7_75t_L g8172 ( 
.A(n_8114),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_8117),
.Y(n_8173)
);

OAI21xp33_ASAP7_75t_L g8174 ( 
.A1(n_8115),
.A2(n_528),
.B(n_529),
.Y(n_8174)
);

AOI22xp5_ASAP7_75t_L g8175 ( 
.A1(n_8142),
.A2(n_8120),
.B1(n_530),
.B2(n_528),
.Y(n_8175)
);

AOI21xp5_ASAP7_75t_L g8176 ( 
.A1(n_8145),
.A2(n_8164),
.B(n_8148),
.Y(n_8176)
);

OAI221xp5_ASAP7_75t_L g8177 ( 
.A1(n_8149),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.C(n_532),
.Y(n_8177)
);

OAI211xp5_ASAP7_75t_L g8178 ( 
.A1(n_8159),
.A2(n_533),
.B(n_531),
.C(n_532),
.Y(n_8178)
);

NAND4xp25_ASAP7_75t_L g8179 ( 
.A(n_8152),
.B(n_536),
.C(n_533),
.D(n_534),
.Y(n_8179)
);

NOR2xp67_ASAP7_75t_L g8180 ( 
.A(n_8167),
.B(n_8146),
.Y(n_8180)
);

INVx2_ASAP7_75t_L g8181 ( 
.A(n_8160),
.Y(n_8181)
);

NAND4xp25_ASAP7_75t_L g8182 ( 
.A(n_8157),
.B(n_537),
.C(n_534),
.D(n_536),
.Y(n_8182)
);

NOR2xp33_ASAP7_75t_L g8183 ( 
.A(n_8151),
.B(n_537),
.Y(n_8183)
);

NAND3xp33_ASAP7_75t_L g8184 ( 
.A(n_8166),
.B(n_538),
.C(n_540),
.Y(n_8184)
);

AOI221xp5_ASAP7_75t_L g8185 ( 
.A1(n_8165),
.A2(n_538),
.B1(n_540),
.B2(n_541),
.C(n_542),
.Y(n_8185)
);

OAI32xp33_ASAP7_75t_L g8186 ( 
.A1(n_8153),
.A2(n_541),
.A3(n_543),
.B1(n_544),
.B2(n_545),
.Y(n_8186)
);

AOI21xp5_ASAP7_75t_L g8187 ( 
.A1(n_8144),
.A2(n_543),
.B(n_547),
.Y(n_8187)
);

NOR2x1_ASAP7_75t_L g8188 ( 
.A(n_8168),
.B(n_547),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_8160),
.Y(n_8189)
);

NOR4xp25_ASAP7_75t_L g8190 ( 
.A(n_8170),
.B(n_548),
.C(n_549),
.D(n_550),
.Y(n_8190)
);

AOI22xp33_ASAP7_75t_L g8191 ( 
.A1(n_8139),
.A2(n_548),
.B1(n_550),
.B2(n_551),
.Y(n_8191)
);

AND2x2_ASAP7_75t_L g8192 ( 
.A(n_8154),
.B(n_551),
.Y(n_8192)
);

OAI21xp5_ASAP7_75t_SL g8193 ( 
.A1(n_8156),
.A2(n_552),
.B(n_553),
.Y(n_8193)
);

O2A1O1Ixp5_ASAP7_75t_L g8194 ( 
.A1(n_8155),
.A2(n_553),
.B(n_554),
.C(n_555),
.Y(n_8194)
);

OA22x2_ASAP7_75t_L g8195 ( 
.A1(n_8158),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_8195)
);

AOI22xp5_ASAP7_75t_L g8196 ( 
.A1(n_8169),
.A2(n_557),
.B1(n_558),
.B2(n_559),
.Y(n_8196)
);

NAND4xp25_ASAP7_75t_SL g8197 ( 
.A(n_8162),
.B(n_558),
.C(n_559),
.D(n_560),
.Y(n_8197)
);

O2A1O1Ixp33_ASAP7_75t_L g8198 ( 
.A1(n_8171),
.A2(n_560),
.B(n_561),
.C(n_562),
.Y(n_8198)
);

NAND2xp5_ASAP7_75t_SL g8199 ( 
.A(n_8161),
.B(n_562),
.Y(n_8199)
);

AOI22xp5_ASAP7_75t_L g8200 ( 
.A1(n_8150),
.A2(n_564),
.B1(n_565),
.B2(n_566),
.Y(n_8200)
);

OAI21xp5_ASAP7_75t_L g8201 ( 
.A1(n_8174),
.A2(n_565),
.B(n_568),
.Y(n_8201)
);

NOR4xp25_ASAP7_75t_L g8202 ( 
.A(n_8172),
.B(n_570),
.C(n_571),
.D(n_572),
.Y(n_8202)
);

OAI22xp33_ASAP7_75t_L g8203 ( 
.A1(n_8173),
.A2(n_570),
.B1(n_571),
.B2(n_573),
.Y(n_8203)
);

AOI222xp33_ASAP7_75t_L g8204 ( 
.A1(n_8143),
.A2(n_573),
.B1(n_574),
.B2(n_576),
.C1(n_578),
.C2(n_579),
.Y(n_8204)
);

AOI211xp5_ASAP7_75t_L g8205 ( 
.A1(n_8147),
.A2(n_574),
.B(n_578),
.C(n_579),
.Y(n_8205)
);

INVx2_ASAP7_75t_L g8206 ( 
.A(n_8140),
.Y(n_8206)
);

A2O1A1Ixp33_ASAP7_75t_L g8207 ( 
.A1(n_8141),
.A2(n_580),
.B(n_581),
.C(n_582),
.Y(n_8207)
);

OAI211xp5_ASAP7_75t_L g8208 ( 
.A1(n_8163),
.A2(n_580),
.B(n_583),
.C(n_584),
.Y(n_8208)
);

NOR3xp33_ASAP7_75t_L g8209 ( 
.A(n_8189),
.B(n_585),
.C(n_586),
.Y(n_8209)
);

NAND2xp5_ASAP7_75t_L g8210 ( 
.A(n_8192),
.B(n_587),
.Y(n_8210)
);

AOI22xp5_ASAP7_75t_L g8211 ( 
.A1(n_8197),
.A2(n_587),
.B1(n_588),
.B2(n_589),
.Y(n_8211)
);

OAI222xp33_ASAP7_75t_L g8212 ( 
.A1(n_8199),
.A2(n_588),
.B1(n_590),
.B2(n_591),
.C1(n_592),
.C2(n_593),
.Y(n_8212)
);

INVx1_ASAP7_75t_L g8213 ( 
.A(n_8188),
.Y(n_8213)
);

OAI221xp5_ASAP7_75t_L g8214 ( 
.A1(n_8185),
.A2(n_591),
.B1(n_594),
.B2(n_595),
.C(n_597),
.Y(n_8214)
);

NAND4xp25_ASAP7_75t_L g8215 ( 
.A(n_8194),
.B(n_594),
.C(n_598),
.D(n_599),
.Y(n_8215)
);

OAI211xp5_ASAP7_75t_L g8216 ( 
.A1(n_8202),
.A2(n_599),
.B(n_600),
.C(n_601),
.Y(n_8216)
);

AOI21xp5_ASAP7_75t_L g8217 ( 
.A1(n_8181),
.A2(n_600),
.B(n_601),
.Y(n_8217)
);

AOI22xp5_ASAP7_75t_L g8218 ( 
.A1(n_8180),
.A2(n_602),
.B1(n_605),
.B2(n_606),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_8184),
.Y(n_8219)
);

HB1xp67_ASAP7_75t_L g8220 ( 
.A(n_8190),
.Y(n_8220)
);

OAI211xp5_ASAP7_75t_SL g8221 ( 
.A1(n_8176),
.A2(n_602),
.B(n_606),
.C(n_607),
.Y(n_8221)
);

NAND4xp75_ASAP7_75t_L g8222 ( 
.A(n_8175),
.B(n_607),
.C(n_608),
.D(n_611),
.Y(n_8222)
);

OAI21xp5_ASAP7_75t_L g8223 ( 
.A1(n_8178),
.A2(n_608),
.B(n_611),
.Y(n_8223)
);

NOR2xp67_ASAP7_75t_L g8224 ( 
.A(n_8179),
.B(n_612),
.Y(n_8224)
);

NAND2xp5_ASAP7_75t_SL g8225 ( 
.A(n_8204),
.B(n_8205),
.Y(n_8225)
);

INVx2_ASAP7_75t_L g8226 ( 
.A(n_8195),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_8183),
.Y(n_8227)
);

AOI21xp33_ASAP7_75t_L g8228 ( 
.A1(n_8177),
.A2(n_612),
.B(n_613),
.Y(n_8228)
);

A2O1A1O1Ixp25_ASAP7_75t_L g8229 ( 
.A1(n_8208),
.A2(n_613),
.B(n_614),
.C(n_615),
.D(n_616),
.Y(n_8229)
);

NOR2xp33_ASAP7_75t_SL g8230 ( 
.A(n_8182),
.B(n_614),
.Y(n_8230)
);

OAI22xp5_ASAP7_75t_L g8231 ( 
.A1(n_8196),
.A2(n_615),
.B1(n_616),
.B2(n_617),
.Y(n_8231)
);

O2A1O1Ixp33_ASAP7_75t_L g8232 ( 
.A1(n_8198),
.A2(n_617),
.B(n_619),
.C(n_623),
.Y(n_8232)
);

NOR2xp33_ASAP7_75t_L g8233 ( 
.A(n_8193),
.B(n_619),
.Y(n_8233)
);

INVx1_ASAP7_75t_L g8234 ( 
.A(n_8201),
.Y(n_8234)
);

AOI22xp33_ASAP7_75t_SL g8235 ( 
.A1(n_8206),
.A2(n_624),
.B1(n_625),
.B2(n_626),
.Y(n_8235)
);

INVx1_ASAP7_75t_L g8236 ( 
.A(n_8210),
.Y(n_8236)
);

NOR3x1_ASAP7_75t_L g8237 ( 
.A(n_8222),
.B(n_8187),
.C(n_8186),
.Y(n_8237)
);

AOI31xp33_ASAP7_75t_L g8238 ( 
.A1(n_8220),
.A2(n_8191),
.A3(n_8203),
.B(n_8207),
.Y(n_8238)
);

AOI21xp5_ASAP7_75t_L g8239 ( 
.A1(n_8213),
.A2(n_8225),
.B(n_8232),
.Y(n_8239)
);

INVx1_ASAP7_75t_L g8240 ( 
.A(n_8211),
.Y(n_8240)
);

NOR3xp33_ASAP7_75t_L g8241 ( 
.A(n_8219),
.B(n_8200),
.C(n_625),
.Y(n_8241)
);

AND2x2_ASAP7_75t_L g8242 ( 
.A(n_8226),
.B(n_8224),
.Y(n_8242)
);

INVx1_ASAP7_75t_L g8243 ( 
.A(n_8216),
.Y(n_8243)
);

NOR3x1_ASAP7_75t_L g8244 ( 
.A(n_8215),
.B(n_624),
.C(n_627),
.Y(n_8244)
);

AOI221xp5_ASAP7_75t_L g8245 ( 
.A1(n_8228),
.A2(n_627),
.B1(n_628),
.B2(n_629),
.C(n_630),
.Y(n_8245)
);

OAI211xp5_ASAP7_75t_SL g8246 ( 
.A1(n_8234),
.A2(n_629),
.B(n_631),
.C(n_633),
.Y(n_8246)
);

NOR3xp33_ASAP7_75t_L g8247 ( 
.A(n_8214),
.B(n_633),
.C(n_635),
.Y(n_8247)
);

NOR2xp33_ASAP7_75t_SL g8248 ( 
.A(n_8212),
.B(n_635),
.Y(n_8248)
);

INVx1_ASAP7_75t_L g8249 ( 
.A(n_8229),
.Y(n_8249)
);

NAND3xp33_ASAP7_75t_SL g8250 ( 
.A(n_8223),
.B(n_636),
.C(n_638),
.Y(n_8250)
);

NOR3xp33_ASAP7_75t_L g8251 ( 
.A(n_8227),
.B(n_636),
.C(n_639),
.Y(n_8251)
);

INVx1_ASAP7_75t_L g8252 ( 
.A(n_8233),
.Y(n_8252)
);

NAND2xp5_ASAP7_75t_L g8253 ( 
.A(n_8209),
.B(n_639),
.Y(n_8253)
);

NOR2xp33_ASAP7_75t_L g8254 ( 
.A(n_8230),
.B(n_640),
.Y(n_8254)
);

AOI211xp5_ASAP7_75t_L g8255 ( 
.A1(n_8221),
.A2(n_641),
.B(n_642),
.C(n_644),
.Y(n_8255)
);

NAND3xp33_ASAP7_75t_L g8256 ( 
.A(n_8217),
.B(n_641),
.C(n_642),
.Y(n_8256)
);

OAI22xp33_ASAP7_75t_L g8257 ( 
.A1(n_8218),
.A2(n_644),
.B1(n_645),
.B2(n_646),
.Y(n_8257)
);

NAND2xp5_ASAP7_75t_L g8258 ( 
.A(n_8235),
.B(n_646),
.Y(n_8258)
);

NOR2xp33_ASAP7_75t_L g8259 ( 
.A(n_8231),
.B(n_647),
.Y(n_8259)
);

NAND2xp5_ASAP7_75t_SL g8260 ( 
.A(n_8211),
.B(n_647),
.Y(n_8260)
);

OAI21xp33_ASAP7_75t_L g8261 ( 
.A1(n_8249),
.A2(n_648),
.B(n_649),
.Y(n_8261)
);

NAND2xp5_ASAP7_75t_L g8262 ( 
.A(n_8251),
.B(n_648),
.Y(n_8262)
);

NAND2xp5_ASAP7_75t_L g8263 ( 
.A(n_8255),
.B(n_651),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_8258),
.Y(n_8264)
);

NAND4xp25_ASAP7_75t_L g8265 ( 
.A(n_8244),
.B(n_651),
.C(n_652),
.D(n_653),
.Y(n_8265)
);

AOI21xp5_ASAP7_75t_L g8266 ( 
.A1(n_8260),
.A2(n_653),
.B(n_654),
.Y(n_8266)
);

NAND4xp25_ASAP7_75t_L g8267 ( 
.A(n_8237),
.B(n_655),
.C(n_656),
.D(n_657),
.Y(n_8267)
);

OR2x2_ASAP7_75t_L g8268 ( 
.A(n_8250),
.B(n_655),
.Y(n_8268)
);

INVxp67_ASAP7_75t_SL g8269 ( 
.A(n_8253),
.Y(n_8269)
);

OR2x2_ASAP7_75t_L g8270 ( 
.A(n_8256),
.B(n_657),
.Y(n_8270)
);

NOR4xp25_ASAP7_75t_L g8271 ( 
.A(n_8243),
.B(n_659),
.C(n_660),
.D(n_662),
.Y(n_8271)
);

OAI211xp5_ASAP7_75t_SL g8272 ( 
.A1(n_8239),
.A2(n_659),
.B(n_660),
.C(n_664),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_8254),
.Y(n_8273)
);

NAND2x1_ASAP7_75t_L g8274 ( 
.A(n_8238),
.B(n_665),
.Y(n_8274)
);

OAI21xp5_ASAP7_75t_SL g8275 ( 
.A1(n_8245),
.A2(n_8242),
.B(n_8240),
.Y(n_8275)
);

HB1xp67_ASAP7_75t_L g8276 ( 
.A(n_8259),
.Y(n_8276)
);

INVx1_ASAP7_75t_L g8277 ( 
.A(n_8246),
.Y(n_8277)
);

NAND2xp5_ASAP7_75t_L g8278 ( 
.A(n_8257),
.B(n_665),
.Y(n_8278)
);

BUFx4f_ASAP7_75t_SL g8279 ( 
.A(n_8236),
.Y(n_8279)
);

INVx1_ASAP7_75t_L g8280 ( 
.A(n_8248),
.Y(n_8280)
);

NOR2xp33_ASAP7_75t_L g8281 ( 
.A(n_8252),
.B(n_666),
.Y(n_8281)
);

NAND2xp5_ASAP7_75t_L g8282 ( 
.A(n_8247),
.B(n_666),
.Y(n_8282)
);

AOI221xp5_ASAP7_75t_L g8283 ( 
.A1(n_8241),
.A2(n_667),
.B1(n_668),
.B2(n_669),
.C(n_670),
.Y(n_8283)
);

NOR3x1_ASAP7_75t_L g8284 ( 
.A(n_8250),
.B(n_667),
.C(n_668),
.Y(n_8284)
);

AOI222xp33_ASAP7_75t_L g8285 ( 
.A1(n_8250),
.A2(n_670),
.B1(n_671),
.B2(n_672),
.C1(n_673),
.C2(n_674),
.Y(n_8285)
);

OAI211xp5_ASAP7_75t_L g8286 ( 
.A1(n_8245),
.A2(n_671),
.B(n_674),
.C(n_675),
.Y(n_8286)
);

NAND3xp33_ASAP7_75t_L g8287 ( 
.A(n_8245),
.B(n_676),
.C(n_678),
.Y(n_8287)
);

AOI211x1_ASAP7_75t_L g8288 ( 
.A1(n_8238),
.A2(n_678),
.B(n_679),
.C(n_680),
.Y(n_8288)
);

AND2x2_ASAP7_75t_L g8289 ( 
.A(n_8249),
.B(n_679),
.Y(n_8289)
);

NAND2xp5_ASAP7_75t_L g8290 ( 
.A(n_8251),
.B(n_680),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_8289),
.Y(n_8291)
);

NAND2xp5_ASAP7_75t_L g8292 ( 
.A(n_8261),
.B(n_681),
.Y(n_8292)
);

NOR3xp33_ASAP7_75t_SL g8293 ( 
.A(n_8275),
.B(n_681),
.C(n_682),
.Y(n_8293)
);

OAI211xp5_ASAP7_75t_L g8294 ( 
.A1(n_8285),
.A2(n_683),
.B(n_686),
.C(n_687),
.Y(n_8294)
);

OAI211xp5_ASAP7_75t_L g8295 ( 
.A1(n_8274),
.A2(n_686),
.B(n_688),
.C(n_689),
.Y(n_8295)
);

XNOR2x2_ASAP7_75t_L g8296 ( 
.A(n_8288),
.B(n_691),
.Y(n_8296)
);

NOR3xp33_ASAP7_75t_L g8297 ( 
.A(n_8280),
.B(n_693),
.C(n_695),
.Y(n_8297)
);

AOI22xp5_ASAP7_75t_L g8298 ( 
.A1(n_8272),
.A2(n_695),
.B1(n_696),
.B2(n_697),
.Y(n_8298)
);

NOR2xp33_ASAP7_75t_L g8299 ( 
.A(n_8265),
.B(n_697),
.Y(n_8299)
);

XNOR2x1_ASAP7_75t_L g8300 ( 
.A(n_8268),
.B(n_698),
.Y(n_8300)
);

NAND2xp5_ASAP7_75t_SL g8301 ( 
.A(n_8271),
.B(n_699),
.Y(n_8301)
);

AND2x4_ASAP7_75t_L g8302 ( 
.A(n_8284),
.B(n_699),
.Y(n_8302)
);

AOI211x1_ASAP7_75t_L g8303 ( 
.A1(n_8287),
.A2(n_700),
.B(n_701),
.C(n_703),
.Y(n_8303)
);

INVx2_ASAP7_75t_SL g8304 ( 
.A(n_8270),
.Y(n_8304)
);

NOR3x1_ASAP7_75t_L g8305 ( 
.A(n_8267),
.B(n_700),
.C(n_704),
.Y(n_8305)
);

NAND3xp33_ASAP7_75t_L g8306 ( 
.A(n_8283),
.B(n_8282),
.C(n_8266),
.Y(n_8306)
);

OAI21xp5_ASAP7_75t_L g8307 ( 
.A1(n_8263),
.A2(n_705),
.B(n_706),
.Y(n_8307)
);

NOR3xp33_ASAP7_75t_L g8308 ( 
.A(n_8264),
.B(n_705),
.C(n_706),
.Y(n_8308)
);

NOR2x1_ASAP7_75t_L g8309 ( 
.A(n_8286),
.B(n_707),
.Y(n_8309)
);

AOI21xp5_ASAP7_75t_L g8310 ( 
.A1(n_8262),
.A2(n_707),
.B(n_708),
.Y(n_8310)
);

AND2x2_ASAP7_75t_L g8311 ( 
.A(n_8277),
.B(n_708),
.Y(n_8311)
);

NAND4xp25_ASAP7_75t_SL g8312 ( 
.A(n_8290),
.B(n_709),
.C(n_710),
.D(n_711),
.Y(n_8312)
);

NOR2xp67_ASAP7_75t_SL g8313 ( 
.A(n_8276),
.B(n_710),
.Y(n_8313)
);

INVxp33_ASAP7_75t_L g8314 ( 
.A(n_8281),
.Y(n_8314)
);

NAND2xp5_ASAP7_75t_L g8315 ( 
.A(n_8273),
.B(n_712),
.Y(n_8315)
);

INVx1_ASAP7_75t_L g8316 ( 
.A(n_8313),
.Y(n_8316)
);

NOR2x1_ASAP7_75t_L g8317 ( 
.A(n_8312),
.B(n_8278),
.Y(n_8317)
);

NOR3xp33_ASAP7_75t_L g8318 ( 
.A(n_8311),
.B(n_8269),
.C(n_8279),
.Y(n_8318)
);

NOR2x1_ASAP7_75t_L g8319 ( 
.A(n_8295),
.B(n_713),
.Y(n_8319)
);

XNOR2x1_ASAP7_75t_L g8320 ( 
.A(n_8296),
.B(n_713),
.Y(n_8320)
);

NOR2xp33_ASAP7_75t_L g8321 ( 
.A(n_8294),
.B(n_714),
.Y(n_8321)
);

NOR2x1_ASAP7_75t_L g8322 ( 
.A(n_8301),
.B(n_714),
.Y(n_8322)
);

OAI21xp33_ASAP7_75t_L g8323 ( 
.A1(n_8293),
.A2(n_715),
.B(n_716),
.Y(n_8323)
);

NAND3xp33_ASAP7_75t_SL g8324 ( 
.A(n_8307),
.B(n_715),
.C(n_716),
.Y(n_8324)
);

INVx2_ASAP7_75t_L g8325 ( 
.A(n_8315),
.Y(n_8325)
);

AND2x2_ASAP7_75t_L g8326 ( 
.A(n_8305),
.B(n_717),
.Y(n_8326)
);

INVx1_ASAP7_75t_L g8327 ( 
.A(n_8292),
.Y(n_8327)
);

NAND2xp5_ASAP7_75t_L g8328 ( 
.A(n_8297),
.B(n_718),
.Y(n_8328)
);

NAND4xp75_ASAP7_75t_L g8329 ( 
.A(n_8309),
.B(n_718),
.C(n_720),
.D(n_723),
.Y(n_8329)
);

NOR2x1_ASAP7_75t_L g8330 ( 
.A(n_8300),
.B(n_720),
.Y(n_8330)
);

NAND2xp5_ASAP7_75t_L g8331 ( 
.A(n_8308),
.B(n_729),
.Y(n_8331)
);

NOR2x1_ASAP7_75t_L g8332 ( 
.A(n_8291),
.B(n_2415),
.Y(n_8332)
);

NOR3x1_ASAP7_75t_L g8333 ( 
.A(n_8306),
.B(n_736),
.C(n_737),
.Y(n_8333)
);

AOI221xp5_ASAP7_75t_L g8334 ( 
.A1(n_8323),
.A2(n_8303),
.B1(n_8299),
.B2(n_8302),
.C(n_8314),
.Y(n_8334)
);

OAI311xp33_ASAP7_75t_L g8335 ( 
.A1(n_8316),
.A2(n_8298),
.A3(n_8302),
.B1(n_8304),
.C1(n_8310),
.Y(n_8335)
);

AOI211xp5_ASAP7_75t_L g8336 ( 
.A1(n_8324),
.A2(n_738),
.B(n_2815),
.C(n_2804),
.Y(n_8336)
);

NAND2xp5_ASAP7_75t_L g8337 ( 
.A(n_8326),
.B(n_2745),
.Y(n_8337)
);

AOI22xp5_ASAP7_75t_L g8338 ( 
.A1(n_8318),
.A2(n_2804),
.B1(n_2763),
.B2(n_2784),
.Y(n_8338)
);

INVx1_ASAP7_75t_SL g8339 ( 
.A(n_8320),
.Y(n_8339)
);

OAI21xp5_ASAP7_75t_L g8340 ( 
.A1(n_8330),
.A2(n_2187),
.B(n_2457),
.Y(n_8340)
);

NOR3xp33_ASAP7_75t_SL g8341 ( 
.A(n_8335),
.B(n_8321),
.C(n_8327),
.Y(n_8341)
);

NOR3xp33_ASAP7_75t_L g8342 ( 
.A(n_8339),
.B(n_8325),
.C(n_8322),
.Y(n_8342)
);

NOR3xp33_ASAP7_75t_L g8343 ( 
.A(n_8334),
.B(n_8317),
.C(n_8328),
.Y(n_8343)
);

NOR2x1p5_ASAP7_75t_L g8344 ( 
.A(n_8337),
.B(n_8329),
.Y(n_8344)
);

NAND2xp5_ASAP7_75t_L g8345 ( 
.A(n_8336),
.B(n_8319),
.Y(n_8345)
);

AND2x2_ASAP7_75t_L g8346 ( 
.A(n_8341),
.B(n_8331),
.Y(n_8346)
);

AOI22xp5_ASAP7_75t_L g8347 ( 
.A1(n_8342),
.A2(n_8343),
.B1(n_8344),
.B2(n_8345),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_8345),
.Y(n_8348)
);

AND2x4_ASAP7_75t_L g8349 ( 
.A(n_8341),
.B(n_8333),
.Y(n_8349)
);

AOI22xp5_ASAP7_75t_L g8350 ( 
.A1(n_8342),
.A2(n_8338),
.B1(n_8332),
.B2(n_8340),
.Y(n_8350)
);

NAND4xp75_ASAP7_75t_L g8351 ( 
.A(n_8341),
.B(n_2168),
.C(n_2175),
.D(n_2176),
.Y(n_8351)
);

INVx1_ASAP7_75t_L g8352 ( 
.A(n_8345),
.Y(n_8352)
);

INVxp67_ASAP7_75t_L g8353 ( 
.A(n_8345),
.Y(n_8353)
);

INVx1_ASAP7_75t_L g8354 ( 
.A(n_8345),
.Y(n_8354)
);

NOR2x1_ASAP7_75t_SL g8355 ( 
.A(n_8345),
.B(n_2815),
.Y(n_8355)
);

NAND2xp33_ASAP7_75t_L g8356 ( 
.A(n_8348),
.B(n_2815),
.Y(n_8356)
);

XNOR2xp5_ASAP7_75t_L g8357 ( 
.A(n_8347),
.B(n_8349),
.Y(n_8357)
);

INVx2_ASAP7_75t_L g8358 ( 
.A(n_8351),
.Y(n_8358)
);

BUFx6f_ASAP7_75t_L g8359 ( 
.A(n_8346),
.Y(n_8359)
);

XNOR2x1_ASAP7_75t_L g8360 ( 
.A(n_8352),
.B(n_2745),
.Y(n_8360)
);

NOR2xp67_ASAP7_75t_L g8361 ( 
.A(n_8353),
.B(n_2312),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_8355),
.Y(n_8362)
);

NAND2xp5_ASAP7_75t_SL g8363 ( 
.A(n_8354),
.B(n_2815),
.Y(n_8363)
);

NOR2x1_ASAP7_75t_L g8364 ( 
.A(n_8350),
.B(n_2168),
.Y(n_8364)
);

NOR3xp33_ASAP7_75t_L g8365 ( 
.A(n_8353),
.B(n_2276),
.C(n_2372),
.Y(n_8365)
);

HB1xp67_ASAP7_75t_L g8366 ( 
.A(n_8349),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_8355),
.Y(n_8367)
);

INVx2_ASAP7_75t_L g8368 ( 
.A(n_8351),
.Y(n_8368)
);

NOR2x1_ASAP7_75t_L g8369 ( 
.A(n_8351),
.B(n_2168),
.Y(n_8369)
);

BUFx2_ASAP7_75t_L g8370 ( 
.A(n_8349),
.Y(n_8370)
);

NOR4xp25_ASAP7_75t_L g8371 ( 
.A(n_8362),
.B(n_2276),
.C(n_2372),
.D(n_2175),
.Y(n_8371)
);

NAND3xp33_ASAP7_75t_SL g8372 ( 
.A(n_8370),
.B(n_2276),
.C(n_2372),
.Y(n_8372)
);

AOI21xp5_ASAP7_75t_L g8373 ( 
.A1(n_8357),
.A2(n_2312),
.B(n_2457),
.Y(n_8373)
);

AOI211xp5_ASAP7_75t_L g8374 ( 
.A1(n_8366),
.A2(n_2175),
.B(n_2176),
.C(n_2213),
.Y(n_8374)
);

INVx2_ASAP7_75t_SL g8375 ( 
.A(n_8359),
.Y(n_8375)
);

NAND4xp25_ASAP7_75t_L g8376 ( 
.A(n_8365),
.B(n_2457),
.C(n_2312),
.D(n_2175),
.Y(n_8376)
);

NAND2xp5_ASAP7_75t_L g8377 ( 
.A(n_8375),
.B(n_8359),
.Y(n_8377)
);

OR2x2_ASAP7_75t_L g8378 ( 
.A(n_8376),
.B(n_8360),
.Y(n_8378)
);

AOI22x1_ASAP7_75t_L g8379 ( 
.A1(n_8373),
.A2(n_8368),
.B1(n_8358),
.B2(n_8367),
.Y(n_8379)
);

AOI22xp5_ASAP7_75t_L g8380 ( 
.A1(n_8372),
.A2(n_8363),
.B1(n_8369),
.B2(n_8356),
.Y(n_8380)
);

NAND2xp5_ASAP7_75t_L g8381 ( 
.A(n_8374),
.B(n_8361),
.Y(n_8381)
);

OAI22xp5_ASAP7_75t_L g8382 ( 
.A1(n_8377),
.A2(n_8380),
.B1(n_8379),
.B2(n_8378),
.Y(n_8382)
);

INVx2_ASAP7_75t_L g8383 ( 
.A(n_8381),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_8377),
.Y(n_8384)
);

INVx2_ASAP7_75t_L g8385 ( 
.A(n_8379),
.Y(n_8385)
);

NAND2xp5_ASAP7_75t_L g8386 ( 
.A(n_8377),
.B(n_8364),
.Y(n_8386)
);

OR2x2_ASAP7_75t_L g8387 ( 
.A(n_8377),
.B(n_8371),
.Y(n_8387)
);

INVx2_ASAP7_75t_L g8388 ( 
.A(n_8379),
.Y(n_8388)
);

XOR2x2_ASAP7_75t_L g8389 ( 
.A(n_8377),
.B(n_2276),
.Y(n_8389)
);

AOI22xp33_ASAP7_75t_L g8390 ( 
.A1(n_8379),
.A2(n_2763),
.B1(n_2784),
.B2(n_2804),
.Y(n_8390)
);

NAND2xp5_ASAP7_75t_L g8391 ( 
.A(n_8377),
.B(n_2299),
.Y(n_8391)
);

INVxp67_ASAP7_75t_L g8392 ( 
.A(n_8377),
.Y(n_8392)
);

INVx1_ASAP7_75t_L g8393 ( 
.A(n_8377),
.Y(n_8393)
);

AOI22x1_ASAP7_75t_L g8394 ( 
.A1(n_8378),
.A2(n_2305),
.B1(n_2300),
.B2(n_2328),
.Y(n_8394)
);

INVx4_ASAP7_75t_L g8395 ( 
.A(n_8378),
.Y(n_8395)
);

OA22x2_ASAP7_75t_L g8396 ( 
.A1(n_8384),
.A2(n_2213),
.B1(n_2206),
.B2(n_2200),
.Y(n_8396)
);

BUFx2_ASAP7_75t_L g8397 ( 
.A(n_8392),
.Y(n_8397)
);

AO21x2_ASAP7_75t_L g8398 ( 
.A1(n_8393),
.A2(n_2205),
.B(n_2222),
.Y(n_8398)
);

NOR2x1_ASAP7_75t_L g8399 ( 
.A(n_8385),
.B(n_2299),
.Y(n_8399)
);

OA21x2_ASAP7_75t_L g8400 ( 
.A1(n_8388),
.A2(n_2213),
.B(n_2206),
.Y(n_8400)
);

BUFx2_ASAP7_75t_L g8401 ( 
.A(n_8395),
.Y(n_8401)
);

INVx1_ASAP7_75t_L g8402 ( 
.A(n_8389),
.Y(n_8402)
);

CKINVDCx20_ASAP7_75t_R g8403 ( 
.A(n_8382),
.Y(n_8403)
);

XOR2xp5_ASAP7_75t_L g8404 ( 
.A(n_8383),
.B(n_2305),
.Y(n_8404)
);

INVx4_ASAP7_75t_L g8405 ( 
.A(n_8387),
.Y(n_8405)
);

INVx3_ASAP7_75t_L g8406 ( 
.A(n_8401),
.Y(n_8406)
);

NAND2xp5_ASAP7_75t_L g8407 ( 
.A(n_8397),
.B(n_8391),
.Y(n_8407)
);

INVx2_ASAP7_75t_SL g8408 ( 
.A(n_8403),
.Y(n_8408)
);

NAND2xp5_ASAP7_75t_L g8409 ( 
.A(n_8404),
.B(n_8386),
.Y(n_8409)
);

NOR2xp33_ASAP7_75t_L g8410 ( 
.A(n_8405),
.B(n_8390),
.Y(n_8410)
);

AOI22xp5_ASAP7_75t_L g8411 ( 
.A1(n_8402),
.A2(n_8394),
.B1(n_2372),
.B2(n_2213),
.Y(n_8411)
);

INVx1_ASAP7_75t_L g8412 ( 
.A(n_8399),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_8398),
.Y(n_8413)
);

NAND2xp5_ASAP7_75t_L g8414 ( 
.A(n_8406),
.B(n_8400),
.Y(n_8414)
);

AOI21xp5_ASAP7_75t_L g8415 ( 
.A1(n_8408),
.A2(n_8396),
.B(n_2457),
.Y(n_8415)
);

AOI22xp5_ASAP7_75t_L g8416 ( 
.A1(n_8410),
.A2(n_2175),
.B1(n_2176),
.B2(n_2213),
.Y(n_8416)
);

NAND2xp5_ASAP7_75t_L g8417 ( 
.A(n_8407),
.B(n_2299),
.Y(n_8417)
);

INVx1_ASAP7_75t_SL g8418 ( 
.A(n_8414),
.Y(n_8418)
);

INVx1_ASAP7_75t_L g8419 ( 
.A(n_8417),
.Y(n_8419)
);

NAND2xp5_ASAP7_75t_L g8420 ( 
.A(n_8418),
.B(n_8409),
.Y(n_8420)
);

NOR2xp33_ASAP7_75t_L g8421 ( 
.A(n_8419),
.B(n_8413),
.Y(n_8421)
);

AOI222xp33_ASAP7_75t_L g8422 ( 
.A1(n_8420),
.A2(n_8412),
.B1(n_8415),
.B2(n_8411),
.C1(n_8416),
.C2(n_2176),
.Y(n_8422)
);

OAI21xp5_ASAP7_75t_L g8423 ( 
.A1(n_8421),
.A2(n_2312),
.B(n_2457),
.Y(n_8423)
);

AOI22xp33_ASAP7_75t_L g8424 ( 
.A1(n_8421),
.A2(n_2176),
.B1(n_2328),
.B2(n_2305),
.Y(n_8424)
);

NAND2xp5_ASAP7_75t_L g8425 ( 
.A(n_8422),
.B(n_2200),
.Y(n_8425)
);

AOI221xp5_ASAP7_75t_L g8426 ( 
.A1(n_8424),
.A2(n_2300),
.B1(n_2299),
.B2(n_2305),
.C(n_2328),
.Y(n_8426)
);

AOI22xp5_ASAP7_75t_L g8427 ( 
.A1(n_8423),
.A2(n_2200),
.B1(n_2206),
.B2(n_2299),
.Y(n_8427)
);

OAI21xp5_ASAP7_75t_L g8428 ( 
.A1(n_8425),
.A2(n_8427),
.B(n_8426),
.Y(n_8428)
);

OAI21xp5_ASAP7_75t_L g8429 ( 
.A1(n_8425),
.A2(n_2312),
.B(n_2205),
.Y(n_8429)
);

OAI21xp33_ASAP7_75t_SL g8430 ( 
.A1(n_8425),
.A2(n_2300),
.B(n_2305),
.Y(n_8430)
);

AOI21xp33_ASAP7_75t_SL g8431 ( 
.A1(n_8425),
.A2(n_2222),
.B(n_2205),
.Y(n_8431)
);

AOI31xp67_ASAP7_75t_L g8432 ( 
.A1(n_8428),
.A2(n_2222),
.A3(n_2205),
.B(n_2271),
.Y(n_8432)
);

OAI21xp5_ASAP7_75t_L g8433 ( 
.A1(n_8430),
.A2(n_2222),
.B(n_2205),
.Y(n_8433)
);

AOI21xp5_ASAP7_75t_L g8434 ( 
.A1(n_8429),
.A2(n_2222),
.B(n_2328),
.Y(n_8434)
);

AOI22xp33_ASAP7_75t_L g8435 ( 
.A1(n_8434),
.A2(n_8431),
.B1(n_2328),
.B2(n_2300),
.Y(n_8435)
);

AOI222xp33_ASAP7_75t_L g8436 ( 
.A1(n_8433),
.A2(n_2300),
.B1(n_2200),
.B2(n_2206),
.C1(n_2241),
.C2(n_2251),
.Y(n_8436)
);

NOR2x1p5_ASAP7_75t_L g8437 ( 
.A(n_8432),
.B(n_2206),
.Y(n_8437)
);

AO21x2_ASAP7_75t_L g8438 ( 
.A1(n_8437),
.A2(n_2275),
.B(n_2271),
.Y(n_8438)
);

NOR2xp33_ASAP7_75t_L g8439 ( 
.A(n_8435),
.B(n_2200),
.Y(n_8439)
);

AOI221xp5_ASAP7_75t_L g8440 ( 
.A1(n_8439),
.A2(n_8436),
.B1(n_2241),
.B2(n_2251),
.C(n_2261),
.Y(n_8440)
);

AOI22xp33_ASAP7_75t_L g8441 ( 
.A1(n_8440),
.A2(n_8438),
.B1(n_2275),
.B2(n_2271),
.Y(n_8441)
);

AOI211xp5_ASAP7_75t_L g8442 ( 
.A1(n_8441),
.A2(n_2277),
.B(n_2241),
.C(n_2251),
.Y(n_8442)
);


endmodule