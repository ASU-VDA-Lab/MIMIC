module real_jpeg_13818_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_65),
.B1(n_67),
.B2(n_72),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_72),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_8),
.A2(n_65),
.B1(n_67),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_8),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_91),
.Y(n_110)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_34),
.B(n_35),
.C(n_40),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_10),
.A2(n_37),
.B1(n_65),
.B2(n_67),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_10),
.A2(n_48),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_10),
.B(n_81),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_60),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_11),
.A2(n_60),
.B1(n_65),
.B2(n_67),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_60),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_13),
.A2(n_52),
.B1(n_65),
.B2(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_14),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_65),
.B1(n_67),
.B2(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_83),
.Y(n_139)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_114),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_112),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_94),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_46),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_21)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_23),
.B(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_23),
.A2(n_27),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_23),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_24),
.A2(n_25),
.B1(n_87),
.B2(n_88),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_24),
.B(n_37),
.C(n_88),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_24),
.B(n_143),
.Y(n_142)
);

CKINVDCx6p67_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_27),
.B(n_110),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_48),
.B(n_49),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_37),
.B(n_39),
.CON(n_107),
.SN(n_107)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_37),
.B(n_48),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_37),
.B(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_39),
.B1(n_64),
.B2(n_68),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_38),
.B(n_65),
.C(n_68),
.Y(n_108)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.C(n_57),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_53),
.B1(n_54),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_51),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_137),
.B1(n_145),
.B2(n_146),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_70),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_62),
.B1(n_81),
.B2(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_71),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

OA22x2_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_67),
.B(n_106),
.C(n_108),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_67),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_67),
.B(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B(n_92),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_101),
.B1(n_103),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_103),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_85),
.A2(n_103),
.B1(n_122),
.B2(n_132),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.C(n_104),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_104),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_102),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_109),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_123),
.B(n_168),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_118),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_121),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_163),
.B(n_167),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_152),
.B(n_162),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_140),
.B(n_151),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_135),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_133),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_146),
.B(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_147),
.B(n_150),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_154),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_158),
.C(n_161),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_166),
.Y(n_167)
);


endmodule