module fake_jpeg_11227_n_638 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_638);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_638;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_64),
.B(n_118),
.Y(n_146)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_30),
.A2(n_9),
.B(n_1),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_68),
.B(n_45),
.C(n_46),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_70),
.Y(n_174)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_77),
.B(n_92),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_89),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_10),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_31),
.B(n_10),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_15),
.Y(n_134)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_100),
.Y(n_194)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_31),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_126),
.Y(n_144)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_105),
.Y(n_197)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_114),
.B(n_119),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_22),
.Y(n_120)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_32),
.Y(n_123)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_33),
.B(n_8),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_134),
.B(n_13),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_140),
.B(n_158),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_38),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_145),
.B(n_171),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_72),
.A2(n_21),
.B1(n_45),
.B2(n_56),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_149),
.A2(n_195),
.B1(n_198),
.B2(n_204),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_73),
.A2(n_21),
.B1(n_39),
.B2(n_54),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_150),
.A2(n_155),
.B1(n_162),
.B2(n_212),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_74),
.A2(n_60),
.B1(n_59),
.B2(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_33),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_55),
.B1(n_53),
.B2(n_47),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_161),
.A2(n_183),
.B(n_189),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_75),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_50),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_169),
.B(n_177),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_50),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_104),
.B(n_46),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_202),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_56),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_65),
.A2(n_55),
.B1(n_53),
.B2(n_47),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_67),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_84),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_76),
.A2(n_42),
.B1(n_41),
.B2(n_0),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_99),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_106),
.B(n_11),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_112),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_122),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_213),
.Y(n_279)
);

HAxp5_ASAP7_75t_SL g209 ( 
.A(n_67),
.B(n_11),
.CON(n_209),
.SN(n_209)
);

NAND2x1_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_117),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_81),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_SL g314 ( 
.A(n_218),
.B(n_166),
.C(n_15),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_149),
.A2(n_87),
.B1(n_86),
.B2(n_83),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_219),
.A2(n_234),
.B1(n_247),
.B2(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_220),
.Y(n_319)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_221),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_223),
.Y(n_305)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_224),
.Y(n_316)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_226),
.Y(n_330)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_227),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_107),
.B1(n_116),
.B2(n_115),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g341 ( 
.A1(n_228),
.A2(n_253),
.B1(n_266),
.B2(n_280),
.Y(n_341)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_130),
.B(n_123),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_230),
.Y(n_302)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_231),
.Y(n_321)
);

NAND2x1_ASAP7_75t_SL g233 ( 
.A(n_210),
.B(n_78),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_233),
.A2(n_283),
.B(n_0),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_127),
.B1(n_124),
.B2(n_120),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_93),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_237),
.B(n_249),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_146),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_238),
.B(n_243),
.Y(n_293)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_239),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_164),
.Y(n_240)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_242),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_205),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g342 ( 
.A(n_246),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_204),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_248),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_139),
.B(n_16),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_250),
.Y(n_333)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_157),
.A2(n_160),
.B1(n_209),
.B2(n_147),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_144),
.B(n_108),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_254),
.B(n_256),
.Y(n_318)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_132),
.Y(n_255)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_18),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_138),
.B(n_18),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_259),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_133),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_156),
.B(n_102),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_270),
.Y(n_317)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_191),
.B(n_118),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_148),
.B(n_118),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_186),
.A2(n_113),
.B1(n_117),
.B2(n_70),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_136),
.Y(n_268)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_183),
.A2(n_36),
.B1(n_78),
.B2(n_7),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_133),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_154),
.B(n_5),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_271),
.B(n_273),
.Y(n_328)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_131),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_272),
.A2(n_277),
.B1(n_284),
.B2(n_285),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_197),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_170),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_186),
.A2(n_36),
.B1(n_5),
.B2(n_8),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_161),
.B(n_5),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_286),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_179),
.B(n_215),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_168),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_288),
.Y(n_324)
);

CKINVDCx12_ASAP7_75t_R g288 ( 
.A(n_136),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_193),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_291),
.Y(n_327)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_181),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_181),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_201),
.B1(n_182),
.B2(n_190),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_196),
.B1(n_153),
.B2(n_189),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_344),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_198),
.B(n_192),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_296),
.A2(n_285),
.B(n_272),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_219),
.A2(n_153),
.B1(n_196),
.B2(n_135),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_299),
.A2(n_306),
.B1(n_242),
.B2(n_268),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_234),
.A2(n_176),
.B1(n_194),
.B2(n_141),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_312),
.A2(n_343),
.B1(n_351),
.B2(n_229),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_230),
.C(n_218),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_274),
.A2(n_233),
.B1(n_278),
.B2(n_232),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_338),
.A2(n_340),
.B1(n_230),
.B2(n_262),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_241),
.B(n_201),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_345),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_220),
.A2(n_182),
.B1(n_142),
.B2(n_143),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g343 ( 
.A1(n_247),
.A2(n_180),
.B1(n_206),
.B2(n_143),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_222),
.B(n_0),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_279),
.B(n_15),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_240),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_292),
.A2(n_289),
.B1(n_263),
.B2(n_218),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_353),
.A2(n_374),
.B(n_389),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_397),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_329),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_355),
.B(n_356),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_358),
.A2(n_335),
.B1(n_350),
.B2(n_348),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_303),
.A2(n_291),
.B1(n_286),
.B2(n_284),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_359),
.A2(n_396),
.B1(n_295),
.B2(n_342),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_324),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_360),
.B(n_361),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_300),
.A2(n_217),
.B1(n_227),
.B2(n_226),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_363),
.A2(n_366),
.B1(n_330),
.B2(n_331),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_319),
.A2(n_283),
.B(n_262),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_364),
.A2(n_372),
.B(n_376),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_300),
.A2(n_224),
.B1(n_225),
.B2(n_255),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_319),
.B(n_264),
.C(n_236),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_371),
.C(n_381),
.Y(n_420)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_264),
.C(n_236),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_373),
.B(n_377),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_324),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_294),
.Y(n_375)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_296),
.A2(n_261),
.B(n_265),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_307),
.B(n_267),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_341),
.A2(n_235),
.B1(n_277),
.B2(n_231),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_378),
.Y(n_436)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_379),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_313),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_380),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_221),
.C(n_239),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_341),
.A2(n_250),
.B1(n_290),
.B2(n_223),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_383),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_293),
.B(n_248),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_384),
.B(n_385),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_248),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_328),
.B(n_246),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_387),
.B(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_316),
.Y(n_388)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_308),
.A2(n_295),
.B1(n_323),
.B2(n_337),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_336),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_394),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_303),
.A2(n_323),
.B(n_337),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_392),
.A2(n_301),
.B(n_346),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_317),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_395),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_349),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_297),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_295),
.A2(n_343),
.B1(n_312),
.B2(n_308),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_321),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_304),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_401),
.B(n_426),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_403),
.A2(n_406),
.B1(n_412),
.B2(n_422),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_356),
.B(n_298),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_418),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_396),
.A2(n_326),
.B1(n_342),
.B2(n_309),
.Y(n_406)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_391),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_411),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_314),
.B1(n_310),
.B2(n_322),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_315),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_358),
.B1(n_363),
.B2(n_366),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_353),
.A2(n_322),
.B1(n_335),
.B2(n_346),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_352),
.B(n_393),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_428),
.A2(n_372),
.B(n_392),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_347),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_364),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_357),
.B(n_394),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_434),
.Y(n_469)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_376),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_404),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_451),
.Y(n_487)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_442),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_443),
.A2(n_449),
.B(n_453),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_369),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_444),
.B(n_446),
.C(n_458),
.Y(n_484)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_398),
.A2(n_365),
.B(n_361),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_412),
.A2(n_365),
.B1(n_360),
.B2(n_374),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_450),
.A2(n_464),
.B(n_439),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_427),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_400),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_452),
.B(n_455),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g453 ( 
.A1(n_431),
.A2(n_365),
.B(n_354),
.Y(n_453)
);

XOR2x1_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_373),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_429),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_400),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_407),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_460),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_377),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_398),
.A2(n_433),
.B1(n_402),
.B2(n_431),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_459),
.A2(n_466),
.B1(n_442),
.B2(n_438),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_434),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_403),
.A2(n_381),
.B1(n_395),
.B2(n_362),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_463),
.A2(n_420),
.B1(n_435),
.B2(n_405),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_422),
.A2(n_367),
.B1(n_355),
.B2(n_382),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_421),
.A2(n_384),
.B(n_387),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_465),
.A2(n_417),
.B(n_425),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_402),
.A2(n_385),
.B1(n_359),
.B2(n_379),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_432),
.Y(n_467)
);

NAND2x1_ASAP7_75t_SL g473 ( 
.A(n_467),
.B(n_432),
.Y(n_473)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_468),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_390),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_470),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_414),
.B(n_401),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_472),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_473),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_474),
.A2(n_478),
.B1(n_489),
.B2(n_463),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_475),
.A2(n_479),
.B1(n_482),
.B2(n_452),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_476),
.B(n_497),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_459),
.A2(n_437),
.B1(n_439),
.B2(n_441),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_453),
.A2(n_421),
.B1(n_436),
.B2(n_399),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_457),
.A2(n_436),
.B1(n_417),
.B2(n_406),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_458),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_486),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_409),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_488),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_471),
.A2(n_417),
.B1(n_424),
.B2(n_415),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_413),
.C(n_415),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_496),
.C(n_460),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_413),
.C(n_424),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_430),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_504),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_456),
.B(n_380),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_501),
.B(n_505),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_430),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_440),
.B(n_370),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_503),
.Y(n_506)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_506),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_509),
.A2(n_523),
.B1(n_525),
.B2(n_529),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_454),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_511),
.B(n_521),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_493),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_513),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_450),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_455),
.Y(n_514)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_514),
.Y(n_551)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_503),
.Y(n_515)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_515),
.Y(n_558)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_480),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_519),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_517),
.A2(n_528),
.B1(n_533),
.B2(n_478),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_518),
.B(n_520),
.Y(n_548)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_475),
.B(n_469),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_469),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_500),
.B(n_440),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_524),
.Y(n_540)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_486),
.B(n_467),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_526),
.B(n_535),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_504),
.B(n_470),
.C(n_457),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_490),
.C(n_497),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_482),
.A2(n_437),
.B1(n_466),
.B2(n_447),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_487),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_487),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_530),
.A2(n_495),
.B1(n_492),
.B2(n_499),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_473),
.B(n_447),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_531),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_479),
.A2(n_443),
.B1(n_468),
.B2(n_448),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_465),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_536),
.B(n_549),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_506),
.A2(n_494),
.B1(n_477),
.B2(n_474),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_538),
.A2(n_559),
.B1(n_397),
.B2(n_332),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_539),
.A2(n_552),
.B1(n_514),
.B2(n_532),
.Y(n_570)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_545),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_508),
.A2(n_491),
.B(n_477),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_546),
.A2(n_553),
.B(n_526),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_521),
.B(n_498),
.C(n_491),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_512),
.B(n_489),
.C(n_488),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_550),
.B(n_507),
.C(n_513),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_SL g552 ( 
.A1(n_522),
.A2(n_494),
.B(n_464),
.C(n_495),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_451),
.B(n_462),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_528),
.A2(n_425),
.B1(n_416),
.B2(n_410),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g563 ( 
.A(n_554),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_518),
.B(n_416),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_556),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_410),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_534),
.A2(n_388),
.B1(n_386),
.B2(n_397),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_375),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_510),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_544),
.A2(n_517),
.B1(n_533),
.B2(n_527),
.Y(n_561)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_561),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_562),
.B(n_568),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_565),
.A2(n_571),
.B(n_549),
.Y(n_584)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_537),
.Y(n_566)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_566),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_557),
.B(n_510),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_573),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_570),
.A2(n_552),
.B1(n_556),
.B2(n_542),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_551),
.A2(n_520),
.B(n_507),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_555),
.B(n_333),
.C(n_334),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_572),
.B(n_576),
.Y(n_595)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_553),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_578),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_547),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_321),
.Y(n_577)
);

CKINVDCx14_ASAP7_75t_R g592 ( 
.A(n_577),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_333),
.C(n_332),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_538),
.A2(n_332),
.B1(n_313),
.B2(n_305),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_563),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_541),
.B(n_320),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_580),
.B(n_552),
.Y(n_583)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_574),
.Y(n_581)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_581),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_570),
.A2(n_558),
.B1(n_536),
.B2(n_550),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_585),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_583),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_584),
.B(n_589),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_565),
.A2(n_552),
.B(n_557),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_564),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_548),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_560),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_590),
.B(n_579),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_593),
.A2(n_561),
.B1(n_568),
.B2(n_564),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_575),
.A2(n_542),
.B(n_543),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_596),
.B(n_562),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_598),
.B(n_600),
.Y(n_621)
);

INVx11_ASAP7_75t_L g601 ( 
.A(n_592),
.Y(n_601)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_601),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_584),
.A2(n_571),
.B(n_578),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_602),
.A2(n_606),
.B(n_609),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_595),
.B(n_589),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_607),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_610),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_543),
.C(n_567),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_609),
.A2(n_586),
.B(n_591),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_583),
.A2(n_572),
.B1(n_569),
.B2(n_567),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_301),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_594),
.C(n_587),
.Y(n_616)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_603),
.A2(n_585),
.B(n_596),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_613),
.A2(n_598),
.B(n_599),
.Y(n_624)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_614),
.A2(n_619),
.B(n_607),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_606),
.B(n_587),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_615),
.B(n_616),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_604),
.A2(n_586),
.B(n_581),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_620),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_624),
.B(n_628),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_621),
.B(n_601),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_625),
.Y(n_630)
);

AO21x1_ASAP7_75t_L g626 ( 
.A1(n_618),
.A2(n_591),
.B(n_607),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_626),
.A2(n_588),
.B1(n_590),
.B2(n_593),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g631 ( 
.A1(n_627),
.A2(n_612),
.B(n_617),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_621),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_622),
.C(n_623),
.Y(n_633)
);

OAI211xp5_ASAP7_75t_L g634 ( 
.A1(n_632),
.A2(n_610),
.B(n_608),
.C(n_611),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_633),
.A2(n_634),
.B1(n_629),
.B2(n_630),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_635),
.A2(n_320),
.B(n_330),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_636),
.A2(n_331),
.B(n_347),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_637),
.B(n_305),
.Y(n_638)
);


endmodule