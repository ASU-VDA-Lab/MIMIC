module fake_jpeg_31986_n_82 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_5),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_14),
.B1(n_26),
.B2(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_42),
.Y(n_44)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_13),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_39),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_34),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_29),
.C(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_55),
.Y(n_66)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_6),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_28),
.C(n_40),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_36),
.A3(n_46),
.B1(n_15),
.B2(n_9),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_60),
.C(n_57),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_36),
.B(n_16),
.C(n_27),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_65),
.B1(n_7),
.B2(n_23),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_69),
.C(n_11),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_73),
.B(n_74),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_62),
.Y(n_75)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_61),
.B(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_72),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_68),
.B1(n_64),
.B2(n_19),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_12),
.B(n_18),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_20),
.Y(n_82)
);


endmodule