module real_aes_8345_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_617;
wire n_552;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g485 ( .A(n_1), .Y(n_485) );
INVx1_ASAP7_75t_L g198 ( .A(n_2), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_3), .A2(n_36), .B1(n_170), .B2(n_494), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g209 ( .A1(n_4), .A2(n_127), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_5), .B(n_157), .Y(n_477) );
AND2x6_ASAP7_75t_L g132 ( .A(n_6), .B(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_7), .A2(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_37), .Y(n_113) );
INVx1_ASAP7_75t_L g742 ( .A(n_8), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_9), .B(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g215 ( .A(n_10), .Y(n_215) );
INVx1_ASAP7_75t_L g153 ( .A(n_11), .Y(n_153) );
INVx1_ASAP7_75t_L g481 ( .A(n_12), .Y(n_481) );
INVx1_ASAP7_75t_L g186 ( .A(n_13), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_14), .B(n_201), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_15), .B(n_149), .Y(n_544) );
AOI222xp33_ASAP7_75t_L g114 ( .A1(n_16), .A2(n_65), .B1(n_115), .B2(n_722), .C1(n_723), .C2(n_726), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_16), .Y(n_722) );
AO32x2_ASAP7_75t_L g491 ( .A1(n_17), .A2(n_148), .A3(n_157), .B1(n_463), .B2(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_18), .B(n_170), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_19), .B(n_143), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_20), .B(n_149), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_21), .A2(n_47), .B1(n_170), .B2(n_494), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_22), .B(n_127), .Y(n_126) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_23), .A2(n_74), .B1(n_170), .B2(n_201), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_24), .B(n_170), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_25), .B(n_208), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_26), .A2(n_183), .B(n_185), .C(n_187), .Y(n_182) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_28), .B(n_161), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_29), .B(n_168), .Y(n_199) );
INVx1_ASAP7_75t_L g225 ( .A(n_30), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_31), .B(n_161), .Y(n_507) );
INVx2_ASAP7_75t_L g130 ( .A(n_32), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_33), .B(n_170), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_34), .B(n_161), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_35), .A2(n_132), .B(n_135), .C(n_138), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_37), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g223 ( .A(n_38), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_39), .B(n_168), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_40), .B(n_170), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_41), .A2(n_84), .B1(n_146), .B2(n_494), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_42), .B(n_170), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_43), .B(n_170), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_44), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_45), .B(n_461), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_46), .B(n_127), .Y(n_171) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_48), .A2(n_58), .B1(n_170), .B2(n_201), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_49), .A2(n_135), .B1(n_201), .B2(n_222), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_50), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_51), .B(n_170), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_52), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_53), .B(n_170), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_54), .A2(n_213), .B(n_214), .C(n_216), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_55), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_56), .Y(n_106) );
INVx1_ASAP7_75t_L g211 ( .A(n_57), .Y(n_211) );
INVx1_ASAP7_75t_L g133 ( .A(n_59), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_60), .B(n_170), .Y(n_486) );
INVx1_ASAP7_75t_L g152 ( .A(n_61), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_62), .Y(n_104) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_63), .A2(n_100), .B1(n_737), .B2(n_748), .Y(n_99) );
AO32x2_ASAP7_75t_L g527 ( .A1(n_64), .A2(n_157), .A3(n_160), .B1(n_463), .B2(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g459 ( .A(n_66), .Y(n_459) );
INVx1_ASAP7_75t_L g502 ( .A(n_67), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_SL g233 ( .A1(n_68), .A2(n_143), .B(n_216), .C(n_234), .Y(n_233) );
INVxp67_ASAP7_75t_L g235 ( .A(n_69), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_70), .B(n_201), .Y(n_503) );
INVx1_ASAP7_75t_L g747 ( .A(n_71), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_72), .Y(n_228) );
INVx1_ASAP7_75t_L g256 ( .A(n_73), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_75), .A2(n_132), .B(n_135), .C(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_76), .B(n_494), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_77), .B(n_201), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_78), .B(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g150 ( .A(n_79), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_80), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_81), .B(n_201), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_82), .A2(n_132), .B(n_135), .C(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g109 ( .A(n_83), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g118 ( .A(n_83), .B(n_111), .Y(n_118) );
INVx2_ASAP7_75t_L g446 ( .A(n_83), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_85), .A2(n_98), .B1(n_201), .B2(n_202), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_86), .A2(n_119), .B1(n_732), .B2(n_733), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_86), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_87), .B(n_161), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_88), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_89), .A2(n_132), .B(n_135), .C(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_90), .Y(n_173) );
INVx1_ASAP7_75t_L g232 ( .A(n_91), .Y(n_232) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_92), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_93), .B(n_140), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_94), .B(n_201), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_95), .B(n_157), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_96), .A2(n_127), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_97), .B(n_747), .Y(n_746) );
AOI22x1_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_114), .B1(n_729), .B2(n_730), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g729 ( .A(n_103), .Y(n_729) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_105), .A2(n_731), .B(n_734), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_109), .Y(n_736) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_110), .B(n_446), .Y(n_725) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g445 ( .A(n_111), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_112), .B(n_446), .C(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_119), .B1(n_443), .B2(n_447), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_118), .A2(n_443), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_119), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_119), .Y(n_732) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_412), .Y(n_119) );
NOR3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_305), .C(n_378), .Y(n_120) );
OAI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_190), .B(n_237), .C(n_289), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_158), .Y(n_123) );
AND2x2_ASAP7_75t_L g253 ( .A(n_124), .B(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g272 ( .A(n_124), .Y(n_272) );
INVx2_ASAP7_75t_L g287 ( .A(n_124), .Y(n_287) );
INVx1_ASAP7_75t_L g317 ( .A(n_124), .Y(n_317) );
AND2x2_ASAP7_75t_L g367 ( .A(n_124), .B(n_288), .Y(n_367) );
AOI32xp33_ASAP7_75t_L g394 ( .A1(n_124), .A2(n_322), .A3(n_395), .B1(n_397), .B2(n_398), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_124), .B(n_243), .Y(n_400) );
AND2x2_ASAP7_75t_L g427 ( .A(n_124), .B(n_270), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_124), .B(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_154), .Y(n_124) );
AOI21xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_134), .B(n_147), .Y(n_125) );
BUFx2_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_128), .B(n_132), .Y(n_195) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g461 ( .A(n_129), .Y(n_461) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g202 ( .A(n_130), .Y(n_202) );
INVx1_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx3_ASAP7_75t_L g141 ( .A(n_131), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_131), .Y(n_143) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
INVx4_ASAP7_75t_SL g188 ( .A(n_132), .Y(n_188) );
BUFx3_ASAP7_75t_L g463 ( .A(n_132), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_132), .A2(n_470), .B(n_473), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_132), .A2(n_480), .B(n_484), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_132), .A2(n_501), .B(n_504), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_132), .A2(n_510), .B(n_514), .Y(n_509) );
INVx5_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx3_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
INVx1_ASAP7_75t_L g494 ( .A(n_136), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_142), .B(n_144), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_140), .A2(n_198), .B(n_199), .C(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_140), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_140), .A2(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g476 ( .A(n_140), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_SL g501 ( .A1(n_140), .A2(n_216), .B(n_502), .C(n_503), .Y(n_501) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_141), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_141), .B(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g528 ( .A1(n_141), .A2(n_168), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g513 ( .A(n_143), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_144), .A2(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
INVx1_ASAP7_75t_L g261 ( .A(n_147), .Y(n_261) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_147), .A2(n_454), .B(n_464), .Y(n_453) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_147), .A2(n_479), .B(n_487), .Y(n_478) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_148), .A2(n_193), .B(n_203), .Y(n_192) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_148), .A2(n_220), .B(n_227), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_148), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_150), .B(n_151), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_SL g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx3_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
AO21x1_ASAP7_75t_L g539 ( .A1(n_156), .A2(n_540), .B(n_543), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_156), .B(n_463), .C(n_540), .Y(n_564) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_157), .A2(n_230), .B(n_236), .Y(n_229) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_157), .A2(n_469), .B(n_477), .Y(n_468) );
AND2x2_ASAP7_75t_L g316 ( .A(n_158), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g338 ( .A(n_158), .Y(n_338) );
AND2x2_ASAP7_75t_L g423 ( .A(n_158), .B(n_253), .Y(n_423) );
AND2x2_ASAP7_75t_L g426 ( .A(n_158), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_175), .Y(n_158) );
INVx2_ASAP7_75t_L g245 ( .A(n_159), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_159), .B(n_270), .Y(n_276) );
AND2x2_ASAP7_75t_L g286 ( .A(n_159), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g322 ( .A(n_159), .Y(n_322) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_172), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_161), .A2(n_177), .B(n_189), .Y(n_176) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_161), .A2(n_500), .B(n_507), .Y(n_499) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_161), .A2(n_509), .B(n_517), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_171), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_169), .Y(n_164) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g213 ( .A(n_168), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_168), .A2(n_476), .B1(n_493), .B2(n_495), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_168), .A2(n_476), .B1(n_541), .B2(n_542), .Y(n_540) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g216 ( .A(n_170), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_174), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_174), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g264 ( .A(n_175), .B(n_245), .Y(n_264) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
AND2x2_ASAP7_75t_L g288 ( .A(n_176), .B(n_270), .Y(n_288) );
AND2x2_ASAP7_75t_L g357 ( .A(n_176), .B(n_254), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_188), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_181), .A2(n_188), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_181), .A2(n_188), .B(n_232), .C(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_183), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g483 ( .A(n_183), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_183), .A2(n_505), .B(n_506), .Y(n_504) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g222 ( .A1(n_184), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_222) );
INVx2_ASAP7_75t_L g224 ( .A(n_184), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_188), .A2(n_195), .B1(n_221), .B2(n_226), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_205), .Y(n_190) );
OR2x2_ASAP7_75t_L g251 ( .A(n_191), .B(n_219), .Y(n_251) );
INVx1_ASAP7_75t_L g330 ( .A(n_191), .Y(n_330) );
AND2x2_ASAP7_75t_L g344 ( .A(n_191), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_191), .B(n_218), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_191), .B(n_342), .Y(n_396) );
AND2x2_ASAP7_75t_L g404 ( .A(n_191), .B(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g241 ( .A(n_192), .Y(n_241) );
AND2x2_ASAP7_75t_L g311 ( .A(n_192), .B(n_219), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_195), .A2(n_256), .B(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_200), .A2(n_481), .B(n_482), .C(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_205), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g438 ( .A(n_205), .Y(n_438) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_218), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_206), .B(n_282), .Y(n_304) );
OR2x2_ASAP7_75t_L g333 ( .A(n_206), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g365 ( .A(n_206), .B(n_345), .Y(n_365) );
INVx1_ASAP7_75t_SL g385 ( .A(n_206), .Y(n_385) );
AND2x2_ASAP7_75t_L g389 ( .A(n_206), .B(n_250), .Y(n_389) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_SL g242 ( .A(n_207), .B(n_218), .Y(n_242) );
AND2x2_ASAP7_75t_L g249 ( .A(n_207), .B(n_229), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_207), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g292 ( .A(n_207), .B(n_274), .Y(n_292) );
INVx1_ASAP7_75t_SL g299 ( .A(n_207), .Y(n_299) );
BUFx2_ASAP7_75t_L g310 ( .A(n_207), .Y(n_310) );
AND2x2_ASAP7_75t_L g326 ( .A(n_207), .B(n_241), .Y(n_326) );
AND2x2_ASAP7_75t_L g341 ( .A(n_207), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g405 ( .A(n_207), .B(n_219), .Y(n_405) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_217), .Y(n_207) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_213), .A2(n_459), .B(n_460), .C(n_462), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_213), .A2(n_515), .B(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_218), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g329 ( .A(n_218), .B(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_218), .A2(n_347), .B1(n_350), .B2(n_353), .C(n_358), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_218), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
INVx3_ASAP7_75t_L g274 ( .A(n_219), .Y(n_274) );
BUFx2_ASAP7_75t_L g284 ( .A(n_229), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_229), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g315 ( .A(n_229), .Y(n_315) );
OR2x2_ASAP7_75t_L g334 ( .A(n_229), .B(n_274), .Y(n_334) );
INVx3_ASAP7_75t_L g342 ( .A(n_229), .Y(n_342) );
AND2x2_ASAP7_75t_L g345 ( .A(n_229), .B(n_274), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_243), .B1(n_247), .B2(n_252), .C(n_265), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_240), .B(n_314), .Y(n_439) );
OR2x2_ASAP7_75t_L g442 ( .A(n_240), .B(n_273), .Y(n_442) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OAI221xp5_ASAP7_75t_SL g265 ( .A1(n_241), .A2(n_266), .B1(n_273), .B2(n_275), .C(n_278), .Y(n_265) );
AND2x2_ASAP7_75t_L g282 ( .A(n_241), .B(n_274), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_241), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_241), .B(n_298), .Y(n_297) );
NAND2x1_ASAP7_75t_L g340 ( .A(n_241), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g392 ( .A(n_241), .B(n_334), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_243), .A2(n_352), .B1(n_381), .B2(n_383), .Y(n_380) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI322xp5_ASAP7_75t_L g289 ( .A1(n_244), .A2(n_253), .A3(n_290), .B1(n_293), .B2(n_296), .C1(n_300), .C2(n_303), .Y(n_289) );
OR2x2_ASAP7_75t_L g301 ( .A(n_244), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_245), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g280 ( .A(n_245), .B(n_254), .Y(n_280) );
INVx1_ASAP7_75t_L g295 ( .A(n_245), .Y(n_295) );
AND2x2_ASAP7_75t_L g361 ( .A(n_245), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g271 ( .A(n_246), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g362 ( .A(n_246), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_246), .B(n_270), .Y(n_436) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_250), .B(n_385), .Y(n_384) );
INVx3_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g336 ( .A(n_251), .B(n_283), .Y(n_336) );
OR2x2_ASAP7_75t_L g433 ( .A(n_251), .B(n_284), .Y(n_433) );
INVx1_ASAP7_75t_L g414 ( .A(n_252), .Y(n_414) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_264), .Y(n_252) );
INVx4_ASAP7_75t_L g302 ( .A(n_253), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_253), .B(n_321), .Y(n_327) );
INVx2_ASAP7_75t_L g270 ( .A(n_254), .Y(n_270) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_261), .B(n_262), .Y(n_254) );
INVx1_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_264), .B(n_324), .Y(n_393) );
AOI21xp33_ASAP7_75t_L g339 ( .A1(n_266), .A2(n_340), .B(n_343), .Y(n_339) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g324 ( .A(n_270), .Y(n_324) );
INVx1_ASAP7_75t_L g351 ( .A(n_270), .Y(n_351) );
INVx1_ASAP7_75t_L g277 ( .A(n_271), .Y(n_277) );
AND2x2_ASAP7_75t_L g279 ( .A(n_271), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g375 ( .A(n_272), .B(n_361), .Y(n_375) );
AND2x2_ASAP7_75t_L g397 ( .A(n_272), .B(n_357), .Y(n_397) );
BUFx2_ASAP7_75t_L g349 ( .A(n_274), .Y(n_349) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AOI32xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_281), .A3(n_282), .B1(n_283), .B2(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g359 ( .A(n_279), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_279), .A2(n_407), .B1(n_408), .B2(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_282), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_282), .B(n_341), .Y(n_382) );
AND2x2_ASAP7_75t_L g429 ( .A(n_282), .B(n_314), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_283), .B(n_330), .Y(n_377) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g430 ( .A(n_285), .Y(n_430) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g355 ( .A(n_286), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_288), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g402 ( .A(n_288), .B(n_322), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_288), .B(n_317), .Y(n_409) );
INVx1_ASAP7_75t_SL g391 ( .A(n_290), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_291), .B(n_342), .Y(n_369) );
NOR4xp25_ASAP7_75t_L g415 ( .A(n_291), .B(n_314), .C(n_416), .D(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_292), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_L g372 ( .A(n_295), .Y(n_372) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_298), .A2(n_389), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g314 ( .A(n_299), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND4xp25_ASAP7_75t_SL g305 ( .A(n_306), .B(n_331), .C(n_346), .D(n_366), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_312), .B(n_316), .C(n_318), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g398 ( .A(n_311), .B(n_341), .Y(n_398) );
AND2x2_ASAP7_75t_L g407 ( .A(n_311), .B(n_385), .Y(n_407) );
INVx3_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_314), .B(n_349), .Y(n_411) );
AND2x2_ASAP7_75t_L g323 ( .A(n_317), .B(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_325), .B1(n_327), .B2(n_328), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
AND2x2_ASAP7_75t_L g421 ( .A(n_321), .B(n_367), .Y(n_421) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_323), .B(n_372), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_324), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_337), .C(n_339), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_332), .A2(n_367), .B1(n_368), .B2(n_370), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_340), .A2(n_425), .B1(n_428), .B2(n_430), .C(n_431), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_341), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_349), .B(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g379 ( .A(n_351), .Y(n_379) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_354), .A2(n_374), .B1(n_376), .B2(n_377), .Y(n_373) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B(n_364), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_363), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_374), .A2(n_400), .B1(n_438), .B2(n_439), .C(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_380), .B(n_386), .C(n_406), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_390), .C(n_399), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_393), .C(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g418 ( .A(n_396), .Y(n_418) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_397), .A2(n_423), .B(n_441), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_403), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g432 ( .A1(n_409), .A2(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_424), .C(n_437), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_420), .C(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx14_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g728 ( .A(n_447), .Y(n_728) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR3x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_650), .C(n_699), .Y(n_448) );
NAND5xp2_ASAP7_75t_L g449 ( .A(n_450), .B(n_565), .C(n_593), .D(n_623), .E(n_637), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_488), .B1(n_518), .B2(n_523), .C(n_532), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_465), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_452), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g545 ( .A(n_453), .Y(n_545) );
AND2x2_ASAP7_75t_L g553 ( .A(n_453), .B(n_468), .Y(n_553) );
AND2x2_ASAP7_75t_L g576 ( .A(n_453), .B(n_467), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_453), .B(n_478), .Y(n_591) );
OR2x2_ASAP7_75t_L g600 ( .A(n_453), .B(n_539), .Y(n_600) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_453), .Y(n_603) );
AND2x2_ASAP7_75t_L g711 ( .A(n_453), .B(n_539), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B(n_463), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_460), .A2(n_476), .B(n_485), .C(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_465), .B(n_603), .Y(n_659) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
OAI311xp33_ASAP7_75t_L g601 ( .A1(n_466), .A2(n_602), .A3(n_603), .B1(n_604), .C1(n_619), .Y(n_601) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_478), .Y(n_466) );
AND2x2_ASAP7_75t_L g562 ( .A(n_467), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g569 ( .A(n_467), .Y(n_569) );
AND2x2_ASAP7_75t_L g690 ( .A(n_467), .B(n_522), .Y(n_690) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_468), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g546 ( .A(n_468), .B(n_478), .Y(n_546) );
AND2x2_ASAP7_75t_L g598 ( .A(n_468), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g612 ( .A(n_468), .B(n_545), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_476), .Y(n_473) );
INVx2_ASAP7_75t_L g522 ( .A(n_478), .Y(n_522) );
AND2x2_ASAP7_75t_L g561 ( .A(n_478), .B(n_545), .Y(n_561) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
OR2x2_ASAP7_75t_L g656 ( .A(n_489), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_489), .B(n_662), .Y(n_673) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_490), .B(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
AND2x2_ASAP7_75t_L g597 ( .A(n_491), .B(n_527), .Y(n_597) );
AND2x2_ASAP7_75t_L g608 ( .A(n_491), .B(n_508), .Y(n_608) );
AND2x2_ASAP7_75t_L g617 ( .A(n_491), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_496), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_496), .B(n_558), .Y(n_602) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g589 ( .A(n_497), .B(n_548), .Y(n_589) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
INVx2_ASAP7_75t_L g525 ( .A(n_498), .Y(n_525) );
AND2x2_ASAP7_75t_L g616 ( .A(n_498), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g535 ( .A(n_499), .Y(n_535) );
OR2x2_ASAP7_75t_L g633 ( .A(n_499), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_499), .Y(n_696) );
AND2x2_ASAP7_75t_L g536 ( .A(n_508), .B(n_531), .Y(n_536) );
INVx1_ASAP7_75t_L g556 ( .A(n_508), .Y(n_556) );
AND2x2_ASAP7_75t_L g577 ( .A(n_508), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g618 ( .A(n_508), .Y(n_618) );
INVx1_ASAP7_75t_L g634 ( .A(n_508), .Y(n_634) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_508), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_513), .Y(n_510) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_520), .B(n_622), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_520), .A2(n_607), .B1(n_656), .B2(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
OAI211xp5_ASAP7_75t_SL g699 ( .A1(n_521), .A2(n_700), .B(n_702), .C(n_720), .Y(n_699) );
INVx2_ASAP7_75t_L g552 ( .A(n_522), .Y(n_552) );
AND2x2_ASAP7_75t_L g610 ( .A(n_522), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g621 ( .A(n_522), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_523), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AND2x2_ASAP7_75t_L g594 ( .A(n_524), .B(n_558), .Y(n_594) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g626 ( .A(n_525), .B(n_617), .Y(n_626) );
AND2x2_ASAP7_75t_L g645 ( .A(n_525), .B(n_559), .Y(n_645) );
AND2x4_ASAP7_75t_L g581 ( .A(n_526), .B(n_555), .Y(n_581) );
AND2x2_ASAP7_75t_L g719 ( .A(n_526), .B(n_695), .Y(n_719) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_527), .Y(n_548) );
INVx1_ASAP7_75t_L g559 ( .A(n_527), .Y(n_559) );
INVx1_ASAP7_75t_L g658 ( .A(n_527), .Y(n_658) );
OR2x2_ASAP7_75t_L g549 ( .A(n_531), .B(n_535), .Y(n_549) );
AND2x2_ASAP7_75t_L g558 ( .A(n_531), .B(n_559), .Y(n_558) );
NOR2xp67_ASAP7_75t_L g578 ( .A(n_531), .B(n_579), .Y(n_578) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_537), .B1(n_547), .B2(n_550), .C(n_554), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_534), .A2(n_555), .B(n_557), .C(n_560), .Y(n_554) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g579 ( .A(n_535), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_535), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_535), .B(n_556), .Y(n_662) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_535), .Y(n_669) );
AND2x2_ASAP7_75t_L g587 ( .A(n_536), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g624 ( .A(n_536), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_546), .Y(n_537) );
INVx2_ASAP7_75t_L g615 ( .A(n_538), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_538), .A2(n_548), .B1(n_665), .B2(n_667), .C1(n_668), .C2(n_670), .Y(n_664) );
AND2x2_ASAP7_75t_L g721 ( .A(n_538), .B(n_690), .Y(n_721) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
INVx1_ASAP7_75t_L g611 ( .A(n_539), .Y(n_611) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g563 ( .A(n_544), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g649 ( .A(n_546), .B(n_583), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_547), .A2(n_661), .B(n_663), .Y(n_660) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g588 ( .A(n_548), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_548), .B(n_555), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_548), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx3_ASAP7_75t_L g614 ( .A(n_552), .Y(n_614) );
OR2x2_ASAP7_75t_L g666 ( .A(n_552), .B(n_588), .Y(n_666) );
AND2x2_ASAP7_75t_L g582 ( .A(n_553), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g620 ( .A(n_553), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_553), .B(n_614), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_553), .B(n_610), .Y(n_636) );
AND2x2_ASAP7_75t_L g640 ( .A(n_553), .B(n_622), .Y(n_640) );
INVxp67_ASAP7_75t_L g572 ( .A(n_555), .Y(n_572) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_557), .A2(n_630), .B1(n_635), .B2(n_636), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_557), .B(n_662), .Y(n_692) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g678 ( .A(n_558), .B(n_669), .Y(n_678) );
AND2x2_ASAP7_75t_L g707 ( .A(n_558), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_558), .B(n_662), .Y(n_712) );
INVx1_ASAP7_75t_L g625 ( .A(n_559), .Y(n_625) );
BUFx2_ASAP7_75t_L g631 ( .A(n_559), .Y(n_631) );
INVx1_ASAP7_75t_L g716 ( .A(n_560), .Y(n_716) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND2x1p5_ASAP7_75t_L g567 ( .A(n_561), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g592 ( .A(n_562), .Y(n_592) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_563), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_563), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g584 ( .A(n_563), .Y(n_584) );
INVx3_ASAP7_75t_L g622 ( .A(n_563), .Y(n_622) );
OR2x2_ASAP7_75t_L g688 ( .A(n_563), .B(n_689), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_570), .B(n_573), .C(n_585), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_566), .A2(n_703), .B1(n_710), .B2(n_712), .C(n_713), .Y(n_702) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_574), .B(n_580), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_576), .B(n_614), .Y(n_628) );
AND2x2_ASAP7_75t_L g670 ( .A(n_576), .B(n_610), .Y(n_670) );
INVx1_ASAP7_75t_SL g683 ( .A(n_577), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_577), .B(n_631), .Y(n_686) );
INVx1_ASAP7_75t_L g704 ( .A(n_578), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_582), .A2(n_672), .B1(n_674), .B2(n_678), .C(n_679), .Y(n_671) );
AND2x2_ASAP7_75t_L g698 ( .A(n_583), .B(n_690), .Y(n_698) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g682 ( .A(n_584), .Y(n_682) );
AOI21xp33_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_589), .B(n_590), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g653 ( .A(n_588), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g639 ( .A(n_589), .Y(n_639) );
INVx1_ASAP7_75t_L g667 ( .A(n_590), .Y(n_667) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_598), .C(n_601), .Y(n_593) );
OAI31xp33_ASAP7_75t_L g720 ( .A1(n_594), .A2(n_632), .A3(n_719), .B(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g694 ( .A(n_597), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g715 ( .A(n_597), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_599), .B(n_614), .Y(n_642) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g717 ( .A(n_600), .B(n_614), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_609), .B1(n_613), .B2(n_616), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_608), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g644 ( .A(n_608), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_608), .B(n_631), .Y(n_647) );
AND2x2_ASAP7_75t_L g701 ( .A(n_608), .B(n_696), .Y(n_701) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g676 ( .A(n_612), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OAI32xp33_ASAP7_75t_L g679 ( .A1(n_614), .A2(n_648), .A3(n_680), .B1(n_682), .B2(n_683), .Y(n_679) );
INVx1_ASAP7_75t_L g654 ( .A(n_617), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_617), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g677 ( .A(n_621), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_627), .C(n_629), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_625), .B(n_662), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_626), .A2(n_638), .B1(n_639), .B2(n_640), .C(n_641), .Y(n_637) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_636), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_646), .B2(n_648), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND4xp25_ASAP7_75t_SL g703 ( .A(n_646), .B(n_704), .C(n_705), .D(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
NAND4xp25_ASAP7_75t_SL g650 ( .A(n_651), .B(n_664), .C(n_671), .D(n_684), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B(n_659), .C(n_660), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g681 ( .A(n_657), .Y(n_681) );
INVx2_ASAP7_75t_L g705 ( .A(n_662), .Y(n_705) );
OR2x2_ASAP7_75t_L g714 ( .A(n_669), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_691), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g710 ( .A(n_690), .B(n_711), .Y(n_710) );
AOI21xp33_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_693), .B(n_697), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
CKINVDCx16_ASAP7_75t_R g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g748 ( .A(n_739), .Y(n_748) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx14_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule