module fake_netlist_5_2367_n_1243 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_10, n_24, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1243);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_10;
input n_24;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1243;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_546;
wire n_731;
wire n_371;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_582;
wire n_512;
wire n_322;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1123;
wire n_1047;
wire n_634;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_922;
wire n_816;
wire n_591;
wire n_631;
wire n_479;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_384;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1113;
wire n_1226;
wire n_722;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_846;
wire n_465;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_215),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_201),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_25),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_206),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_52),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_246),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_217),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_247),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_109),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_150),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_66),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_216),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_12),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_53),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_60),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_296),
.Y(n_344)
);

BUFx2_ASAP7_75t_SL g345 ( 
.A(n_197),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_240),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_208),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_162),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_130),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_34),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_144),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_200),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_170),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_220),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_80),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_18),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_222),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_180),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_279),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_272),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_218),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_183),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_149),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_17),
.B(n_51),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_174),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_122),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_54),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_230),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_7),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_108),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_317),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_195),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_108),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_214),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_184),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_292),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_312),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_226),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_137),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_54),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_155),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_104),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_38),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_251),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_280),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_127),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_287),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_125),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_207),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_139),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_3),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_16),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_14),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_104),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_223),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_244),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_132),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_284),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_81),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_266),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_229),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_45),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_293),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_124),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_213),
.Y(n_413)
);

BUFx10_ASAP7_75t_L g414 ( 
.A(n_3),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_320),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_138),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_120),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_51),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_306),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_237),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_25),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_189),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_188),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_56),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_55),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_187),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_182),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_43),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_131),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_40),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_211),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_277),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_304),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_178),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_262),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_205),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_56),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_135),
.B(n_298),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_286),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_4),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_110),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_129),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_126),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_299),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_142),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_45),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_318),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_245),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_267),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_303),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_128),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_241),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_18),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_305),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_212),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_113),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_291),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_136),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_193),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_231),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_121),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_73),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_152),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_209),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_254),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_36),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_238),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_9),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_154),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_141),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_23),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_311),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_199),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_264),
.B(n_19),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_15),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_110),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_310),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_140),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_243),
.B(n_210),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_309),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_64),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_0),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_350),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_330),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_373),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_333),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_376),
.B(n_1),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_333),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_414),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_330),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_450),
.Y(n_495)
);

AOI22x1_ASAP7_75t_SL g496 ( 
.A1(n_425),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_430),
.A2(n_6),
.B1(n_2),
.B2(n_5),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

OAI22x1_ASAP7_75t_SL g499 ( 
.A1(n_425),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_378),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_395),
.B(n_422),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_123),
.Y(n_505)
);

AOI22x1_ASAP7_75t_SL g506 ( 
.A1(n_437),
.A2(n_466),
.B1(n_335),
.B2(n_339),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_468),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_350),
.B(n_8),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_441),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_331),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_337),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_340),
.Y(n_517)
);

CKINVDCx6p67_ASAP7_75t_R g518 ( 
.A(n_385),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_475),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_452),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_364),
.A2(n_9),
.B(n_10),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_437),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_364),
.B(n_10),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_452),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_408),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_472),
.B(n_11),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_341),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_472),
.B(n_13),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g530 ( 
.A1(n_365),
.A2(n_369),
.B(n_366),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_481),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_466),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_365),
.B(n_19),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_436),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_324),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_474),
.B(n_20),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_352),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_358),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_446),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_360),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_326),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_375),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_369),
.B(n_21),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_397),
.B(n_22),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_327),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_379),
.B(n_23),
.Y(n_546)
);

BUFx12f_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_417),
.B(n_24),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_363),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_332),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_336),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_486),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_488),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_525),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_329),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_536),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_518),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_500),
.B(n_477),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_483),
.B(n_536),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_505),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_483),
.B(n_338),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_525),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_491),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_511),
.A2(n_370),
.B(n_438),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_549),
.B(n_464),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_525),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_501),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_527),
.B(n_338),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_527),
.B(n_368),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_495),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_486),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_495),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_494),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_537),
.B(n_345),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_515),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_551),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_494),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_535),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_494),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_485),
.A2(n_534),
.B1(n_526),
.B2(n_511),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_549),
.B(n_464),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_SL g586 ( 
.A(n_490),
.B(n_368),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_532),
.A2(n_371),
.B1(n_380),
.B2(n_377),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_529),
.B(n_371),
.Y(n_588)
);

NOR2x1p5_ASAP7_75t_L g589 ( 
.A(n_492),
.B(n_462),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_547),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_545),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_559),
.Y(n_592)
);

INVx8_ASAP7_75t_L g593 ( 
.A(n_557),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_560),
.B(n_538),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_516),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_581),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_582),
.B(n_570),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_585),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_556),
.B(n_505),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_555),
.B(n_589),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_591),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_562),
.A2(n_517),
.B1(n_508),
.B2(n_353),
.Y(n_602)
);

BUFx12f_ASAP7_75t_L g603 ( 
.A(n_558),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_554),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_566),
.B(n_517),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_561),
.B(n_529),
.Y(n_607)
);

OAI21xp33_ASAP7_75t_L g608 ( 
.A1(n_583),
.A2(n_539),
.B(n_484),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_570),
.B(n_552),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_566),
.B(n_552),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_554),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_566),
.A2(n_530),
.B1(n_522),
.B2(n_524),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_570),
.B(n_528),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_553),
.B(n_540),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_578),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_565),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_563),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_567),
.A2(n_530),
.B(n_533),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_574),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_563),
.B(n_512),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_564),
.B(n_520),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_580),
.B(n_489),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_571),
.B(n_489),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_586),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_571),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_572),
.B(n_520),
.Y(n_627)
);

AO221x1_ASAP7_75t_L g628 ( 
.A1(n_587),
.A2(n_503),
.B1(n_502),
.B2(n_342),
.C(n_348),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_586),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_572),
.B(n_504),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_575),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_588),
.B(n_510),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_558),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_577),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_557),
.B(n_504),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_557),
.B(n_550),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_579),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_610),
.A2(n_618),
.B(n_612),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_594),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_592),
.A2(n_562),
.B1(n_548),
.B2(n_546),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_594),
.A2(n_561),
.B1(n_392),
.B2(n_457),
.Y(n_642)
);

AO32x1_ASAP7_75t_L g643 ( 
.A1(n_625),
.A2(n_349),
.A3(n_351),
.B1(n_347),
.B2(n_343),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_595),
.B(n_614),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_624),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_610),
.B(n_584),
.Y(n_646)
);

AO22x1_ASAP7_75t_L g647 ( 
.A1(n_606),
.A2(n_544),
.B1(n_543),
.B2(n_399),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_608),
.A2(n_543),
.B(n_544),
.C(n_546),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_596),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_612),
.B(n_627),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_638),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_629),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_613),
.B(n_577),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_598),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_601),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_629),
.B(n_497),
.C(n_590),
.Y(n_656)
);

A2O1A1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_630),
.A2(n_479),
.B(n_354),
.C(n_359),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_627),
.B(n_577),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_622),
.Y(n_660)
);

CKINVDCx8_ASAP7_75t_R g661 ( 
.A(n_634),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_623),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_630),
.B(n_355),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_607),
.A2(n_633),
.B(n_600),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_628),
.A2(n_372),
.B1(n_384),
.B2(n_382),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_636),
.A2(n_388),
.B(n_386),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_602),
.B(n_577),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_636),
.A2(n_394),
.B(n_391),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_605),
.B(n_523),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_635),
.A2(n_356),
.B1(n_380),
.B2(n_377),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_616),
.B(n_398),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_620),
.A2(n_479),
.B(n_409),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_631),
.B(n_632),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_603),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_637),
.B(n_403),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_626),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_617),
.B(n_420),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_621),
.A2(n_426),
.B(n_429),
.C(n_423),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_605),
.B(n_523),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_609),
.A2(n_432),
.B(n_431),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_621),
.A2(n_442),
.B(n_439),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_597),
.B(n_619),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_593),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_593),
.A2(n_448),
.B(n_445),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_626),
.Y(n_687)
);

OA22x2_ASAP7_75t_L g688 ( 
.A1(n_628),
.A2(n_539),
.B1(n_471),
.B2(n_325),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_592),
.B(n_403),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_592),
.B(n_482),
.C(n_569),
.Y(n_690)
);

OAI321xp33_ASAP7_75t_L g691 ( 
.A1(n_592),
.A2(n_531),
.A3(n_521),
.B1(n_458),
.B2(n_455),
.C(n_459),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_622),
.Y(n_692)
);

INVx3_ASAP7_75t_SL g693 ( 
.A(n_634),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_592),
.B(n_463),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_595),
.B(n_569),
.Y(n_695)
);

AOI21xp33_ASAP7_75t_L g696 ( 
.A1(n_592),
.A2(n_415),
.B(n_383),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_599),
.A2(n_470),
.B(n_467),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_610),
.A2(n_323),
.B(n_322),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_592),
.A2(n_434),
.B1(n_499),
.B2(n_334),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_595),
.B(n_487),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_626),
.Y(n_702)
);

AOI22x1_ASAP7_75t_L g703 ( 
.A1(n_618),
.A2(n_344),
.B1(n_346),
.B2(n_328),
.Y(n_703)
);

INVx11_ASAP7_75t_L g704 ( 
.A(n_603),
.Y(n_704)
);

BUFx4f_ASAP7_75t_L g705 ( 
.A(n_593),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_633),
.B(n_493),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_SL g707 ( 
.A(n_607),
.B(n_357),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_592),
.B(n_434),
.Y(n_708)
);

O2A1O1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_592),
.A2(n_509),
.B(n_519),
.C(n_498),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_592),
.A2(n_362),
.B1(n_367),
.B2(n_361),
.Y(n_710)
);

OA22x2_ASAP7_75t_L g711 ( 
.A1(n_628),
.A2(n_424),
.B1(n_428),
.B2(n_421),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_592),
.B(n_374),
.Y(n_712)
);

BUFx8_ASAP7_75t_L g713 ( 
.A(n_603),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_596),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_605),
.B(n_509),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_592),
.A2(n_513),
.B(n_514),
.C(n_507),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_592),
.B(n_440),
.Y(n_717)
);

O2A1O1Ixp5_ASAP7_75t_L g718 ( 
.A1(n_610),
.A2(n_513),
.B(n_514),
.C(n_507),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_592),
.B(n_381),
.Y(n_719)
);

NOR4xp25_ASAP7_75t_L g720 ( 
.A(n_708),
.B(n_496),
.C(n_506),
.D(n_461),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_718),
.A2(n_396),
.B(n_393),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_640),
.A2(n_405),
.B1(n_406),
.B2(n_404),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_650),
.A2(n_412),
.B1(n_413),
.B2(n_411),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_649),
.Y(n_724)
);

OAI22x1_ASAP7_75t_L g725 ( 
.A1(n_699),
.A2(n_419),
.B1(n_427),
.B2(n_416),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_717),
.A2(n_435),
.B1(n_443),
.B2(n_433),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_712),
.B(n_444),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_644),
.Y(n_728)
);

OA21x2_ASAP7_75t_L g729 ( 
.A1(n_639),
.A2(n_449),
.B(n_447),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_654),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_646),
.A2(n_454),
.B(n_451),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_655),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_666),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_700),
.B(n_662),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_689),
.B(n_460),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_694),
.A2(n_469),
.B1(n_473),
.B2(n_465),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_719),
.B(n_478),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_695),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_714),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_687),
.Y(n_740)
);

A2O1A1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_696),
.A2(n_480),
.B(n_27),
.C(n_24),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_675),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_645),
.B(n_26),
.Y(n_743)
);

CKINVDCx11_ASAP7_75t_R g744 ( 
.A(n_661),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_658),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_690),
.B(n_26),
.C(n_27),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_28),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_641),
.B(n_642),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_641),
.B(n_28),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_685),
.B(n_133),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_647),
.B(n_29),
.Y(n_751)
);

AOI21xp33_ASAP7_75t_L g752 ( 
.A1(n_698),
.A2(n_29),
.B(n_30),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_687),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_665),
.B(n_134),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_660),
.B(n_30),
.Y(n_755)
);

AND3x4_ASAP7_75t_L g756 ( 
.A(n_656),
.B(n_31),
.C(n_32),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_687),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_668),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_758)
);

AOI21xp33_ASAP7_75t_L g759 ( 
.A1(n_659),
.A2(n_33),
.B(n_35),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_706),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_652),
.A2(n_145),
.B1(n_146),
.B2(n_143),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_648),
.A2(n_148),
.B(n_147),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_702),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_651),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_664),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_697),
.A2(n_153),
.B(n_151),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_670),
.B(n_37),
.Y(n_767)
);

NOR2x1_ASAP7_75t_SL g768 ( 
.A(n_685),
.B(n_156),
.Y(n_768)
);

BUFx8_ASAP7_75t_L g769 ( 
.A(n_702),
.Y(n_769)
);

OAI21x1_ASAP7_75t_SL g770 ( 
.A1(n_674),
.A2(n_158),
.B(n_157),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_716),
.A2(n_160),
.B(n_159),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_701),
.Y(n_772)
);

OAI21xp33_ASAP7_75t_L g773 ( 
.A1(n_677),
.A2(n_38),
.B(n_39),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_693),
.Y(n_774)
);

OAI21x1_ASAP7_75t_SL g775 ( 
.A1(n_686),
.A2(n_163),
.B(n_161),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_669),
.A2(n_692),
.B1(n_684),
.B2(n_710),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_703),
.A2(n_165),
.B(n_164),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_702),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_678),
.Y(n_779)
);

AO21x1_ASAP7_75t_L g780 ( 
.A1(n_683),
.A2(n_41),
.B(n_42),
.Y(n_780)
);

AOI211x1_ASAP7_75t_L g781 ( 
.A1(n_682),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_709),
.A2(n_167),
.B(n_166),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_679),
.A2(n_169),
.B(n_168),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_667),
.A2(n_672),
.B1(n_705),
.B2(n_673),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_691),
.A2(n_172),
.B(n_171),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_705),
.A2(n_175),
.B1(n_176),
.B2(n_173),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_713),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_653),
.B(n_177),
.Y(n_788)
);

AO31x2_ASAP7_75t_L g789 ( 
.A1(n_680),
.A2(n_47),
.A3(n_44),
.B(n_46),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_711),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_671),
.B(n_47),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_681),
.B(n_48),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_715),
.B(n_179),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_688),
.A2(n_185),
.B1(n_186),
.B2(n_181),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_699),
.B(n_49),
.Y(n_795)
);

AO21x1_ASAP7_75t_L g796 ( 
.A1(n_643),
.A2(n_49),
.B(n_50),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_676),
.B(n_190),
.Y(n_797)
);

AO31x2_ASAP7_75t_L g798 ( 
.A1(n_643),
.A2(n_55),
.A3(n_52),
.B(n_53),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_707),
.B(n_57),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_643),
.B(n_57),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_713),
.B(n_58),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_704),
.A2(n_192),
.B(n_191),
.Y(n_802)
);

AOI21xp33_ASAP7_75t_L g803 ( 
.A1(n_708),
.A2(n_58),
.B(n_59),
.Y(n_803)
);

OA22x2_ASAP7_75t_L g804 ( 
.A1(n_699),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_644),
.B(n_61),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_640),
.B(n_62),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_640),
.B(n_62),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_640),
.A2(n_196),
.B1(n_198),
.B2(n_194),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_640),
.B(n_63),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_644),
.B(n_65),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_708),
.B(n_66),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_693),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_700),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_689),
.B(n_67),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_708),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_692),
.B(n_202),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_685),
.B(n_203),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_644),
.B(n_68),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_644),
.B(n_69),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_700),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_685),
.B(n_204),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_644),
.B(n_70),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_640),
.B(n_70),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_708),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_640),
.B(n_71),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_640),
.B(n_72),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_SL g827 ( 
.A(n_640),
.B(n_74),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_640),
.B(n_74),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_689),
.B(n_75),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_687),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_640),
.B(n_75),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_644),
.Y(n_832)
);

AO31x2_ASAP7_75t_L g833 ( 
.A1(n_650),
.A2(n_76),
.A3(n_77),
.B(n_78),
.Y(n_833)
);

AO31x2_ASAP7_75t_L g834 ( 
.A1(n_650),
.A2(n_76),
.A3(n_77),
.B(n_78),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_640),
.B(n_79),
.Y(n_835)
);

BUFx5_ASAP7_75t_L g836 ( 
.A(n_649),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_693),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_708),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_640),
.A2(n_239),
.B1(n_314),
.B2(n_313),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_649),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_649),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_650),
.A2(n_82),
.A3(n_83),
.B(n_84),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_700),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_718),
.A2(n_221),
.B(n_219),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_644),
.B(n_82),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_734),
.B(n_83),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_728),
.B(n_84),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_724),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_778),
.B(n_224),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_811),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_748),
.A2(n_752),
.B1(n_749),
.B2(n_767),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_795),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_730),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_732),
.Y(n_854)
);

NAND2x1_ASAP7_75t_L g855 ( 
.A(n_740),
.B(n_225),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_739),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_733),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_762),
.A2(n_88),
.B(n_89),
.C(n_90),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_774),
.B(n_88),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_832),
.Y(n_860)
);

AO21x2_ASAP7_75t_L g861 ( 
.A1(n_844),
.A2(n_249),
.B(n_302),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_776),
.A2(n_248),
.B1(n_301),
.B2(n_300),
.Y(n_862)
);

OAI22xp33_ASAP7_75t_L g863 ( 
.A1(n_814),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_SL g864 ( 
.A1(n_754),
.A2(n_242),
.B(n_295),
.C(n_294),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_742),
.B(n_806),
.Y(n_865)
);

AOI221xp5_ASAP7_75t_L g866 ( 
.A1(n_803),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_769),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_759),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.C(n_96),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_742),
.A2(n_236),
.B1(n_289),
.B2(n_288),
.Y(n_869)
);

BUFx4_ASAP7_75t_SL g870 ( 
.A(n_837),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_727),
.A2(n_235),
.B(n_285),
.Y(n_871)
);

OAI21x1_ASAP7_75t_SL g872 ( 
.A1(n_768),
.A2(n_234),
.B(n_283),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_738),
.Y(n_873)
);

AOI21xp33_ASAP7_75t_L g874 ( 
.A1(n_735),
.A2(n_95),
.B(n_96),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_790),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_758),
.B(n_97),
.C(n_98),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_807),
.A2(n_233),
.B1(n_275),
.B2(n_274),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_840),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_809),
.B(n_97),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_782),
.A2(n_232),
.B(n_273),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_813),
.B(n_98),
.Y(n_881)
);

OAI21x1_ASAP7_75t_SL g882 ( 
.A1(n_768),
.A2(n_250),
.B(n_271),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_823),
.A2(n_826),
.B(n_825),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_SL g884 ( 
.A1(n_828),
.A2(n_835),
.B(n_831),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_745),
.Y(n_885)
);

AOI222xp33_ASAP7_75t_SL g886 ( 
.A1(n_756),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C1(n_102),
.C2(n_103),
.Y(n_886)
);

OAI21x1_ASAP7_75t_SL g887 ( 
.A1(n_770),
.A2(n_775),
.B(n_771),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_820),
.B(n_99),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_744),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_843),
.B(n_100),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_765),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_740),
.B(n_228),
.Y(n_892)
);

BUFx2_ASAP7_75t_SL g893 ( 
.A(n_753),
.Y(n_893)
);

BUFx8_ASAP7_75t_L g894 ( 
.A(n_787),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_760),
.B(n_805),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_755),
.B(n_101),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_777),
.A2(n_252),
.B(n_270),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_836),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_737),
.A2(n_227),
.B1(n_269),
.B2(n_268),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_812),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_836),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_769),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_773),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.C(n_106),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_753),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_753),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_731),
.A2(n_261),
.B1(n_260),
.B2(n_259),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_764),
.B(n_105),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_743),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_757),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_747),
.A2(n_258),
.B(n_257),
.Y(n_910)
);

OR2x6_ASAP7_75t_L g911 ( 
.A(n_763),
.B(n_106),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_763),
.B(n_256),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_757),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_779),
.A2(n_253),
.B1(n_111),
.B2(n_112),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_757),
.B(n_107),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_830),
.Y(n_916)
);

AOI22x1_ASAP7_75t_L g917 ( 
.A1(n_721),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_772),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_793),
.A2(n_114),
.B(n_115),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_816),
.B(n_115),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_810),
.Y(n_921)
);

INVx3_ASAP7_75t_SL g922 ( 
.A(n_791),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_788),
.B(n_116),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_SL g924 ( 
.A1(n_815),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_L g925 ( 
.A(n_784),
.B(n_121),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_827),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_SL g927 ( 
.A1(n_792),
.A2(n_829),
.B1(n_804),
.B2(n_791),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_818),
.B(n_845),
.Y(n_928)
);

BUFx2_ASAP7_75t_SL g929 ( 
.A(n_819),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_822),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_751),
.Y(n_931)
);

OAI222xp33_ASAP7_75t_L g932 ( 
.A1(n_794),
.A2(n_761),
.B1(n_723),
.B2(n_800),
.C1(n_786),
.C2(n_722),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_725),
.B(n_720),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_729),
.A2(n_766),
.B(n_785),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_726),
.B(n_736),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_746),
.B(n_799),
.Y(n_936)
);

AO21x2_ASAP7_75t_L g937 ( 
.A1(n_802),
.A2(n_783),
.B(n_839),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_750),
.A2(n_817),
.B(n_821),
.Y(n_938)
);

AO31x2_ASAP7_75t_L g939 ( 
.A1(n_780),
.A2(n_838),
.A3(n_824),
.B(n_741),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_808),
.A2(n_801),
.B(n_781),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_789),
.B(n_833),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_798),
.A2(n_797),
.B(n_833),
.Y(n_942)
);

AOI221xp5_ASAP7_75t_L g943 ( 
.A1(n_833),
.A2(n_708),
.B1(n_583),
.B2(n_689),
.C(n_811),
.Y(n_943)
);

CKINVDCx8_ASAP7_75t_R g944 ( 
.A(n_834),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_834),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_842),
.A2(n_650),
.B(n_640),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_842),
.B(n_778),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_753),
.Y(n_948)
);

OA21x2_ASAP7_75t_L g949 ( 
.A1(n_844),
.A2(n_639),
.B(n_762),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_728),
.B(n_689),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_811),
.A2(n_762),
.B(n_640),
.Y(n_951)
);

OA21x2_ASAP7_75t_L g952 ( 
.A1(n_844),
.A2(n_639),
.B(n_762),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_811),
.A2(n_708),
.B(n_640),
.C(n_717),
.Y(n_953)
);

AO31x2_ASAP7_75t_L g954 ( 
.A1(n_796),
.A2(n_610),
.A3(n_657),
.B(n_780),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_728),
.B(n_708),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_733),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_841),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_728),
.B(n_689),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_811),
.A2(n_708),
.B1(n_717),
.B2(n_640),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_724),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_724),
.Y(n_961)
);

OA21x2_ASAP7_75t_L g962 ( 
.A1(n_844),
.A2(n_639),
.B(n_762),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_724),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_728),
.B(n_708),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_811),
.A2(n_708),
.B1(n_748),
.B2(n_640),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_742),
.B(n_640),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_841),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_733),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_769),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_848),
.Y(n_970)
);

AOI21xp33_ASAP7_75t_SL g971 ( 
.A1(n_955),
.A2(n_964),
.B(n_922),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_913),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_857),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_860),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_948),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_900),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_853),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_898),
.B(n_901),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_854),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_856),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_856),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_950),
.B(n_958),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_895),
.B(n_846),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_956),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_SL g985 ( 
.A1(n_917),
.A2(n_876),
.B1(n_920),
.B2(n_925),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_878),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_873),
.B(n_968),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_875),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_961),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_921),
.B(n_847),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_948),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_963),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_885),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_969),
.Y(n_994)
);

OA21x2_ASAP7_75t_L g995 ( 
.A1(n_934),
.A2(n_942),
.B(n_946),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_891),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_960),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_957),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_904),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_867),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_967),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_966),
.B(n_928),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_918),
.Y(n_1003)
);

INVx8_ASAP7_75t_L g1004 ( 
.A(n_849),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_865),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_905),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_907),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_904),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_908),
.B(n_930),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_965),
.B(n_959),
.Y(n_1010)
);

INVx6_ASAP7_75t_L g1011 ( 
.A(n_894),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_903),
.A2(n_866),
.B1(n_868),
.B2(n_943),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_947),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_888),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_894),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_855),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_890),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_953),
.B(n_851),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_931),
.B(n_929),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_927),
.B(n_923),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_941),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_923),
.B(n_936),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_949),
.A2(n_962),
.B(n_952),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_945),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_909),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_916),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_896),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_883),
.B(n_884),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_870),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_879),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_936),
.B(n_915),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_949),
.A2(n_962),
.B(n_952),
.Y(n_1032)
);

AO21x1_ASAP7_75t_SL g1033 ( 
.A1(n_932),
.A2(n_862),
.B(n_850),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_915),
.B(n_902),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_889),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_951),
.A2(n_887),
.B(n_937),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_924),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_938),
.B(n_933),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_893),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_926),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_917),
.A2(n_852),
.B1(n_874),
.B2(n_863),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_940),
.A2(n_858),
.B(n_935),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_912),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_939),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_914),
.A2(n_906),
.B(n_919),
.C(n_910),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_911),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_911),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_881),
.B(n_859),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_939),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_939),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_859),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_944),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_886),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_872),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_882),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_877),
.A2(n_899),
.B1(n_869),
.B2(n_871),
.C(n_864),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_954),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_861),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_880),
.B(n_897),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_892),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_934),
.A2(n_942),
.B(n_946),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_892),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1005),
.B(n_979),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_972),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_982),
.B(n_1002),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_1027),
.B(n_987),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_984),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1030),
.B(n_983),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1031),
.B(n_990),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_974),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1022),
.B(n_1020),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_974),
.B(n_984),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_972),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1009),
.B(n_1019),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1010),
.B(n_1014),
.Y(n_1075)
);

INVx4_ASAP7_75t_R g1076 ( 
.A(n_976),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1010),
.B(n_1017),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1053),
.A2(n_1012),
.B1(n_1033),
.B2(n_1041),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_970),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1018),
.B(n_1007),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1006),
.B(n_998),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_973),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_988),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_971),
.B(n_1004),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_993),
.B(n_996),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_997),
.B(n_1025),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1048),
.B(n_1034),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1013),
.B(n_977),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_980),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1026),
.B(n_1001),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_981),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_986),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_989),
.B(n_992),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1024),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1028),
.B(n_1060),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1062),
.B(n_1038),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1062),
.B(n_976),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1052),
.B(n_1046),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1039),
.B(n_1035),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_985),
.B(n_1041),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_985),
.B(n_1012),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_1000),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1021),
.B(n_1049),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1037),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1044),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1000),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1053),
.B(n_1051),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1050),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1042),
.B(n_1057),
.Y(n_1113)
);

BUFx8_ASAP7_75t_L g1114 ( 
.A(n_1029),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1042),
.B(n_1057),
.Y(n_1115)
);

INVxp67_ASAP7_75t_R g1116 ( 
.A(n_1015),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_978),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1095),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1065),
.B(n_999),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1079),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1090),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1092),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1078),
.A2(n_1045),
.B1(n_1056),
.B2(n_994),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1097),
.B(n_1055),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1107),
.B(n_1036),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1080),
.B(n_999),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1093),
.Y(n_1127)
);

INVxp33_ASAP7_75t_L g1128 ( 
.A(n_1069),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1080),
.B(n_999),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1094),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1075),
.B(n_1023),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1113),
.B(n_1061),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1072),
.B(n_1066),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1113),
.B(n_995),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1115),
.B(n_1023),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1115),
.B(n_995),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1077),
.B(n_1032),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1063),
.B(n_1032),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1081),
.B(n_1059),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1068),
.B(n_1008),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1067),
.B(n_1054),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1070),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_1084),
.B(n_975),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1109),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1112),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1085),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1110),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1074),
.B(n_1008),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1089),
.B(n_1058),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1105),
.B(n_991),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_1064),
.B(n_1016),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1144),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1145),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1123),
.B(n_1104),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1133),
.B(n_1070),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1118),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1120),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1121),
.Y(n_1158)
);

OAI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1128),
.A2(n_1078),
.B(n_1096),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1122),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1127),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1147),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1128),
.B(n_1150),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1146),
.B(n_1103),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1124),
.B(n_1099),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1125),
.B(n_1132),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1124),
.B(n_1099),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1134),
.B(n_1136),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1142),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1139),
.B(n_1086),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1151),
.B(n_1117),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1152),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1166),
.B(n_1138),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1153),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1172),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1156),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1157),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_1165),
.B(n_1131),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1170),
.B(n_1130),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1162),
.Y(n_1181)
);

OAI33xp33_ASAP7_75t_L g1182 ( 
.A1(n_1155),
.A2(n_1141),
.A3(n_1140),
.B1(n_1119),
.B2(n_1108),
.B3(n_1148),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1166),
.B(n_1149),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1158),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1159),
.B(n_1015),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1154),
.B(n_1126),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1167),
.B(n_1135),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1160),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1165),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1169),
.B(n_1135),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1161),
.Y(n_1191)
);

AO21x1_ASAP7_75t_SL g1192 ( 
.A1(n_1180),
.A2(n_1137),
.B(n_1164),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1186),
.A2(n_1154),
.B(n_1111),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1173),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1186),
.B(n_1163),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1175),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1177),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1187),
.B(n_1163),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1187),
.B(n_1190),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1178),
.Y(n_1200)
);

NAND2x1_ASAP7_75t_L g1201 ( 
.A(n_1176),
.B(n_1076),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1185),
.A2(n_1045),
.B(n_1143),
.C(n_1073),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1179),
.A2(n_1129),
.B(n_1171),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1181),
.A2(n_1168),
.B1(n_1071),
.B2(n_1011),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1181),
.A2(n_1056),
.B(n_1172),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1184),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1194),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1195),
.B(n_1190),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1198),
.B(n_1203),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1199),
.B(n_1174),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1196),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1197),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1192),
.B(n_1174),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1193),
.A2(n_1182),
.B(n_1179),
.C(n_1100),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1214),
.B(n_1193),
.C(n_1202),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1209),
.B(n_1200),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1211),
.A2(n_1205),
.B1(n_1212),
.B2(n_1208),
.C(n_1207),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1213),
.A2(n_1204),
.B(n_1205),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1213),
.A2(n_1206),
.B1(n_1191),
.B2(n_1188),
.C(n_1083),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1216),
.B(n_1210),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1217),
.B(n_1210),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1215),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1218),
.B(n_1011),
.Y(n_1223)
);

NOR2x1_ASAP7_75t_L g1224 ( 
.A(n_1219),
.B(n_1201),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1217),
.B(n_1183),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1222),
.B(n_1101),
.C(n_1088),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1223),
.B(n_1064),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1221),
.B(n_1176),
.Y(n_1228)
);

AND4x2_ASAP7_75t_L g1229 ( 
.A(n_1228),
.B(n_1224),
.C(n_1011),
.D(n_1225),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1227),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1230),
.B(n_1226),
.Y(n_1231)
);

OA22x2_ASAP7_75t_L g1232 ( 
.A1(n_1231),
.A2(n_1229),
.B1(n_1220),
.B2(n_1176),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1232),
.A2(n_1179),
.B1(n_1114),
.B2(n_1073),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1232),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1234),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1233),
.A2(n_1082),
.B(n_1102),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1235),
.A2(n_1236),
.B(n_1189),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1235),
.A2(n_1116),
.B1(n_1114),
.B2(n_1110),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1237),
.B(n_1238),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1238),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1240),
.B(n_1239),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_SL g1242 ( 
.A(n_1241),
.B(n_1106),
.C(n_1098),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1242),
.A2(n_1087),
.B(n_1091),
.Y(n_1243)
);


endmodule