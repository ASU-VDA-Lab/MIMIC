module real_jpeg_4549_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_0),
.A2(n_50),
.B1(n_115),
.B2(n_252),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_0),
.A2(n_50),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_0),
.A2(n_50),
.B1(n_452),
.B2(n_454),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_134),
.B1(n_138),
.B2(n_141),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_1),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_141),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_1),
.A2(n_141),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_2),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_2),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_92),
.B1(n_95),
.B2(n_99),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_3),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_99),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_99),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_4),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_4),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_5),
.A2(n_51),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_5),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_5),
.A2(n_236),
.B1(n_259),
.B2(n_289),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_5),
.A2(n_259),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_5),
.A2(n_259),
.B1(n_390),
.B2(n_448),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_6),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_6),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_6),
.B(n_88),
.C(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_6),
.B(n_116),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_6),
.B(n_295),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_6),
.B(n_90),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_6),
.B(n_152),
.Y(n_357)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g420 ( 
.A(n_7),
.Y(n_420)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_8),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_9),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_9),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_9),
.A2(n_215),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_9),
.A2(n_215),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_9),
.A2(n_131),
.B1(n_180),
.B2(n_215),
.Y(n_359)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_12),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_13),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_13),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_13),
.A2(n_129),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_13),
.A2(n_129),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_13),
.A2(n_129),
.B1(n_399),
.B2(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_15),
.A2(n_33),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_15),
.A2(n_60),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_15),
.A2(n_60),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_15),
.A2(n_60),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_16),
.A2(n_249),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_16),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_16),
.A2(n_304),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_16),
.A2(n_304),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_16),
.A2(n_58),
.B1(n_304),
.B2(n_475),
.Y(n_474)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_18),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_521),
.B(n_523),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_220),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_219),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_163),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_24),
.B(n_163),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_142),
.B2(n_143),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_61),
.C(n_100),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_27),
.A2(n_144),
.B1(n_145),
.B2(n_162),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_27),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_28),
.A2(n_55),
.B1(n_57),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_28),
.A2(n_257),
.B(n_260),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_28),
.A2(n_55),
.B1(n_257),
.B2(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_29),
.B(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_29),
.A2(n_443),
.B(n_444),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_39),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.Y(n_39)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_37),
.Y(n_422)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_42),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_42),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_42),
.Y(n_156)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_45),
.Y(n_180)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_49),
.B(n_56),
.Y(n_212)
);

INVx8_ASAP7_75t_L g427 ( 
.A(n_51),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_55),
.B(n_274),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_55),
.A2(n_213),
.B(n_474),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_56),
.B(n_214),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g443 ( 
.A1(n_58),
.A2(n_274),
.B(n_425),
.Y(n_443)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_62),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_62),
.B1(n_100),
.B2(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_89),
.B(n_91),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_63),
.A2(n_271),
.B(n_275),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_63),
.A2(n_89),
.B1(n_303),
.B2(n_348),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_63),
.A2(n_275),
.B(n_348),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_63),
.A2(n_89),
.B1(n_451),
.B2(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_64),
.A2(n_90),
.B1(n_169),
.B2(n_175),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_64),
.A2(n_90),
.B1(n_169),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_64),
.A2(n_90),
.B1(n_204),
.B2(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_64),
.B(n_276),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_78),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_68),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_69),
.Y(n_206)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_SL g249 ( 
.A(n_75),
.Y(n_249)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_76),
.Y(n_453)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_78),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_84),
.B2(n_87),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_81),
.Y(n_299)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_83),
.Y(n_236)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_85),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_86),
.Y(n_285)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_89),
.A2(n_306),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_90),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_94),
.B(n_112),
.Y(n_376)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_95),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_97),
.Y(n_372)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_98),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_98),
.Y(n_278)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_124),
.B1(n_132),
.B2(n_133),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_132),
.B1(n_133),
.B2(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_102),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_102),
.A2(n_132),
.B1(n_179),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_102),
.A2(n_132),
.B1(n_387),
.B2(n_447),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_116),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_111),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_116),
.A2(n_125),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22x1_ASAP7_75t_L g477 ( 
.A1(n_116),
.A2(n_177),
.B1(n_394),
.B2(n_478),
.Y(n_477)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g305 ( 
.A(n_118),
.Y(n_305)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_123),
.Y(n_375)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g389 ( 
.A(n_128),
.Y(n_389)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_132),
.B(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_132),
.A2(n_387),
.B(n_393),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_137),
.Y(n_392)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_157),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_156),
.Y(n_355)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_156),
.Y(n_414)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_156),
.Y(n_424)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_156),
.Y(n_449)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_183),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_164),
.B(n_167),
.CI(n_183),
.CON(n_222),
.SN(n_222)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_167),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g282 ( 
.A(n_174),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_177),
.A2(n_354),
.B(n_358),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_177),
.B(n_394),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_177),
.A2(n_358),
.B(n_494),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B(n_211),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_203),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_211),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_185),
.A2(n_203),
.B1(n_228),
.B2(n_463),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_194),
.B(n_197),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_186),
.A2(n_197),
.B1(n_235),
.B2(n_240),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_186),
.A2(n_288),
.B(n_293),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_186),
.A2(n_274),
.B(n_293),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_186),
.A2(n_430),
.B1(n_431),
.B2(n_434),
.Y(n_429)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_187),
.B(n_296),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_187),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_187),
.A2(n_363),
.B1(n_398),
.B2(n_401),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_187),
.A2(n_435),
.B1(n_469),
.B2(n_470),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_193),
.Y(n_292)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_198),
.Y(n_399)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_200),
.Y(n_436)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_201),
.Y(n_365)
);

BUFx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_202),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_203),
.Y(n_463)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_261),
.B(n_520),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_222),
.B(n_223),
.Y(n_520)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_222),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.C(n_232),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_229),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_232),
.B(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_250),
.C(n_256),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_233),
.B(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_234),
.B(n_244),
.Y(n_488)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_235),
.Y(n_469)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_243),
.Y(n_433)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_245),
.Y(n_467)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_249),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_250),
.B(n_256),
.Y(n_461)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_251),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_260),
.Y(n_444)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI311xp33_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_457),
.A3(n_496),
.B1(n_514),
.C1(n_519),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_405),
.B(n_456),
.Y(n_264)
);

AO21x1_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_378),
.B(n_404),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_342),
.B(n_377),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_309),
.B(n_341),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_286),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_269),
.B(n_286),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_280),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_270),
.A2(n_280),
.B1(n_281),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_270),
.Y(n_339)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_SL g354 ( 
.A1(n_274),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_274),
.B(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_279),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_284),
.Y(n_400)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_300),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_301),
.C(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_291),
.Y(n_366)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_307),
.B2(n_308),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_332),
.B(n_340),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_318),
.B(n_331),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_330),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_330),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_326),
.B(n_329),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_328),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_362),
.B(n_367),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_338),
.Y(n_340)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_344),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_360),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_352),
.B2(n_353),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_352),
.C(n_360),
.Y(n_379)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI32xp33_ASAP7_75t_L g368 ( 
.A1(n_357),
.A2(n_369),
.A3(n_370),
.B1(n_373),
.B2(n_376),
.Y(n_368)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_368),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_368),
.Y(n_384)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_380),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_385),
.B2(n_403),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_384),
.C(n_403),
.Y(n_406)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_395),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_396),
.C(n_397),
.Y(n_437)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_406),
.B(n_407),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_440),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.Y(n_408)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_428),
.B2(n_429),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_411),
.B(n_428),
.Y(n_492)
);

OAI32xp33_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_415),
.A3(n_418),
.B1(n_421),
.B2(n_425),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_437),
.B(n_438),
.C(n_440),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_442),
.B1(n_445),
.B2(n_455),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_441),
.B(n_446),
.C(n_450),
.Y(n_505)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_450),
.Y(n_445)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_447),
.Y(n_494)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_482),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_458),
.A2(n_482),
.B(n_515),
.C(n_518),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_479),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_459),
.B(n_479),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.C(n_464),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_460),
.B(n_462),
.CI(n_464),
.CON(n_495),
.SN(n_495)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_472),
.C(n_477),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_468),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_468),
.Y(n_504)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_472),
.A2(n_473),
.B1(n_477),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_477),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_495),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_495),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_488),
.C(n_489),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_484),
.A2(n_485),
.B1(n_488),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_488),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_507),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.C(n_493),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_490),
.A2(n_491),
.B1(n_493),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_495),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_509),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_498),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_506),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_506),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_503),
.C(n_505),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_512),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_505),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_511),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_511),
.Y(n_516)
);

INVx8_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx13_ASAP7_75t_L g525 ( 
.A(n_522),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);


endmodule