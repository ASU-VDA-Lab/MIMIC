module fake_jpeg_31949_n_205 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_51),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_44),
.Y(n_72)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_56),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_48),
.B1(n_52),
.B2(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_32),
.B1(n_23),
.B2(n_29),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_23),
.B(n_22),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_32),
.B(n_26),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_33),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_42),
.B1(n_50),
.B2(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_32),
.B1(n_23),
.B2(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_84),
.B1(n_90),
.B2(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_43),
.C(n_46),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_62),
.C(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_31),
.Y(n_115)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_43),
.B(n_26),
.C(n_28),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_95),
.B1(n_99),
.B2(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_45),
.B1(n_29),
.B2(n_22),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_101),
.B1(n_70),
.B2(n_61),
.Y(n_116)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_21),
.B1(n_35),
.B2(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_95),
.B(n_103),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_49),
.B1(n_35),
.B2(n_31),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_56),
.A2(n_62),
.A3(n_69),
.B1(n_66),
.B2(n_72),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_72),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_73),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_105),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_103),
.B(n_88),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_129),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_121),
.B1(n_127),
.B2(n_131),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_61),
.B1(n_80),
.B2(n_67),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_82),
.B(n_106),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_2),
.B(n_3),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_73),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_102),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_79),
.B1(n_60),
.B2(n_67),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_73),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_104),
.C(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_136),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_85),
.B(n_91),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_128),
.B(n_125),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_128),
.B1(n_119),
.B2(n_110),
.C(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_98),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_3),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_92),
.C(n_82),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_94),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_97),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_126),
.B1(n_125),
.B2(n_5),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_87),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_49),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_129),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_60),
.B1(n_49),
.B2(n_89),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_117),
.B1(n_126),
.B2(n_114),
.Y(n_161)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

NOR2x1_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_16),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_R g166 ( 
.A(n_150),
.B(n_12),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_121),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_156),
.C(n_167),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_129),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_159),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_163),
.B(n_166),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_149),
.B1(n_148),
.B2(n_133),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_145),
.B1(n_141),
.B2(n_163),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_137),
.C(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_147),
.C(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_132),
.C(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_165),
.B1(n_162),
.B2(n_7),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_145),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_177),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_167),
.C(n_154),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_4),
.C(n_6),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_176),
.A2(n_158),
.B1(n_164),
.B2(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_6),
.C(n_7),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_186),
.B(n_8),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_173),
.B1(n_168),
.B2(n_10),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_173),
.B1(n_9),
.B2(n_10),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_189),
.B1(n_179),
.B2(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_8),
.B1(n_11),
.B2(n_183),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_11),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_194),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_180),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_191),
.A2(n_184),
.B(n_185),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_198),
.B(n_199),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_198),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_203),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);


endmodule