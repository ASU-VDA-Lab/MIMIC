module fake_jpeg_29735_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_26),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_25),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_52),
.B1(n_56),
.B2(n_53),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_84),
.C(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_85),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_56),
.B1(n_64),
.B2(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_67),
.B1(n_60),
.B2(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_54),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_64),
.B1(n_70),
.B2(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_58),
.B1(n_74),
.B2(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_5),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_58),
.B1(n_72),
.B2(n_71),
.Y(n_113)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_57),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_119),
.C(n_11),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_69),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_118),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_62),
.B1(n_28),
.B2(n_30),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_119),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_23),
.C(n_49),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_33),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_132),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_101),
.B1(n_100),
.B2(n_8),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_130),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_101),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_34),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_139),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_6),
.B(n_9),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_47),
.B(n_51),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_10),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_11),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_42),
.C(n_46),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_12),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_125),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_104),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_38),
.C(n_48),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_134),
.C(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_31),
.C(n_35),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_130),
.B1(n_146),
.B2(n_129),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_158),
.B(n_159),
.C(n_160),
.D(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_149),
.C(n_145),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.C(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_153),
.C(n_152),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_168),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_163),
.B(n_173),
.C(n_165),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_167),
.C(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_147),
.B1(n_138),
.B2(n_133),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_136),
.Y(n_179)
);


endmodule