module fake_jpeg_29854_n_144 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_15),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_31),
.B1(n_35),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_31),
.B1(n_33),
.B2(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_33),
.B1(n_30),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_48),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_35),
.B1(n_30),
.B2(n_34),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_24),
.B(n_14),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_18),
.B(n_21),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_44),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_19),
.C(n_6),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_41),
.B1(n_56),
.B2(n_60),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_75),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_41),
.B1(n_46),
.B2(n_44),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_60),
.B1(n_69),
.B2(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_65),
.B1(n_63),
.B2(n_25),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_58),
.C(n_56),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_94),
.C(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_95),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_93),
.B1(n_74),
.B2(n_76),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_14),
.C(n_19),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_19),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_76),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_84),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_97),
.B(n_111),
.C(n_107),
.D(n_89),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_83),
.B(n_72),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_81),
.B(n_2),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_94),
.C(n_86),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_101),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_92),
.B(n_93),
.C(n_73),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_118),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_100),
.C(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_1),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_19),
.C(n_6),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_110),
.C(n_105),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_5),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_3),
.C2(n_4),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_120),
.B(n_110),
.C(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_118),
.C(n_114),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_127),
.B1(n_113),
.B2(n_115),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_1),
.CI(n_4),
.CON(n_126),
.SN(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_131),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_123),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_135),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_137),
.B(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_131),
.Y(n_139)
);

AOI31xp33_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_122),
.A3(n_121),
.B(n_134),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_141),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_114),
.Y(n_144)
);


endmodule