module fake_jpeg_12643_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_51),
.B(n_60),
.Y(n_117)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_53),
.B(n_80),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_64),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_78),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_31),
.B(n_4),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g145 ( 
.A(n_81),
.Y(n_145)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_92),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_7),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_85),
.B(n_88),
.Y(n_139)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_89),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_43),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_91),
.B(n_94),
.Y(n_144)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_48),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_98),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_103),
.Y(n_126)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_102),
.Y(n_150)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_19),
.B1(n_32),
.B2(n_35),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_105),
.A2(n_115),
.B1(n_124),
.B2(n_128),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_19),
.B1(n_32),
.B2(n_35),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_116),
.B(n_143),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_34),
.B1(n_50),
.B2(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_50),
.B1(n_99),
.B2(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_53),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_80),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_148),
.B(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_63),
.B(n_66),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_71),
.A2(n_80),
.B(n_53),
.C(n_85),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_118),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_69),
.A2(n_81),
.B1(n_39),
.B2(n_52),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_153),
.B1(n_142),
.B2(n_130),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_72),
.A2(n_58),
.B1(n_57),
.B2(n_69),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_144),
.B(n_126),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_159),
.B(n_161),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_163),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_129),
.A2(n_137),
.B1(n_153),
.B2(n_119),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_173),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_155),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_117),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_172),
.Y(n_197)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_104),
.B(n_113),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_168),
.B(n_174),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_125),
.C(n_155),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_134),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_108),
.B(n_138),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_176),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_108),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_185),
.Y(n_199)
);

AO22x1_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_152),
.B1(n_118),
.B2(n_133),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_174),
.B(n_179),
.C(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_154),
.B(n_122),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_188),
.Y(n_202)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_165),
.B1(n_174),
.B2(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_122),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_193),
.Y(n_205)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_127),
.B(n_154),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_127),
.CI(n_160),
.CON(n_204),
.SN(n_204)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_210),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_158),
.B(n_164),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_221),
.B(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_213),
.B1(n_182),
.B2(n_178),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_219),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_163),
.B1(n_195),
.B2(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_157),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_209),
.B(n_170),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_229),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_178),
.C(n_163),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_210),
.C(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_238),
.B1(n_218),
.B2(n_220),
.Y(n_252)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_235),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_199),
.A2(n_182),
.B1(n_167),
.B2(n_188),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_233),
.B(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_193),
.B1(n_211),
.B2(n_200),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_242),
.B1(n_219),
.B2(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_216),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_198),
.B1(n_205),
.B2(n_206),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_250),
.Y(n_266)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_233),
.B(n_236),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_258),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_200),
.B1(n_199),
.B2(n_208),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_220),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_226),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_218),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_254),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_267),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_248),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_268),
.C(n_257),
.Y(n_275)
);

OA21x2_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_204),
.B(n_229),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_227),
.B1(n_246),
.B2(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_266),
.C(n_264),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_263),
.B(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_247),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_265),
.B1(n_251),
.B2(n_196),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_204),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_268),
.C(n_255),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_279),
.B(n_270),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_285),
.C(n_205),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_280),
.B1(n_276),
.B2(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_271),
.B1(n_237),
.B2(n_220),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_273),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_295),
.B1(n_293),
.B2(n_273),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_266),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_260),
.Y(n_298)
);


endmodule