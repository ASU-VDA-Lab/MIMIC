module real_jpeg_6148_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_105;
wire n_40;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_1),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_173),
.B1(n_177),
.B2(n_181),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_3),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_95),
.B1(n_122),
.B2(n_131),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_194),
.C(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_4),
.B(n_119),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_4),
.B(n_29),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_4),
.B(n_99),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_81),
.B1(n_101),
.B2(n_104),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_5),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_5),
.A2(n_104),
.B1(n_173),
.B2(n_199),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_6),
.A2(n_38),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_38),
.B1(n_82),
.B2(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_8),
.Y(n_228)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_11),
.A2(n_94),
.B1(n_152),
.B2(n_157),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_11),
.A2(n_94),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_185),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_183),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_141),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_16),
.B(n_141),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_70),
.C(n_105),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_17),
.B(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_18),
.B(n_41),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_28),
.B(n_30),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_20),
.A2(n_31),
.B1(n_33),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_21),
.Y(n_221)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_24),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_28),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_30),
.A2(n_220),
.B(n_226),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_31),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_31),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_37),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_39),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_84)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.A3(n_54),
.B1(n_59),
.B2(n_64),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_48),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_48),
.Y(n_156)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_70),
.A2(n_105),
.B1(n_106),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_91),
.B1(n_98),
.B2(n_100),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_71),
.A2(n_100),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_71),
.A2(n_145),
.B(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_72),
.B(n_146),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_84),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_75),
.B(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_84),
.A2(n_91),
.B(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_127),
.B(n_133),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_117),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_119),
.Y(n_140)
);

AO22x2_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_131),
.B(n_132),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_131),
.A2(n_200),
.B(n_201),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_151),
.B(n_158),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_149),
.B2(n_182),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_160),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_171),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_243),
.B(n_248),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_209),
.B(n_242),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_196),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_204),
.C(n_208),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_231),
.B(n_241),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_218),
.B(n_230),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_229),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_229),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_239),
.Y(n_241)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);


endmodule