module fake_netlist_6_1965_n_1710 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1710);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1710;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_56),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_42),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx11_ASAP7_75t_R g160 ( 
.A(n_67),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_52),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_28),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_21),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_88),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_13),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_30),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_42),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_34),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_31),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_15),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_21),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_58),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_22),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_76),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_72),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_66),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_53),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_51),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_107),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_39),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_65),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_79),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_4),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_0),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_69),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_98),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_70),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_29),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_150),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_83),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_51),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_12),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_115),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_71),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_103),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_81),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_94),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_96),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_110),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_19),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_55),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_92),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_140),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_19),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_9),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_50),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_61),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_108),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_44),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_24),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_113),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_11),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_129),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_25),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_26),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_85),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_30),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_130),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_10),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_101),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_133),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_62),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_73),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_93),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_111),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_5),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_28),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_105),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_32),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_32),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_16),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_80),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_29),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_152),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_77),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_114),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_91),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_23),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_127),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_40),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_13),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_134),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_119),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_104),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_89),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_59),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_17),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_131),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_78),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_23),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_102),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_84),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_68),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_20),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_100),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_9),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_2),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_18),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_138),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_40),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_53),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_149),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_3),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_251),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_160),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_191),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_200),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_180),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_241),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_241),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_231),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_284),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_166),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_215),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_195),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_156),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_178),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_166),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_170),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_162),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_226),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_174),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_265),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_181),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_199),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_192),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_212),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_166),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_182),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_201),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_226),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_228),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_226),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_243),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_252),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_244),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_203),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_245),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_255),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_207),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_230),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_267),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_182),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_210),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_276),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_277),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_182),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_159),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_172),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_240),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_226),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_213),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_294),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_295),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_240),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_214),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_307),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_221),
.Y(n_391)
);

NOR2x1_ASAP7_75t_L g392 ( 
.A(n_314),
.B(n_172),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_316),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_318),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_335),
.A2(n_184),
.B1(n_232),
.B2(n_308),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_221),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g409 ( 
.A(n_332),
.B(n_161),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_370),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_339),
.B(n_155),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_380),
.B(n_240),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_380),
.B(n_155),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_339),
.B(n_254),
.Y(n_416)
);

OAI21x1_ASAP7_75t_L g417 ( 
.A1(n_349),
.A2(n_176),
.B(n_161),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_330),
.B(n_254),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_324),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_340),
.Y(n_423)
);

AND2x2_ASAP7_75t_SL g424 ( 
.A(n_333),
.B(n_176),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_179),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_330),
.B(n_208),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_334),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

INVx6_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_331),
.B(n_179),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_329),
.A2(n_281),
.B1(n_308),
.B2(n_177),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_354),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_311),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_336),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_353),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_343),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_359),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_353),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_355),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_320),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_331),
.B(n_157),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_320),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_321),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_321),
.A2(n_220),
.B(n_185),
.Y(n_456)
);

XNOR2x2_ASAP7_75t_L g457 ( 
.A(n_356),
.B(n_185),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_325),
.A2(n_177),
.B1(n_173),
.B2(n_304),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_361),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_337),
.B(n_157),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_447),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_438),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_444),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_369),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_373),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_437),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_409),
.B(n_385),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_438),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_409),
.B(n_385),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_437),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_426),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_426),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_457),
.A2(n_364),
.B1(n_326),
.B2(n_348),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_423),
.Y(n_491)
);

INVx8_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_424),
.B(n_357),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_412),
.B(n_358),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_412),
.B(n_391),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_395),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_416),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_L g500 ( 
.A1(n_458),
.A2(n_227),
.B1(n_198),
.B2(n_234),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_424),
.B(n_366),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_419),
.B(n_391),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_406),
.B(n_343),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_389),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_424),
.B(n_372),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_406),
.B(n_230),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_442),
.B(n_429),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_416),
.B(n_343),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_457),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_420),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_457),
.A2(n_220),
.B1(n_343),
.B2(n_383),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_416),
.B(n_343),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_390),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_429),
.B(n_407),
.Y(n_520)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_456),
.A2(n_194),
.B(n_188),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_407),
.B(n_382),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_206),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_393),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_416),
.B(n_343),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_399),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

NOR2x1p5_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_312),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_437),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_400),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_450),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_394),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_400),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_394),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_451),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_456),
.A2(n_235),
.B(n_197),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_451),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_451),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_437),
.B(n_343),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_418),
.B(n_337),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_392),
.B(n_343),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_418),
.B(n_338),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_417),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_417),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_415),
.B(n_386),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_414),
.B(n_345),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_392),
.B(n_218),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_461),
.B(n_363),
.C(n_361),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_458),
.B(n_158),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_402),
.B(n_219),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_402),
.B(n_222),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_440),
.A2(n_257),
.B1(n_230),
.B2(n_378),
.Y(n_565)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_456),
.A2(n_249),
.B(n_236),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_433),
.B(n_158),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_440),
.B(n_322),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_420),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_401),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_440),
.B(n_322),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_401),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_441),
.A2(n_173),
.B1(n_171),
.B2(n_164),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_402),
.B(n_223),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_451),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_408),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_436),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_404),
.B(n_224),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_408),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_440),
.B(n_261),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_411),
.Y(n_582)
);

AND3x2_ASAP7_75t_L g583 ( 
.A(n_433),
.B(n_271),
.C(n_266),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_436),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_404),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_455),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_439),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_403),
.B(n_164),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_455),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_404),
.Y(n_593)
);

AND2x2_ASAP7_75t_SL g594 ( 
.A(n_446),
.B(n_230),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_455),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_411),
.B(n_323),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_427),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_427),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_413),
.B(n_323),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_441),
.B(n_163),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_460),
.B(n_272),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_413),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_428),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_428),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_446),
.B(n_230),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_403),
.B(n_171),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_455),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_432),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_405),
.B(n_225),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_484),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_478),
.B(n_396),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_495),
.B(n_446),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_512),
.A2(n_279),
.B1(n_290),
.B2(n_285),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_489),
.B(n_163),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_460),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_594),
.B(n_454),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_476),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_594),
.B(n_503),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_594),
.B(n_454),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_485),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_511),
.B(n_257),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_485),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_552),
.Y(n_624)
);

NOR2x1p5_ASAP7_75t_L g625 ( 
.A(n_494),
.B(n_281),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_552),
.B(n_226),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_552),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_570),
.B(n_454),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_533),
.B(n_459),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_502),
.B(n_459),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_556),
.B(n_165),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_570),
.B(n_405),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_487),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_548),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_572),
.B(n_410),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_576),
.B(n_410),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_515),
.B(n_257),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_527),
.B(n_257),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_410),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_518),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_604),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_536),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_548),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_518),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_580),
.B(n_582),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_555),
.B(n_434),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_580),
.B(n_421),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_L g650 ( 
.A(n_501),
.B(n_434),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_475),
.B(n_257),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_496),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_582),
.B(n_421),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_475),
.B(n_226),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_603),
.B(n_421),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_299),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_604),
.B(n_435),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_499),
.B(n_435),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_552),
.B(n_557),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_496),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_504),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_608),
.B(n_445),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_608),
.Y(n_663)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_557),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_504),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_558),
.B(n_445),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_512),
.A2(n_452),
.B(n_449),
.C(n_448),
.Y(n_667)
);

AND2x2_ASAP7_75t_SL g668 ( 
.A(n_514),
.B(n_448),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_499),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_558),
.B(n_449),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_474),
.B(n_165),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_568),
.B(n_571),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_552),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_510),
.B(n_167),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_475),
.B(n_226),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_497),
.B(n_452),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_R g678 ( 
.A(n_473),
.B(n_167),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_475),
.B(n_226),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_492),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_497),
.B(n_246),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_505),
.B(n_248),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_505),
.B(n_506),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_476),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_516),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_571),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_577),
.B(n_242),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_517),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_602),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_488),
.B(n_196),
.C(n_193),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_506),
.B(n_253),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_588),
.B(n_363),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_577),
.B(n_486),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_588),
.B(n_365),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_551),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_528),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_596),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_480),
.B(n_168),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_502),
.B(n_365),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_520),
.A2(n_387),
.B(n_384),
.C(n_378),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_596),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_560),
.A2(n_387),
.B(n_384),
.C(n_375),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_507),
.B(n_256),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_507),
.B(n_519),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_524),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_523),
.A2(n_282),
.B1(n_296),
.B2(n_297),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_577),
.B(n_242),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_525),
.B(n_258),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_599),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_525),
.B(n_270),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_560),
.A2(n_375),
.B(n_374),
.C(n_371),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_494),
.B(n_367),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_528),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_577),
.B(n_242),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_486),
.B(n_242),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_581),
.B(n_601),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_482),
.B(n_374),
.C(n_371),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_523),
.A2(n_282),
.B1(n_296),
.B2(n_297),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_489),
.B(n_367),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_601),
.A2(n_242),
.B1(n_301),
.B2(n_303),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_583),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_493),
.B(n_168),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_523),
.A2(n_169),
.B1(n_183),
.B2(n_186),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_523),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_529),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_526),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_526),
.B(n_274),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_486),
.B(n_242),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_534),
.B(n_169),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_534),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_523),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_532),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_554),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_598),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_492),
.B(n_187),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_492),
.B(n_189),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_567),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_492),
.B(n_483),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_544),
.B(n_242),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_559),
.B(n_189),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_544),
.B(n_242),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_522),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_492),
.B(n_584),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_584),
.B(n_190),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_601),
.B(n_190),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_489),
.B(n_368),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_535),
.Y(n_751)
);

INVx8_ASAP7_75t_L g752 ( 
.A(n_581),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_535),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_508),
.B(n_280),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_R g755 ( 
.A(n_473),
.B(n_280),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_601),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_553),
.B(n_368),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_489),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_549),
.B(n_287),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_549),
.B(n_287),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_553),
.B(n_288),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_537),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_581),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_465),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_465),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_565),
.A2(n_288),
.B1(n_289),
.B2(n_309),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_467),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_544),
.B(n_550),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_549),
.B(n_289),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_467),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_561),
.A2(n_292),
.B1(n_293),
.B2(n_309),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_581),
.B(n_327),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_581),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_L g774 ( 
.A(n_544),
.B(n_292),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_664),
.B(n_544),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_631),
.B(n_537),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_610),
.Y(n_777)
);

AND2x6_ASAP7_75t_SL g778 ( 
.A(n_611),
.B(n_589),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_746),
.B(n_600),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_610),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_671),
.B(n_668),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_650),
.B(n_569),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_612),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_737),
.B(n_569),
.C(n_573),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_669),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_672),
.B(n_530),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_678),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_680),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_629),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_741),
.B(n_500),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_684),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_692),
.B(n_530),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_694),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_668),
.B(n_538),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_721),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_729),
.B(n_538),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_750),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_621),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_SL g801 ( 
.A1(n_642),
.A2(n_589),
.B1(n_597),
.B2(n_513),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_623),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_619),
.A2(n_566),
.B(n_541),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_701),
.B(n_462),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_680),
.Y(n_805)
);

INVx5_ASAP7_75t_L g806 ( 
.A(n_680),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_757),
.A2(n_606),
.B1(n_509),
.B2(n_573),
.Y(n_807)
);

OAI21xp33_ASAP7_75t_SL g808 ( 
.A1(n_733),
.A2(n_609),
.B(n_562),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_757),
.A2(n_605),
.B1(n_463),
.B2(n_466),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_623),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_678),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_646),
.B(n_491),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_633),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_664),
.B(n_540),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_633),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_755),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_756),
.A2(n_574),
.B1(n_563),
.B2(n_579),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_674),
.B(n_540),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_616),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_664),
.B(n_542),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_635),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_664),
.B(n_542),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_664),
.B(n_463),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_664),
.B(n_544),
.Y(n_824)
);

NOR2x1_ASAP7_75t_R g825 ( 
.A(n_758),
.B(n_293),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_680),
.B(n_479),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_669),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_635),
.B(n_464),
.Y(n_828)
);

AND3x1_ASAP7_75t_L g829 ( 
.A(n_734),
.B(n_327),
.C(n_328),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_634),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_641),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_669),
.B(n_479),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_736),
.B(n_740),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_736),
.B(n_479),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_714),
.B(n_328),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_718),
.B(n_585),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_648),
.B(n_466),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_761),
.A2(n_468),
.B(n_469),
.C(n_477),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_736),
.A2(n_521),
.B1(n_490),
.B2(n_498),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_672),
.B(n_468),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_672),
.B(n_469),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_740),
.B(n_479),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_755),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_695),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_SL g845 ( 
.A(n_625),
.B(n_298),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_695),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_693),
.A2(n_547),
.B(n_490),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_758),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_644),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_689),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_647),
.B(n_477),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_630),
.Y(n_852)
);

OR2x2_ASAP7_75t_SL g853 ( 
.A(n_690),
.B(n_204),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_676),
.A2(n_545),
.B1(n_539),
.B2(n_595),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_683),
.B(n_470),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_645),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_706),
.B(n_470),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_725),
.A2(n_205),
.B1(n_209),
.B2(n_211),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_757),
.A2(n_605),
.B1(n_481),
.B2(n_471),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_724),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_707),
.B(n_471),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_658),
.B(n_657),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_762),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_624),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_752),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_740),
.A2(n_521),
.B1(n_479),
.B2(n_498),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_757),
.A2(n_605),
.B1(n_481),
.B2(n_472),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_752),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_686),
.A2(n_586),
.B1(n_539),
.B2(n_595),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_696),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_708),
.B(n_490),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_658),
.B(n_472),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_490),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_658),
.B(n_490),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_R g875 ( 
.A(n_615),
.B(n_298),
.Y(n_875)
);

OR2x2_ASAP7_75t_SL g876 ( 
.A(n_699),
.B(n_216),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_662),
.B(n_498),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_754),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_752),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_703),
.B(n_498),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_652),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_693),
.A2(n_498),
.B(n_531),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_752),
.B(n_543),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_711),
.B(n_723),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_718),
.B(n_531),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_SL g886 ( 
.A(n_771),
.B(n_614),
.C(n_700),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_677),
.B(n_531),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_726),
.B(n_217),
.C(n_229),
.Y(n_888)
);

AO22x1_ASAP7_75t_L g889 ( 
.A1(n_718),
.A2(n_233),
.B1(n_278),
.B2(n_237),
.Y(n_889)
);

AO22x1_ASAP7_75t_L g890 ( 
.A1(n_719),
.A2(n_238),
.B1(n_275),
.B2(n_239),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_660),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_661),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_757),
.A2(n_605),
.B1(n_247),
.B2(n_259),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_661),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_643),
.B(n_663),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_772),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_772),
.B(n_543),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_667),
.B(n_531),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_624),
.B(n_531),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_624),
.B(n_593),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_SL g901 ( 
.A1(n_766),
.A2(n_260),
.B1(n_262),
.B2(n_269),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_727),
.B(n_300),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_665),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_666),
.B(n_585),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_763),
.B(n_607),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_732),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_757),
.A2(n_605),
.B1(n_607),
.B2(n_575),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_685),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_670),
.B(n_585),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_685),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_749),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_627),
.B(n_593),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_722),
.B(n_300),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_627),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_627),
.B(n_593),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_763),
.B(n_306),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_773),
.A2(n_578),
.B1(n_545),
.B2(n_592),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_673),
.B(n_688),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_681),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_688),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_773),
.B(n_586),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_673),
.B(n_593),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_697),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_659),
.A2(n_578),
.B1(n_546),
.B2(n_592),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_697),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_SL g926 ( 
.A(n_702),
.B(n_306),
.C(n_546),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_673),
.B(n_593),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_698),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_613),
.B(n_591),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_682),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_698),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_715),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_617),
.B(n_591),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_748),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_656),
.B(n_590),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_728),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_620),
.B(n_575),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_747),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_691),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_728),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_735),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_735),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_751),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_705),
.B(n_564),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_753),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_764),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_742),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_632),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_775),
.A2(n_659),
.B(n_768),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_919),
.B(n_781),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_871),
.A2(n_761),
.B(n_626),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_786),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_868),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_798),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_775),
.A2(n_824),
.B(n_823),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_786),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_SL g957 ( 
.A1(n_878),
.A2(n_738),
.B1(n_739),
.B2(n_712),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_868),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_807),
.A2(n_704),
.B1(n_713),
.B2(n_628),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_804),
.B(n_704),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_824),
.A2(n_768),
.B(n_774),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_896),
.B(n_865),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_800),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_777),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_906),
.B(n_744),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_862),
.A2(n_774),
.B(n_626),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_814),
.A2(n_651),
.B(n_717),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_792),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_802),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_792),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_819),
.B(n_710),
.Y(n_971)
);

AO31x2_ASAP7_75t_L g972 ( 
.A1(n_839),
.A2(n_713),
.A3(n_655),
.B(n_637),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_886),
.A2(n_730),
.B1(n_769),
.B2(n_759),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_791),
.A2(n_760),
.B(n_622),
.C(n_639),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_820),
.A2(n_651),
.B(n_717),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_788),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_794),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_780),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_779),
.A2(n_902),
.B(n_791),
.C(n_888),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_799),
.B(n_636),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_850),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_939),
.B(n_765),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_783),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_789),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_930),
.B(n_796),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_SL g986 ( 
.A(n_789),
.B(n_654),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_822),
.A2(n_731),
.B(n_709),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_790),
.B(n_640),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_779),
.A2(n_653),
.B(n_649),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_794),
.B(n_622),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_810),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_L g992 ( 
.A(n_801),
.B(n_731),
.C(n_687),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_844),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_807),
.A2(n_770),
.B1(n_767),
.B2(n_765),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_795),
.A2(n_767),
.B1(n_638),
.B2(n_639),
.Y(n_995)
);

OAI21xp33_ASAP7_75t_L g996 ( 
.A1(n_902),
.A2(n_638),
.B(n_679),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_911),
.A2(n_873),
.B(n_871),
.C(n_913),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_852),
.B(n_679),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_782),
.A2(n_687),
.B(n_654),
.C(n_716),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_815),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_835),
.B(n_675),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_948),
.B(n_675),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_852),
.B(n_793),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_789),
.A2(n_716),
.B(n_709),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_844),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_873),
.A2(n_745),
.B(n_743),
.C(n_564),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_846),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_813),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_808),
.A2(n_605),
.B(n_3),
.C(n_5),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_856),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_884),
.B(n_811),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_816),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_784),
.B(n_1),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_897),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_R g1015 ( 
.A(n_843),
.B(n_848),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_934),
.A2(n_605),
.B1(n_153),
.B2(n_151),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_856),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_805),
.A2(n_147),
.B(n_146),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_805),
.A2(n_142),
.B(n_135),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_907),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_868),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_805),
.A2(n_806),
.B(n_887),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_870),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_858),
.A2(n_11),
.B(n_14),
.C(n_17),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_805),
.B(n_124),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_875),
.A2(n_812),
.B(n_895),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_806),
.A2(n_915),
.B(n_912),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_946),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_830),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_778),
.B(n_121),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_907),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_1031)
);

INVx8_ASAP7_75t_L g1032 ( 
.A(n_883),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_806),
.A2(n_922),
.B(n_833),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_812),
.B(n_24),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_870),
.A2(n_25),
.B(n_27),
.C(n_33),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_809),
.A2(n_864),
.B1(n_867),
.B2(n_859),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_833),
.A2(n_99),
.B(n_97),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_851),
.B(n_90),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_891),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_SL g1040 ( 
.A(n_875),
.B(n_27),
.C(n_33),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_853),
.B(n_34),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_845),
.B(n_82),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_947),
.B(n_75),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_787),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_947),
.B(n_74),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_831),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_818),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_868),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_787),
.A2(n_57),
.B1(n_36),
.B2(n_37),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_947),
.B(n_35),
.Y(n_1050)
);

NAND2x1_ASAP7_75t_SL g1051 ( 
.A(n_865),
.B(n_38),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_879),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_776),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_879),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_860),
.B(n_46),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_923),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_821),
.A2(n_48),
.B(n_49),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_866),
.A2(n_48),
.B(n_49),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_916),
.B(n_54),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_855),
.B(n_54),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_944),
.A2(n_55),
.B(n_877),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_828),
.A2(n_863),
.B(n_945),
.C(n_943),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_901),
.A2(n_840),
.B(n_841),
.C(n_872),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_829),
.A2(n_947),
.B1(n_885),
.B2(n_921),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_889),
.B(n_890),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_847),
.A2(n_882),
.B(n_904),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_876),
.B(n_825),
.Y(n_1068)
);

XNOR2xp5_ASAP7_75t_L g1069 ( 
.A(n_836),
.B(n_883),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_837),
.B(n_880),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_879),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_857),
.B(n_861),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_785),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_883),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_909),
.A2(n_874),
.B(n_842),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_785),
.B(n_827),
.Y(n_1076)
);

NOR2xp67_ASAP7_75t_L g1077 ( 
.A(n_925),
.B(n_942),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_931),
.B(n_885),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_914),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_898),
.A2(n_797),
.B(n_926),
.C(n_933),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_914),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_933),
.A2(n_937),
.B(n_929),
.C(n_838),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_914),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_928),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_918),
.A2(n_929),
.B(n_900),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_893),
.A2(n_941),
.B(n_940),
.C(n_936),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_SL g1087 ( 
.A1(n_817),
.A2(n_937),
.B(n_832),
.C(n_803),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_979),
.A2(n_893),
.B(n_917),
.C(n_869),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1029),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_951),
.A2(n_903),
.A3(n_920),
.B(n_910),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_1062),
.A2(n_826),
.B(n_832),
.C(n_834),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1046),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_957),
.A2(n_938),
.B1(n_921),
.B2(n_905),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_993),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1013),
.A2(n_826),
.B1(n_854),
.B2(n_834),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1087),
.A2(n_924),
.B(n_842),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_997),
.A2(n_1080),
.B(n_959),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1067),
.A2(n_927),
.B(n_900),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_952),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_1009),
.A2(n_899),
.B(n_849),
.C(n_881),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_966),
.A2(n_1072),
.B(n_987),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_967),
.A2(n_931),
.B(n_938),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_996),
.A2(n_932),
.B(n_892),
.C(n_894),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_974),
.A2(n_908),
.B(n_899),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1036),
.A2(n_931),
.B1(n_836),
.B2(n_905),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_975),
.A2(n_935),
.B(n_914),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_980),
.B(n_935),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_968),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_1007),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1003),
.B(n_935),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1011),
.B(n_905),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1070),
.B(n_1026),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_956),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_998),
.B(n_971),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_970),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_954),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1041),
.A2(n_1064),
.B(n_992),
.C(n_1063),
.Y(n_1117)
);

AOI21x1_ASAP7_75t_L g1118 ( 
.A1(n_995),
.A2(n_961),
.B(n_1075),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_SL g1119 ( 
.A(n_1071),
.B(n_984),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_959),
.A2(n_995),
.A3(n_1086),
.B(n_994),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1017),
.B(n_981),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1038),
.A2(n_1002),
.B(n_949),
.Y(n_1122)
);

AOI22x1_ASAP7_75t_L g1123 ( 
.A1(n_1059),
.A2(n_1078),
.B1(n_1033),
.B2(n_955),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_SL g1124 ( 
.A1(n_1024),
.A2(n_1035),
.B1(n_1031),
.B2(n_1020),
.C(n_1054),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_962),
.B(n_1074),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_994),
.A2(n_1006),
.A3(n_1038),
.B(n_1036),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1023),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1017),
.B(n_1005),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1005),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_963),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_1081),
.B(n_953),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_969),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_991),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1027),
.A2(n_1082),
.B(n_1022),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_SL g1135 ( 
.A1(n_1066),
.A2(n_1061),
.B(n_1060),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_999),
.A2(n_1061),
.B(n_973),
.C(n_1001),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_977),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_1002),
.B(n_1004),
.Y(n_1138)
);

AO21x1_ASAP7_75t_L g1139 ( 
.A1(n_1020),
.A2(n_1031),
.B(n_989),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1028),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1000),
.Y(n_1141)
);

BUFx2_ASAP7_75t_R g1142 ( 
.A(n_976),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_962),
.B(n_1074),
.Y(n_1143)
);

NAND3x1_ASAP7_75t_L g1144 ( 
.A(n_1068),
.B(n_1049),
.C(n_1065),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1014),
.B(n_985),
.Y(n_1145)
);

O2A1O1Ixp5_ASAP7_75t_L g1146 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_1050),
.C(n_986),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1083),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1039),
.Y(n_1148)
);

AOI221x1_ASAP7_75t_L g1149 ( 
.A1(n_1047),
.A2(n_1040),
.B1(n_1037),
.B2(n_1018),
.C(n_1019),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_1077),
.A2(n_988),
.B(n_990),
.Y(n_1150)
);

OAI22x1_ASAP7_75t_L g1151 ( 
.A1(n_1034),
.A2(n_1069),
.B1(n_965),
.B2(n_1010),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1015),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1057),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_982),
.B(n_983),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1014),
.B(n_1008),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1053),
.A2(n_1056),
.B(n_1042),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1084),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1074),
.A2(n_1081),
.B1(n_1032),
.B2(n_964),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_978),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1016),
.A2(n_1025),
.B(n_1073),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1079),
.B(n_972),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1076),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1051),
.A2(n_972),
.B(n_1081),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1030),
.A2(n_953),
.B(n_958),
.Y(n_1164)
);

OAI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_958),
.A2(n_1055),
.B(n_1021),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1032),
.A2(n_958),
.B(n_1021),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1021),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1044),
.A2(n_1048),
.B1(n_1052),
.B2(n_1055),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1044),
.A2(n_1048),
.B(n_1052),
.C(n_1055),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1029),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1029),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_979),
.B(n_631),
.C(n_878),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_SL g1173 ( 
.A(n_1071),
.B(n_758),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_950),
.B(n_960),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_L g1175 ( 
.A(n_992),
.B(n_878),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_962),
.B(n_865),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_979),
.A2(n_631),
.B(n_1013),
.C(n_997),
.Y(n_1177)
);

INVxp67_ASAP7_75t_SL g1178 ( 
.A(n_993),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_966),
.A2(n_693),
.B(n_577),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1067),
.A2(n_1085),
.B(n_997),
.Y(n_1180)
);

AND2x2_ASAP7_75t_SL g1181 ( 
.A(n_1013),
.B(n_615),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_957),
.A2(n_878),
.B1(n_501),
.B2(n_335),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_984),
.Y(n_1183)
);

BUFx2_ASAP7_75t_SL g1184 ( 
.A(n_1012),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_979),
.B(n_631),
.C(n_878),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_968),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1085),
.A2(n_1067),
.B(n_949),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_979),
.A2(n_589),
.B(n_555),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_SL g1189 ( 
.A1(n_1058),
.A2(n_951),
.B(n_1059),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1087),
.A2(n_997),
.B(n_974),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_951),
.A2(n_959),
.A3(n_997),
.B(n_1067),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_950),
.B(n_960),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_950),
.B(n_960),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_997),
.A2(n_512),
.B1(n_878),
.B2(n_781),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_979),
.A2(n_997),
.B(n_779),
.C(n_781),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1066),
.A2(n_781),
.B(n_1061),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_997),
.A2(n_512),
.B1(n_878),
.B2(n_781),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1059),
.A2(n_997),
.B1(n_1009),
.B2(n_1062),
.C(n_1013),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1029),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_979),
.A2(n_1059),
.B(n_781),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_997),
.A2(n_512),
.B1(n_878),
.B2(n_781),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_950),
.B(n_878),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1029),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1085),
.A2(n_1067),
.B(n_949),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_968),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_950),
.B(n_781),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1085),
.A2(n_1067),
.B(n_949),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_950),
.B(n_781),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_979),
.B(n_631),
.C(n_878),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1085),
.A2(n_1067),
.B(n_949),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1029),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_968),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_950),
.B(n_781),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_997),
.A2(n_512),
.B1(n_878),
.B2(n_781),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_962),
.B(n_865),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1101),
.A2(n_1122),
.B(n_1179),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1199),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1203),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1167),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1190),
.A2(n_1097),
.B(n_1189),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1089),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1170),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1176),
.B(n_1215),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1181),
.A2(n_1139),
.B1(n_1185),
.B2(n_1209),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1210),
.A2(n_1098),
.B(n_1134),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1190),
.A2(n_1097),
.B(n_1198),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_1188),
.B(n_1172),
.C(n_1177),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1171),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1175),
.A2(n_1202),
.B1(n_1182),
.B2(n_1144),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1174),
.B(n_1192),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_1112),
.A2(n_1194),
.B(n_1201),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1106),
.A2(n_1118),
.B(n_1123),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_1119),
.B(n_1173),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1176),
.Y(n_1234)
);

AO21x2_ASAP7_75t_L g1235 ( 
.A1(n_1096),
.A2(n_1138),
.B(n_1163),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1117),
.A2(n_1195),
.B(n_1136),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1215),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1096),
.A2(n_1138),
.B(n_1200),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1111),
.B(n_1193),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1162),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1099),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1095),
.A2(n_1105),
.B(n_1161),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1108),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1146),
.A2(n_1114),
.B(n_1088),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1194),
.A2(n_1214),
.B1(n_1201),
.B2(n_1197),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1196),
.A2(n_1135),
.B(n_1104),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1104),
.A2(n_1091),
.B(n_1163),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1180),
.A2(n_1161),
.B(n_1105),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1186),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1151),
.A2(n_1214),
.B1(n_1197),
.B2(n_1152),
.Y(n_1250)
);

INVx3_ASAP7_75t_SL g1251 ( 
.A(n_1128),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1211),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1107),
.A2(n_1158),
.B(n_1160),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1092),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1142),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1180),
.A2(n_1149),
.B(n_1158),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1206),
.B(n_1208),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1116),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1130),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1131),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1213),
.B(n_1156),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1184),
.A2(n_1129),
.B1(n_1178),
.B2(n_1109),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1132),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1110),
.A2(n_1093),
.B(n_1166),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1131),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1169),
.B(n_1164),
.Y(n_1266)
);

BUFx2_ASAP7_75t_R g1267 ( 
.A(n_1205),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1125),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1168),
.A2(n_1133),
.B(n_1141),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1090),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1113),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1124),
.A2(n_1103),
.B(n_1155),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_L g1273 ( 
.A(n_1212),
.B(n_1115),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1148),
.A2(n_1159),
.B(n_1157),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1090),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1127),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1153),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1090),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1140),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1137),
.B(n_1099),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1191),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1183),
.A2(n_1145),
.B(n_1147),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1147),
.A2(n_1154),
.B(n_1165),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1100),
.A2(n_1121),
.B(n_1094),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1125),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1150),
.A2(n_1191),
.B(n_1120),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1120),
.A2(n_1126),
.B(n_1150),
.Y(n_1287)
);

INVx2_ASAP7_75t_R g1288 ( 
.A(n_1120),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1126),
.A2(n_1167),
.B(n_1143),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1143),
.B(n_1126),
.Y(n_1290)
);

AOI222xp33_ASAP7_75t_L g1291 ( 
.A1(n_1188),
.A2(n_403),
.B1(n_589),
.B2(n_1181),
.C1(n_414),
.C2(n_784),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1172),
.A2(n_1209),
.B(n_1185),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1129),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1119),
.B(n_865),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1188),
.A2(n_878),
.B1(n_1181),
.B2(n_555),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1187),
.A2(n_1207),
.B(n_1204),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1101),
.A2(n_1122),
.B(n_1179),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1152),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1199),
.Y(n_1299)
);

INVxp33_ASAP7_75t_L g1300 ( 
.A(n_1202),
.Y(n_1300)
);

NOR2xp67_ASAP7_75t_L g1301 ( 
.A(n_1172),
.B(n_976),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1199),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1174),
.B(n_1192),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1152),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1162),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1187),
.A2(n_1207),
.B(n_1204),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1199),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1176),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1177),
.A2(n_979),
.B(n_1188),
.C(n_997),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1172),
.A2(n_1209),
.B(n_1185),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1125),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1188),
.A2(n_878),
.B1(n_1181),
.B2(n_555),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1199),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1176),
.B(n_1215),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1187),
.A2(n_1207),
.B(n_1204),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1181),
.A2(n_1139),
.B1(n_1185),
.B2(n_1172),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1187),
.A2(n_1207),
.B(n_1204),
.Y(n_1317)
);

AOI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1177),
.A2(n_979),
.B(n_1209),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1172),
.A2(n_1209),
.B(n_1185),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1129),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1188),
.B(n_878),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1199),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1199),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1172),
.A2(n_1209),
.B(n_1185),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1174),
.B(n_1192),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1187),
.A2(n_1207),
.B(n_1204),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1188),
.B(n_1185),
.C(n_1172),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1158),
.B(n_1032),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1106),
.A2(n_1102),
.B(n_1118),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1199),
.Y(n_1330)
);

CKINVDCx8_ASAP7_75t_R g1331 ( 
.A(n_1184),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1158),
.B(n_1032),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1251),
.B(n_1239),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1236),
.A2(n_1297),
.B(n_1216),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1251),
.B(n_1293),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1230),
.B(n_1261),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1288),
.B(n_1290),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1293),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1289),
.B(n_1328),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1241),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1229),
.A2(n_1312),
.B1(n_1295),
.B2(n_1245),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1320),
.B(n_1280),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1286),
.B(n_1220),
.Y(n_1343)
);

INVx3_ASAP7_75t_SL g1344 ( 
.A(n_1255),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1220),
.B(n_1226),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1226),
.B(n_1287),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1226),
.B(n_1287),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1320),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1328),
.B(n_1332),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1230),
.B(n_1261),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1271),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1303),
.B(n_1325),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1252),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1245),
.A2(n_1300),
.B1(n_1316),
.B2(n_1224),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1309),
.A2(n_1227),
.B(n_1318),
.C(n_1244),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1300),
.A2(n_1316),
.B1(n_1224),
.B2(n_1327),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1257),
.B(n_1276),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1255),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1262),
.A2(n_1321),
.B1(n_1250),
.B2(n_1301),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1309),
.B(n_1254),
.Y(n_1360)
);

AOI221xp5_ASAP7_75t_L g1361 ( 
.A1(n_1292),
.A2(n_1324),
.B1(n_1319),
.B2(n_1310),
.C(n_1321),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1274),
.Y(n_1362)
);

OA22x2_ASAP7_75t_L g1363 ( 
.A1(n_1266),
.A2(n_1257),
.B1(n_1284),
.B2(n_1332),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1328),
.B(n_1332),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1221),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1266),
.A2(n_1271),
.B1(n_1240),
.B2(n_1305),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1266),
.A2(n_1240),
.B1(n_1305),
.B2(n_1304),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1294),
.A2(n_1233),
.B(n_1314),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1223),
.A2(n_1314),
.B(n_1291),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1298),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1269),
.B(n_1264),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1222),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1232),
.A2(n_1247),
.B(n_1246),
.Y(n_1373)
);

NOR2xp67_ASAP7_75t_L g1374 ( 
.A(n_1243),
.B(n_1279),
.Y(n_1374)
);

O2A1O1Ixp5_ASAP7_75t_L g1375 ( 
.A1(n_1231),
.A2(n_1253),
.B(n_1242),
.C(n_1329),
.Y(n_1375)
);

INVx6_ASAP7_75t_SL g1376 ( 
.A(n_1267),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1217),
.B(n_1218),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1228),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1299),
.B(n_1302),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1264),
.B(n_1268),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1238),
.B(n_1235),
.Y(n_1381)
);

AOI211xp5_ASAP7_75t_L g1382 ( 
.A1(n_1273),
.A2(n_1249),
.B(n_1258),
.C(n_1259),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1307),
.B(n_1323),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1313),
.B(n_1322),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1298),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1256),
.A2(n_1248),
.B(n_1225),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1330),
.B(n_1277),
.Y(n_1387)
);

O2A1O1Ixp5_ASAP7_75t_L g1388 ( 
.A1(n_1281),
.A2(n_1275),
.B(n_1270),
.C(n_1278),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1263),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1304),
.A2(n_1331),
.B1(n_1233),
.B2(n_1311),
.Y(n_1390)
);

NOR3xp33_ASAP7_75t_L g1391 ( 
.A(n_1234),
.B(n_1308),
.C(n_1237),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_SL g1392 ( 
.A(n_1219),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1294),
.A2(n_1272),
.B(n_1285),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1311),
.A2(n_1234),
.B1(n_1308),
.B2(n_1237),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1282),
.B(n_1260),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1238),
.B(n_1235),
.Y(n_1396)
);

O2A1O1Ixp5_ASAP7_75t_L g1397 ( 
.A1(n_1281),
.A2(n_1278),
.B(n_1275),
.C(n_1265),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1219),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1399)
);

O2A1O1Ixp5_ASAP7_75t_L g1400 ( 
.A1(n_1296),
.A2(n_1306),
.B(n_1315),
.C(n_1317),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1326),
.A2(n_1188),
.B(n_979),
.C(n_1117),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1229),
.A2(n_878),
.B1(n_1312),
.B2(n_1295),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1236),
.A2(n_1297),
.B(n_1216),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1216),
.A2(n_1190),
.B(n_1297),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1289),
.B(n_1328),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1239),
.B(n_1288),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1230),
.B(n_1261),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1230),
.B(n_1261),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1251),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1251),
.B(n_1239),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1236),
.A2(n_758),
.B(n_997),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1230),
.B(n_1261),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1271),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1362),
.Y(n_1414)
);

OAI332xp33_ASAP7_75t_L g1415 ( 
.A1(n_1341),
.A2(n_1356),
.A3(n_1354),
.B1(n_1402),
.B2(n_1412),
.B3(n_1407),
.C1(n_1336),
.C2(n_1408),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1406),
.B(n_1337),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1395),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1350),
.B(n_1355),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1406),
.B(n_1337),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1338),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1361),
.A2(n_1359),
.B1(n_1355),
.B2(n_1366),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1400),
.A2(n_1334),
.B(n_1403),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1349),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1348),
.B(n_1353),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1388),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1349),
.B(n_1364),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1346),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1360),
.B(n_1365),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1399),
.B(n_1371),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1335),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1372),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1378),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1347),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1339),
.B(n_1405),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1347),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1371),
.B(n_1380),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1345),
.A2(n_1343),
.B(n_1396),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1399),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1381),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1389),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1397),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1387),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1380),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1396),
.B(n_1343),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1339),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1405),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1405),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1357),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1363),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1390),
.B(n_1401),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1352),
.B(n_1385),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1342),
.B(n_1363),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1421),
.A2(n_1333),
.B1(n_1410),
.B2(n_1376),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1421),
.A2(n_1367),
.B1(n_1409),
.B2(n_1382),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1448),
.B(n_1404),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1427),
.B(n_1433),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1414),
.Y(n_1458)
);

NAND2x1_ASAP7_75t_L g1459 ( 
.A(n_1436),
.B(n_1393),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1437),
.B(n_1404),
.Y(n_1460)
);

AOI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1415),
.A2(n_1411),
.B1(n_1375),
.B2(n_1340),
.C(n_1368),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1438),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1442),
.B(n_1384),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1431),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1437),
.B(n_1373),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1444),
.B(n_1383),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1429),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1432),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1444),
.B(n_1379),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1432),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1435),
.B(n_1386),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1452),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1428),
.B(n_1377),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1450),
.A2(n_1376),
.B1(n_1370),
.B2(n_1374),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1464),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1458),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1472),
.B(n_1416),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1461),
.A2(n_1450),
.B(n_1418),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1464),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1461),
.B(n_1452),
.C(n_1418),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1472),
.A2(n_1415),
.B1(n_1449),
.B2(n_1430),
.C(n_1428),
.Y(n_1481)
);

AOI222xp33_ASAP7_75t_L g1482 ( 
.A1(n_1474),
.A2(n_1449),
.B1(n_1451),
.B2(n_1430),
.C1(n_1351),
.C2(n_1413),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1457),
.B(n_1416),
.Y(n_1483)
);

AOI211xp5_ASAP7_75t_L g1484 ( 
.A1(n_1474),
.A2(n_1422),
.B(n_1420),
.C(n_1394),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1467),
.Y(n_1485)
);

AO21x1_ASAP7_75t_SL g1486 ( 
.A1(n_1455),
.A2(n_1446),
.B(n_1447),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1454),
.B(n_1453),
.C(n_1456),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1460),
.A2(n_1441),
.B(n_1425),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1459),
.B(n_1426),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1466),
.Y(n_1490)
);

AND4x1_ASAP7_75t_L g1491 ( 
.A(n_1454),
.B(n_1376),
.C(n_1391),
.D(n_1447),
.Y(n_1491)
);

INVx5_ASAP7_75t_L g1492 ( 
.A(n_1462),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1466),
.B(n_1469),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1457),
.B(n_1419),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1468),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1473),
.B(n_1446),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_R g1497 ( 
.A(n_1453),
.B(n_1358),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1459),
.A2(n_1369),
.B(n_1422),
.C(n_1370),
.Y(n_1498)
);

INVx4_ASAP7_75t_L g1499 ( 
.A(n_1467),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1456),
.A2(n_1441),
.B1(n_1425),
.B2(n_1440),
.C(n_1424),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1470),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1467),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1473),
.A2(n_1429),
.B1(n_1445),
.B2(n_1443),
.C(n_1417),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1467),
.B(n_1434),
.Y(n_1504)
);

AND2x2_ASAP7_75t_SL g1505 ( 
.A(n_1460),
.B(n_1423),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1434),
.Y(n_1506)
);

AOI211xp5_ASAP7_75t_L g1507 ( 
.A1(n_1460),
.A2(n_1422),
.B(n_1344),
.C(n_1443),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1463),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1475),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1479),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1505),
.B(n_1486),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1489),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1492),
.B(n_1462),
.Y(n_1513)
);

INVx8_ASAP7_75t_L g1514 ( 
.A(n_1489),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1500),
.B(n_1455),
.Y(n_1515)
);

AO21x1_ASAP7_75t_L g1516 ( 
.A1(n_1478),
.A2(n_1484),
.B(n_1507),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1488),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_SL g1518 ( 
.A(n_1482),
.B(n_1358),
.C(n_1465),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1492),
.B(n_1489),
.Y(n_1519)
);

INVx4_ASAP7_75t_SL g1520 ( 
.A(n_1489),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1490),
.B(n_1471),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1488),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1488),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1476),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1495),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1492),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1492),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1463),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1501),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1502),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1505),
.B(n_1506),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1511),
.B(n_1506),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1483),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1531),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1529),
.B(n_1496),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1524),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1511),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1531),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1529),
.B(n_1508),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1523),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1515),
.B(n_1508),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1523),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1515),
.B(n_1487),
.C(n_1481),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1519),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1533),
.B(n_1483),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1533),
.B(n_1494),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1504),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1524),
.B(n_1477),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_1493),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1533),
.B(n_1494),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1520),
.B(n_1504),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1523),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1509),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1532),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1510),
.B(n_1525),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1519),
.B(n_1485),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1521),
.B(n_1477),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1516),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1519),
.B(n_1485),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1519),
.B(n_1485),
.Y(n_1563)
);

NAND2xp67_ASAP7_75t_L g1564 ( 
.A(n_1527),
.B(n_1344),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1509),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1532),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_L g1567 ( 
.A(n_1514),
.B(n_1497),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1532),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1520),
.B(n_1504),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1518),
.A2(n_1498),
.B(n_1491),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1519),
.B(n_1499),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1521),
.B(n_1503),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1527),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1519),
.B(n_1499),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1556),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1545),
.B(n_1516),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1539),
.B(n_1520),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1561),
.B(n_1520),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1561),
.B(n_1526),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1561),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1551),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1539),
.B(n_1520),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1551),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1545),
.B(n_1516),
.Y(n_1586)
);

NAND4xp25_ASAP7_75t_L g1587 ( 
.A(n_1570),
.B(n_1518),
.C(n_1498),
.D(n_1512),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1565),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1565),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1570),
.B(n_1522),
.C(n_1517),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1535),
.B(n_1520),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1558),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1535),
.B(n_1512),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1543),
.A2(n_1526),
.B(n_1530),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1557),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1558),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1535),
.B(n_1512),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1566),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1536),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1542),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1536),
.Y(n_1601)
);

NOR2x1p5_ASAP7_75t_SL g1602 ( 
.A(n_1542),
.B(n_1523),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1542),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1540),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1538),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1544),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1540),
.Y(n_1608)
);

NAND3x2_ASAP7_75t_L g1609 ( 
.A(n_1572),
.B(n_1513),
.C(n_1497),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1547),
.B(n_1513),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1582),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1606),
.B(n_1538),
.Y(n_1612)
);

AOI22x1_ASAP7_75t_L g1613 ( 
.A1(n_1581),
.A2(n_1568),
.B1(n_1546),
.B2(n_1573),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1582),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1576),
.B(n_1537),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1586),
.A2(n_1567),
.B1(n_1543),
.B2(n_1537),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1584),
.Y(n_1618)
);

NAND4xp25_ASAP7_75t_L g1619 ( 
.A(n_1590),
.B(n_1541),
.C(n_1572),
.D(n_1568),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1595),
.B(n_1598),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1581),
.B(n_1546),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1578),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1591),
.B(n_1548),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1593),
.B(n_1548),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1578),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1584),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1585),
.B(n_1550),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1580),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1609),
.A2(n_1549),
.B1(n_1554),
.B2(n_1569),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1550),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1593),
.B(n_1548),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1579),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1597),
.B(n_1553),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1609),
.A2(n_1579),
.B1(n_1583),
.B2(n_1597),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1579),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1583),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1553),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1624),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1613),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1616),
.B(n_1583),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1614),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1628),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1612),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1612),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1625),
.B(n_1553),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1619),
.A2(n_1587),
.B(n_1594),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1635),
.B(n_1564),
.Y(n_1648)
);

O2A1O1Ixp5_ASAP7_75t_L g1649 ( 
.A1(n_1621),
.A2(n_1601),
.B(n_1608),
.C(n_1605),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1634),
.A2(n_1592),
.B1(n_1596),
.B2(n_1608),
.C(n_1605),
.Y(n_1650)
);

AOI322xp5_ASAP7_75t_L g1651 ( 
.A1(n_1617),
.A2(n_1637),
.A3(n_1633),
.B1(n_1631),
.B2(n_1621),
.C1(n_1636),
.C2(n_1623),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1631),
.Y(n_1652)
);

XOR2x2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.B(n_1601),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1632),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1613),
.A2(n_1549),
.B1(n_1554),
.B2(n_1569),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1629),
.A2(n_1620),
.B(n_1614),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1638),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1639),
.B(n_1623),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1652),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1647),
.A2(n_1627),
.B1(n_1622),
.B2(n_1546),
.C(n_1630),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1644),
.A2(n_1637),
.B1(n_1633),
.B2(n_1514),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1622),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1653),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1640),
.B(n_1575),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1645),
.B(n_1627),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1642),
.Y(n_1668)
);

AOI222xp33_ASAP7_75t_L g1669 ( 
.A1(n_1665),
.A2(n_1650),
.B1(n_1653),
.B2(n_1640),
.C1(n_1656),
.C2(n_1643),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1667),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1666),
.A2(n_1649),
.B(n_1651),
.C(n_1641),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1660),
.B(n_1639),
.Y(n_1672)
);

OAI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1662),
.A2(n_1641),
.B(n_1648),
.C(n_1642),
.Y(n_1673)
);

OAI322xp33_ASAP7_75t_L g1674 ( 
.A1(n_1659),
.A2(n_1657),
.A3(n_1646),
.B1(n_1618),
.B2(n_1626),
.C1(n_1615),
.C2(n_1630),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1661),
.B(n_1657),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1667),
.B(n_1592),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1673),
.B(n_1664),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1669),
.A2(n_1671),
.B(n_1672),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1670),
.A2(n_1663),
.B1(n_1655),
.B2(n_1577),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1668),
.B(n_1575),
.C(n_1596),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1668),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1681),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1680),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_L g1684 ( 
.A(n_1678),
.B(n_1675),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1677),
.B(n_1676),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1679),
.B(n_1610),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1681),
.B(n_1610),
.Y(n_1687)
);

AO22x2_ASAP7_75t_L g1688 ( 
.A1(n_1683),
.A2(n_1573),
.B1(n_1589),
.B2(n_1588),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1684),
.A2(n_1549),
.B1(n_1569),
.B2(n_1554),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1682),
.B(n_1534),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1685),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1687),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1691),
.B(n_1686),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1690),
.B(n_1588),
.Y(n_1694)
);

AOI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1689),
.A2(n_1674),
.B(n_1589),
.C(n_1559),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1693),
.A2(n_1692),
.B1(n_1688),
.B2(n_1607),
.Y(n_1696)
);

A2O1A1Ixp33_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1695),
.B(n_1694),
.C(n_1602),
.Y(n_1697)
);

OR3x2_ASAP7_75t_L g1698 ( 
.A(n_1697),
.B(n_1560),
.C(n_1552),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1697),
.A2(n_1607),
.B1(n_1604),
.B2(n_1600),
.C(n_1544),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1698),
.A2(n_1604),
.B1(n_1600),
.B2(n_1559),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1699),
.A2(n_1555),
.B1(n_1544),
.B2(n_1571),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_1700),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1701),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1702),
.A2(n_1392),
.B1(n_1398),
.B2(n_1554),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1703),
.Y(n_1705)
);

XNOR2xp5_ASAP7_75t_L g1706 ( 
.A(n_1705),
.B(n_1564),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1704),
.B(n_1555),
.Y(n_1707)
);

AOI322xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1555),
.A3(n_1574),
.B1(n_1571),
.B2(n_1559),
.C1(n_1562),
.C2(n_1563),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1562),
.B1(n_1574),
.B2(n_1571),
.C(n_1563),
.Y(n_1709)
);

AOI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1562),
.B(n_1574),
.C(n_1563),
.Y(n_1710)
);


endmodule