module fake_jpeg_7231_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_27),
.B1(n_33),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_72),
.B1(n_37),
.B2(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_37),
.B1(n_36),
.B2(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_28),
.B1(n_19),
.B2(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_88),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_78),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_84),
.B1(n_64),
.B2(n_52),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_14),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_97),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_99),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_17),
.B(n_20),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_52),
.B1(n_73),
.B2(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_48),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_107),
.B1(n_118),
.B2(n_124),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_0),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_0),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_94),
.B1(n_92),
.B2(n_97),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_53),
.B1(n_50),
.B2(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_127),
.Y(n_143)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_69),
.B1(n_21),
.B2(n_43),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_50),
.B1(n_69),
.B2(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_123),
.Y(n_145)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx5_ASAP7_75t_SL g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_43),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_21),
.B1(n_48),
.B2(n_43),
.Y(n_128)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_91),
.CON(n_130),
.SN(n_130)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_150),
.B(n_125),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_48),
.C(n_62),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_146),
.C(n_155),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_140),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_113),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_122),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_10),
.Y(n_149)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_34),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_95),
.B1(n_82),
.B2(n_89),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_112),
.B1(n_128),
.B2(n_114),
.Y(n_163)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_83),
.B1(n_123),
.B2(n_79),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_42),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_111),
.B1(n_115),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_171),
.B1(n_172),
.B2(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_109),
.B(n_127),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_166),
.B(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_184),
.B1(n_181),
.B2(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_178),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_0),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_150),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_119),
.B(n_104),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_95),
.B1(n_124),
.B2(n_96),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_95),
.B1(n_96),
.B2(n_83),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_63),
.C(n_62),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_136),
.C(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_182),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_83),
.B1(n_91),
.B2(n_79),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_199),
.C(n_202),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_169),
.B1(n_156),
.B2(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_209),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_208),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_135),
.B1(n_138),
.B2(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_145),
.C(n_129),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_171),
.C(n_166),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_145),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_144),
.B1(n_79),
.B2(n_91),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_144),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_210),
.Y(n_228)
);

OR2x4_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_38),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_170),
.B(n_194),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_31),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_63),
.C(n_134),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_157),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_231),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_183),
.B(n_182),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_192),
.B1(n_185),
.B2(n_191),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_232),
.B1(n_235),
.B2(n_214),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_193),
.B1(n_185),
.B2(n_196),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_190),
.B(n_161),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_236),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_184),
.B1(n_163),
.B2(n_170),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_193),
.B1(n_200),
.B2(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_29),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_180),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

XOR2x2_ASAP7_75t_SL g236 ( 
.A(n_190),
.B(n_167),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_211),
.C(n_209),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_189),
.B(n_157),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_24),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_240),
.A2(n_253),
.B1(n_259),
.B2(n_25),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_187),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_243),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_247),
.B1(n_261),
.B2(n_30),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_223),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_202),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_258),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_200),
.B1(n_201),
.B2(n_208),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_250),
.C(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_192),
.C(n_191),
.Y(n_250)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_223),
.C(n_225),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_137),
.C(n_174),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_260),
.C(n_67),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_75),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_234),
.B1(n_216),
.B2(n_236),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_102),
.C(n_75),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_24),
.B1(n_34),
.B2(n_25),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_226),
.C(n_213),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_31),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_230),
.B1(n_233),
.B2(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_228),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_245),
.A2(n_239),
.B1(n_252),
.B2(n_258),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_275),
.B1(n_277),
.B2(n_30),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_226),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_218),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

AO221x1_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_274),
.B1(n_18),
.B2(n_31),
.C(n_3),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_254),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_246),
.B1(n_260),
.B2(n_252),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_30),
.B1(n_31),
.B2(n_42),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_244),
.B1(n_67),
.B2(n_61),
.Y(n_282)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_279),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_295),
.B1(n_18),
.B2(n_35),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_61),
.B1(n_55),
.B2(n_93),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_289),
.B1(n_288),
.B2(n_280),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_277),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_291),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_278),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_61),
.B1(n_55),
.B2(n_93),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_55),
.B1(n_11),
.B2(n_12),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_293),
.Y(n_305)
);

AOI321xp33_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_38),
.A3(n_31),
.B1(n_18),
.B2(n_35),
.C(n_10),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_1),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_294),
.A2(n_263),
.B(n_265),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_263),
.C(n_278),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_15),
.C(n_13),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_307),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_272),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_290),
.B1(n_287),
.B2(n_3),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_16),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_10),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_298),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_15),
.B(n_13),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_306),
.B(n_305),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_1),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_309),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_296),
.B(n_303),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_324),
.A3(n_325),
.B1(n_326),
.B2(n_317),
.C1(n_2),
.C2(n_4),
.Y(n_330)
);

OA21x2_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_307),
.B(n_305),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_313),
.C(n_312),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_332),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_304),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_329),
.A2(n_330),
.B(n_327),
.C(n_5),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_331),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_4),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_334),
.B1(n_6),
.B2(n_8),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_4),
.C(n_6),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_8),
.C(n_9),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_9),
.Y(n_340)
);


endmodule