module fake_aes_1116_n_674 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_674);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_674;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_57), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_10), .Y(n_79) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_44), .B(n_45), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_13), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_74), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_56), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_21), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_76), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_29), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_41), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_54), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_15), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_13), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_75), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_51), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_61), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_20), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_62), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_23), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_40), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_28), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_25), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_55), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_33), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_31), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_71), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_27), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_64), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_43), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_26), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_52), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_10), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_14), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_73), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_38), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_7), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_101), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_101), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_81), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_101), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_79), .B(n_0), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_90), .B(n_34), .Y(n_138) );
INVx6_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_78), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_124), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_124), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_82), .B(n_1), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_92), .B(n_3), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_84), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_96), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_100), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_98), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_110), .B(n_4), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_108), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_109), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_114), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_117), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_148), .B(n_106), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_159), .B(n_118), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_148), .B(n_87), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_148), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_148), .B(n_106), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_140), .A2(n_123), .B1(n_78), .B2(n_119), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_129), .B(n_122), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_129), .B(n_121), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_131), .B(n_120), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_131), .B(n_112), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_159), .B(n_115), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
NAND3xp33_ASAP7_75t_L g190 ( .A(n_146), .B(n_112), .C(n_105), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_143), .B(n_133), .Y(n_191) );
NOR2x1p5_ASAP7_75t_L g192 ( .A(n_134), .B(n_104), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_143), .B(n_80), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_134), .B(n_86), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_155), .B(n_113), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_153), .B(n_165), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_145), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_165), .B(n_102), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_126), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_138), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
BUFx10_ASAP7_75t_L g206 ( .A(n_138), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
INVxp67_ASAP7_75t_SL g208 ( .A(n_157), .Y(n_208) );
NAND2x1p5_ASAP7_75t_L g209 ( .A(n_133), .B(n_91), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_149), .B(n_91), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_158), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_135), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
AND2x6_ASAP7_75t_L g214 ( .A(n_136), .B(n_89), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_126), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_127), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_136), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_130), .Y(n_218) );
AND2x6_ASAP7_75t_L g219 ( .A(n_142), .B(n_89), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_142), .B(n_36), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_149), .B(n_37), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_127), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_137), .B(n_5), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_151), .B(n_35), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_127), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_150), .B(n_42), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_189), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_195), .B(n_144), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_207), .Y(n_238) );
BUFx12f_ASAP7_75t_L g239 ( .A(n_211), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_186), .B(n_150), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_210), .B(n_167), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_178), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_206), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_226), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_202), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_208), .B(n_140), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_197), .B(n_167), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_191), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_195), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_196), .A2(n_151), .B1(n_164), .B2(n_156), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_177), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_183), .A2(n_138), .B1(n_164), .B2(n_162), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_195), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_170), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_170), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_196), .A2(n_162), .B1(n_156), .B2(n_138), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_170), .Y(n_259) );
BUFx2_ASAP7_75t_SL g260 ( .A(n_191), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_192), .B(n_191), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_196), .A2(n_138), .B1(n_154), .B2(n_150), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_202), .B(n_150), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_188), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_188), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_188), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_172), .B(n_163), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_168), .B(n_154), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_179), .A2(n_163), .B(n_161), .C(n_154), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_191), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_191), .A2(n_138), .B1(n_161), .B2(n_152), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_189), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_176), .B(n_166), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_212), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_191), .B(n_166), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_218), .B(n_166), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_201), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_213), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_199), .Y(n_280) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_195), .B(n_166), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_201), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_206), .B(n_166), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_199), .B(n_152), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_187), .B(n_152), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_217), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_227), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
NOR2x1_ASAP7_75t_L g290 ( .A(n_190), .B(n_132), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_214), .A2(n_132), .B1(n_128), .B2(n_127), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_214), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_204), .Y(n_294) );
AND2x4_ASAP7_75t_SL g295 ( .A(n_227), .B(n_132), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_209), .B(n_5), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_224), .B(n_128), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_187), .B(n_132), .Y(n_298) );
CKINVDCx6p67_ASAP7_75t_R g299 ( .A(n_239), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_287), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_252), .B(n_209), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_250), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_244), .B(n_227), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_260), .B(n_227), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_241), .A2(n_258), .B1(n_262), .B2(n_256), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_255), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_296), .A2(n_214), .B1(n_219), .B2(n_193), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_269), .A2(n_185), .B(n_181), .C(n_184), .Y(n_312) );
BUFx12f_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_270), .A2(n_185), .B1(n_184), .B2(n_181), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_241), .A2(n_219), .B1(n_214), .B2(n_193), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_276), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_237), .A2(n_173), .B1(n_219), .B2(n_214), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_245), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_289), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_293), .Y(n_321) );
NAND2xp33_ASAP7_75t_R g322 ( .A(n_251), .B(n_214), .Y(n_322) );
AND2x6_ASAP7_75t_L g323 ( .A(n_293), .B(n_228), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_233), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_240), .A2(n_173), .B(n_221), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_261), .A2(n_219), .B1(n_193), .B2(n_222), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_281), .B(n_221), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_238), .Y(n_328) );
INVx5_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_249), .B(n_219), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_236), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_236), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_276), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_232), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_242), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_254), .A2(n_219), .B(n_193), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_253), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_267), .A2(n_194), .B(n_198), .C(n_231), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_272), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_235), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_257), .B(n_193), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_240), .A2(n_204), .B(n_198), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_237), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_237), .A2(n_193), .B1(n_231), .B2(n_220), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_263), .A2(n_194), .B(n_198), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_280), .B(n_6), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_232), .B(n_194), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_261), .B(n_285), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_320), .Y(n_350) );
AND2x2_ASAP7_75t_SL g351 ( .A(n_319), .B(n_295), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_309), .A2(n_295), .B1(n_271), .B2(n_288), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_331), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_303), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_318), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_300), .B(n_261), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_309), .A2(n_271), .B1(n_254), .B2(n_264), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_338), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_303), .B(n_259), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_300), .A2(n_266), .B1(n_265), .B2(n_267), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_307), .A2(n_248), .B1(n_277), .B2(n_286), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_304), .B(n_268), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_329), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_306), .A2(n_290), .B1(n_263), .B2(n_234), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_301), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_301), .B(n_234), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_302), .B(n_246), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_306), .Y(n_373) );
BUFx4_ASAP7_75t_SL g374 ( .A(n_344), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_307), .A2(n_298), .B1(n_274), .B2(n_291), .Y(n_377) );
AOI21xp5_ASAP7_75t_SL g378 ( .A1(n_337), .A2(n_246), .B(n_273), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_308), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_302), .A2(n_274), .B1(n_298), .B2(n_291), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_364), .A2(n_344), .B1(n_307), .B2(n_315), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_356), .A2(n_310), .B1(n_341), .B2(n_307), .Y(n_382) );
OAI33xp33_ASAP7_75t_L g383 ( .A1(n_364), .A2(n_347), .A3(n_345), .B1(n_341), .B2(n_330), .B3(n_312), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_373), .A2(n_347), .B1(n_315), .B2(n_349), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_365), .A2(n_324), .B1(n_328), .B2(n_311), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_373), .A2(n_349), .B1(n_324), .B2(n_328), .C(n_314), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_356), .B(n_319), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_362), .A2(n_360), .B1(n_363), .B2(n_354), .C(n_350), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_350), .B(n_342), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_377), .A2(n_325), .B(n_327), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_353), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_370), .B(n_336), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_374), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_370), .B(n_316), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_326), .B(n_317), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_352), .A2(n_310), .B1(n_351), .B2(n_313), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_365), .A2(n_352), .B1(n_354), .B2(n_360), .C(n_363), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_365), .A2(n_299), .B1(n_322), .B2(n_319), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_357), .B(n_299), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_361), .A2(n_334), .B1(n_316), .B2(n_336), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_351), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_378), .A2(n_339), .B(n_284), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_357), .B(n_316), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_351), .A2(n_305), .B1(n_329), .B2(n_334), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_361), .A2(n_329), .B1(n_305), .B2(n_323), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
AOI22xp5_ASAP7_75t_SL g409 ( .A1(n_394), .A2(n_374), .B1(n_377), .B2(n_366), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_404), .A2(n_368), .B(n_376), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_359), .B1(n_357), .B2(n_371), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_393), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_397), .A2(n_361), .B1(n_359), .B2(n_366), .Y(n_414) );
OAI222xp33_ASAP7_75t_L g415 ( .A1(n_381), .A2(n_366), .B1(n_376), .B2(n_375), .C1(n_368), .C2(n_355), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_396), .A2(n_361), .B1(n_371), .B2(n_372), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_390), .B(n_402), .Y(n_417) );
OA21x2_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_380), .B(n_376), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_396), .A2(n_361), .B1(n_372), .B2(n_371), .Y(n_419) );
AO21x2_ASAP7_75t_L g420 ( .A1(n_391), .A2(n_375), .B(n_292), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_402), .B(n_375), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_383), .A2(n_372), .B1(n_367), .B2(n_379), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_392), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_393), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_398), .A2(n_379), .B1(n_329), .B2(n_369), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_388), .B(n_379), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_385), .A2(n_380), .B1(n_379), .B2(n_346), .C(n_284), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_386), .B(n_127), .C(n_128), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_392), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_403), .A2(n_369), .B1(n_355), .B2(n_358), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_408), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_408), .B(n_358), .Y(n_432) );
AOI31xp67_ASAP7_75t_L g433 ( .A1(n_389), .A2(n_225), .A3(n_216), .B(n_215), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_384), .A2(n_355), .B1(n_329), .B2(n_335), .C(n_358), .Y(n_434) );
AOI21xp5_ASAP7_75t_SL g435 ( .A1(n_385), .A2(n_358), .B(n_321), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_395), .B(n_358), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_399), .A2(n_291), .B1(n_284), .B2(n_231), .C(n_220), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_382), .B(n_358), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_400), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_407), .A2(n_355), .B1(n_358), .B2(n_333), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_405), .B(n_333), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_431), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_423), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_417), .B(n_405), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_431), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_412), .B(n_387), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_417), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_412), .B(n_401), .Y(n_452) );
OAI31xp33_ASAP7_75t_L g453 ( .A1(n_415), .A2(n_340), .A3(n_348), .B(n_308), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_428), .A2(n_406), .B(n_340), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_442), .B(n_369), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_414), .A2(n_335), .B1(n_348), .B2(n_308), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_429), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_437), .B(n_6), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_421), .B(n_8), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_437), .B(n_8), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_440), .B(n_9), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_437), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_432), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_438), .B(n_60), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_432), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_424), .B(n_9), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_440), .B(n_11), .Y(n_470) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_428), .A2(n_343), .B(n_297), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_409), .A2(n_323), .B1(n_291), .B2(n_284), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_409), .B(n_220), .C(n_180), .D(n_175), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_411), .B(n_11), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_418), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_425), .A2(n_335), .B1(n_348), .B2(n_321), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
NOR3xp33_ASAP7_75t_SL g479 ( .A(n_441), .B(n_297), .C(n_283), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_444), .B(n_12), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_418), .Y(n_481) );
OAI322xp33_ASAP7_75t_L g482 ( .A1(n_411), .A2(n_132), .A3(n_128), .B1(n_18), .B2(n_19), .C1(n_16), .C2(n_17), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_418), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_416), .B(n_16), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_436), .Y(n_486) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_422), .A2(n_171), .B1(n_174), .B2(n_175), .C(n_180), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_433), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_426), .B(n_17), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_426), .B(n_419), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_410), .B(n_420), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_435), .B(n_18), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_434), .B(n_19), .Y(n_494) );
NOR2xp67_ASAP7_75t_L g495 ( .A(n_434), .B(n_22), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_430), .B(n_171), .C(n_174), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_465), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_446), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_495), .B(n_443), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_493), .B(n_128), .C(n_439), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_457), .B(n_435), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_451), .B(n_443), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_495), .B(n_427), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_446), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_484), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_449), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_466), .B(n_420), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_480), .B(n_420), .Y(n_509) );
AOI31xp33_ASAP7_75t_L g510 ( .A1(n_472), .A2(n_433), .A3(n_30), .B(n_32), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_473), .B(n_24), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_480), .B(n_323), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_447), .B(n_46), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_460), .B(n_323), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_458), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_464), .B(n_49), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_466), .B(n_468), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_468), .B(n_50), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_458), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_464), .B(n_461), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_447), .B(n_53), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_469), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g524 ( .A1(n_493), .A2(n_58), .B(n_59), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_460), .B(n_63), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_445), .Y(n_526) );
OAI31xp33_ASAP7_75t_L g527 ( .A1(n_494), .A2(n_283), .A3(n_216), .B(n_225), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_462), .B(n_323), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_448), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_448), .B(n_65), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_475), .A2(n_494), .B(n_491), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_486), .B(n_229), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g534 ( .A(n_455), .B(n_67), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_467), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_462), .B(n_323), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_486), .B(n_69), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_490), .B(n_70), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_490), .B(n_72), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_482), .B(n_294), .C(n_282), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_475), .B(n_169), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_481), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_452), .B(n_169), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_452), .B(n_169), .Y(n_544) );
AOI31xp33_ASAP7_75t_L g545 ( .A1(n_485), .A2(n_459), .A3(n_467), .B(n_470), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_453), .A2(n_273), .B(n_243), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_483), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_489), .Y(n_548) );
INVxp33_ASAP7_75t_SL g549 ( .A(n_485), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_463), .B(n_169), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_506), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_548), .B(n_492), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_532), .B(n_476), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_535), .B(n_467), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_545), .A2(n_459), .B1(n_474), .B2(n_450), .Y(n_556) );
NOR3xp33_ASAP7_75t_SL g557 ( .A(n_524), .B(n_482), .C(n_453), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_548), .Y(n_558) );
AND4x1_ASAP7_75t_L g559 ( .A(n_500), .B(n_479), .C(n_454), .D(n_496), .Y(n_559) );
NOR2xp67_ASAP7_75t_SL g560 ( .A(n_525), .B(n_487), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_517), .B(n_478), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_520), .Y(n_562) );
XNOR2xp5_ASAP7_75t_L g563 ( .A(n_549), .B(n_456), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_498), .B(n_483), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_522), .B(n_492), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_504), .B(n_492), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_549), .A2(n_531), .B1(n_523), .B2(n_534), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_507), .B(n_488), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_501), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_520), .B(n_515), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_537), .B(n_471), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_520), .B(n_477), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_519), .B(n_471), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_533), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_512), .A2(n_471), .B1(n_200), .B2(n_205), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_508), .B(n_182), .Y(n_577) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_537), .B(n_243), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_503), .B(n_182), .C(n_200), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_508), .B(n_200), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_509), .B(n_200), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_533), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_502), .B(n_205), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_516), .B(n_243), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_526), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_510), .A2(n_205), .B(n_229), .C(n_294), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_529), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_205), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_529), .B(n_229), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_542), .B(n_229), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_533), .B(n_278), .Y(n_591) );
NOR3xp33_ASAP7_75t_SL g592 ( .A(n_503), .B(n_278), .C(n_282), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_556), .A2(n_499), .B1(n_538), .B2(n_539), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_552), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_568), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_554), .Y(n_597) );
AO211x2_ASAP7_75t_L g598 ( .A1(n_579), .A2(n_536), .B(n_528), .C(n_541), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_570), .B(n_533), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_570), .B(n_542), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_558), .B(n_511), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
OAI32xp33_ASAP7_75t_L g603 ( .A1(n_575), .A2(n_521), .A3(n_513), .B1(n_499), .B2(n_518), .Y(n_603) );
OAI211xp5_ASAP7_75t_L g604 ( .A1(n_567), .A2(n_527), .B(n_544), .C(n_550), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_571), .B(n_547), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_561), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
AOI311xp33_ASAP7_75t_L g608 ( .A1(n_566), .A2(n_540), .A3(n_546), .B(n_543), .C(n_516), .Y(n_608) );
XOR2x2_ASAP7_75t_L g609 ( .A(n_563), .B(n_516), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_566), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_530), .B(n_518), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_553), .Y(n_612) );
XOR2xp5_ASAP7_75t_L g613 ( .A(n_555), .B(n_543), .Y(n_613) );
OAI322xp33_ASAP7_75t_L g614 ( .A1(n_573), .A2(n_243), .A3(n_247), .B1(n_575), .B2(n_564), .C1(n_572), .C2(n_569), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_591), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_564), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_592), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_569), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_SL g619 ( .A1(n_582), .A2(n_247), .B(n_557), .C(n_585), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_581), .A2(n_247), .B(n_577), .C(n_578), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_582), .A2(n_247), .B(n_584), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_572), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_581), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_583), .B(n_580), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_584), .A2(n_578), .B(n_574), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_560), .A2(n_588), .B1(n_580), .B2(n_577), .Y(n_627) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_574), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_590), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_589), .B(n_576), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_589), .B(n_559), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_565), .B(n_570), .Y(n_632) );
A2O1A1O1Ixp25_ASAP7_75t_L g633 ( .A1(n_552), .A2(n_545), .B(n_531), .C(n_455), .D(n_522), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_552), .B(n_565), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_566), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_556), .B(n_535), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_556), .A2(n_531), .A3(n_557), .B1(n_523), .B2(n_522), .C1(n_570), .C2(n_552), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_552), .B(n_565), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_563), .B(n_394), .Y(n_639) );
NOR2x1p5_ASAP7_75t_L g640 ( .A(n_617), .B(n_633), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_635), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_636), .A2(n_619), .B(n_594), .C(n_631), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_612), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g644 ( .A(n_637), .B(n_608), .C(n_593), .D(n_627), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_614), .B(n_619), .C(n_631), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_635), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_628), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_610), .B(n_602), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_609), .A2(n_639), .B(n_622), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_609), .A2(n_603), .B(n_639), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_597), .Y(n_651) );
NOR4xp25_ASAP7_75t_L g652 ( .A(n_595), .B(n_604), .C(n_607), .D(n_621), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_612), .A2(n_623), .B1(n_599), .B2(n_617), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_652), .A2(n_601), .B(n_615), .C(n_623), .Y(n_654) );
AOI221x1_ASAP7_75t_L g655 ( .A1(n_650), .A2(n_596), .B1(n_601), .B2(n_626), .C(n_618), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_649), .A2(n_611), .B1(n_606), .B2(n_613), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_651), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_644), .A2(n_630), .B(n_624), .C(n_625), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_647), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_648), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_640), .A2(n_638), .B(n_634), .C(n_616), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_658), .B(n_642), .C(n_645), .D(n_653), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_656), .A2(n_645), .B(n_647), .C(n_643), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_657), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_663), .A2(n_656), .B1(n_654), .B2(n_660), .Y(n_666) );
INVx4_ASAP7_75t_L g667 ( .A(n_662), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_664), .A2(n_661), .B1(n_655), .B2(n_646), .C(n_641), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_667), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_666), .Y(n_670) );
XOR2x2_ASAP7_75t_L g671 ( .A(n_669), .B(n_668), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_670), .B1(n_665), .B2(n_632), .C1(n_624), .C2(n_600), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_620), .B1(n_629), .B2(n_605), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_673), .A2(n_598), .B(n_632), .Y(n_674) );
endmodule