module real_jpeg_28061_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_4;
wire n_8;
wire n_6;
wire n_7;
wire n_9;

HAxp5_ASAP7_75t_SL g6 ( 
.A(n_0),
.B(n_7),
.CON(n_6),
.SN(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_SL g8 ( 
.A(n_2),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g3 ( 
.A1(n_4),
.A2(n_8),
.B(n_9),
.Y(n_3)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g4 ( 
.A(n_5),
.Y(n_4)
);

CKINVDCx5p33_ASAP7_75t_R g5 ( 
.A(n_6),
.Y(n_5)
);

BUFx24_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);


endmodule