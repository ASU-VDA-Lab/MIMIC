module real_jpeg_25289_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_206;
wire n_53;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_123),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_110),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_28),
.B(n_43),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_89),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_1),
.A2(n_25),
.B1(n_221),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_1),
.A2(n_64),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_2),
.A2(n_73),
.B1(n_74),
.B2(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_2),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_121),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_121),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_121),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_69),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_76),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_76),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_76),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_6),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_7),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_87),
.B1(n_107),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_87),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_8),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_9),
.A2(n_40),
.B1(n_64),
.B2(n_65),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_11),
.B(n_110),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_13),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_14),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_78),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_78),
.Y(n_241)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_149),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_148),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_20),
.B(n_125),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_21),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_21),
.B(n_153),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_92),
.CI(n_101),
.CON(n_21),
.SN(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_56),
.B1(n_57),
.B2(n_91),
.Y(n_22)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_24),
.B(n_41),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_25),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_25),
.A2(n_95),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_25),
.A2(n_211),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_25),
.A2(n_35),
.B(n_129),
.Y(n_247)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_26),
.B(n_39),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_33),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_26),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_27),
.B(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_31),
.B(n_110),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_51),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_42),
.A2(n_46),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_42),
.B(n_53),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_42),
.A2(n_99),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_42),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_42),
.B(n_110),
.Y(n_219)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_45),
.A2(n_48),
.B(n_110),
.C(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_48),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_47),
.B(n_84),
.Y(n_246)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_48),
.A2(n_64),
.A3(n_83),
.B1(n_239),
.B2(n_246),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_54),
.A2(n_133),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_54),
.A2(n_194),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_54),
.A2(n_202),
.B1(n_203),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_79),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_58),
.B(n_79),
.C(n_91),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_72),
.B2(n_77),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_59),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_59),
.A2(n_77),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_65),
.A3(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_106)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_65),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_65),
.B(n_110),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_73),
.A2(n_109),
.B(n_110),
.Y(n_161)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_88),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_80),
.A2(n_82),
.B1(n_178),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_81),
.B(n_90),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_81),
.A2(n_89),
.B1(n_103),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_81),
.A2(n_89),
.B1(n_163),
.B2(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_86),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_82),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_94),
.A2(n_115),
.B(n_128),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_100),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_99),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_119),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_119),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_112),
.B1(n_113),
.B2(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_106),
.Y(n_173)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_141),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_125),
.Y(n_276)
);

FAx1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.CI(n_147),
.CON(n_125),
.SN(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_146),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_183),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_165),
.B(n_182),
.Y(n_151)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_152),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_164),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_164),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_159),
.B(n_202),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_170),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_176),
.B(n_256),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_179),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_273),
.C(n_274),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_267),
.B(n_272),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_251),
.B(n_266),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_232),
.B(n_250),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_207),
.B(n_231),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_197),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_191),
.B1(n_195),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_205),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_204),
.C(n_205),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_217),
.B(n_230),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_215),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_224),
.B(n_229),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_243),
.C(n_248),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_261),
.C(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);


endmodule