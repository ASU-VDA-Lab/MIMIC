module fake_ariane_3077_n_2063 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2063);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2063;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_13),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_54),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_15),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_10),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_107),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_65),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_153),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_23),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_55),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_55),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g221 ( 
.A(n_173),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_101),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_54),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_48),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_75),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_10),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_85),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_90),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_178),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_72),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_25),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_88),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_191),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_56),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_166),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_24),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_130),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_49),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_78),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_161),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_143),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_113),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_137),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_116),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_32),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_75),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_122),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_8),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_156),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_157),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_115),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_32),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_27),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_169),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_92),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_182),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_105),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_22),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_163),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_95),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_91),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_60),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_56),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_114),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_16),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_74),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_58),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_41),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_62),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_20),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_0),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_82),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_134),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_96),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_72),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_69),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_118),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_13),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_66),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_62),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_21),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_41),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_109),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_20),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_36),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_14),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_87),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_43),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_168),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_144),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_9),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_37),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_138),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_76),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_40),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_18),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_18),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_172),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_27),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_9),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_65),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_16),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_7),
.Y(n_324)
);

BUFx8_ASAP7_75t_SL g325 ( 
.A(n_48),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_184),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_76),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_59),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_8),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_37),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_25),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_181),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_57),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_61),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_73),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_148),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_34),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_149),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_188),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_33),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_170),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_57),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_69),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_0),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_35),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_93),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_14),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_33),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_131),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_71),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_176),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_187),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_51),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_71),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_49),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_174),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_35),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_193),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_102),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_50),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_1),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_141),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_58),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_45),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_68),
.Y(n_367)
);

BUFx8_ASAP7_75t_SL g368 ( 
.A(n_19),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_40),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_6),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_70),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_36),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_164),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_97),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_31),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_127),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_31),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_125),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_64),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_11),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_145),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_81),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_190),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_132),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_89),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_64),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_51),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_42),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_68),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_60),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_42),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_77),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_290),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_325),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_368),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_197),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_252),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_249),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_280),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_272),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_198),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_232),
.Y(n_413)
);

INVxp33_ASAP7_75t_SL g414 ( 
.A(n_389),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_198),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_208),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_238),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_272),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_204),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_270),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_204),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_209),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_214),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_206),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_201),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_206),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_317),
.B(n_1),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_217),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_228),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_199),
.B(n_2),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_207),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_282),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_238),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_317),
.B(n_3),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_197),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_201),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_258),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_287),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_199),
.B(n_3),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_301),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_258),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_230),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_207),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_231),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_212),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_212),
.B(n_4),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_215),
.B(n_4),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_223),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_288),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_331),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_236),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_211),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_223),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_241),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_238),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_238),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_224),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_242),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_R g459 ( 
.A(n_202),
.B(n_80),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_238),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_356),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_247),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_257),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_224),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_235),
.B(n_5),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_259),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_235),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_248),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_211),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_272),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_262),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_374),
.Y(n_472)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_268),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_248),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_374),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_216),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_329),
.B(n_5),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_269),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_274),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_274),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_291),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_216),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_275),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_277),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_275),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_297),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_374),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_302),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_303),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_278),
.B(n_6),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_307),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_278),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_411),
.B(n_415),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_408),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_403),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_436),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_394),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_393),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_413),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_473),
.B(n_281),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_398),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_420),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_395),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_432),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_416),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_411),
.B(n_281),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_417),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_422),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_438),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_415),
.B(n_286),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_440),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_450),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_461),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_419),
.B(n_288),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_423),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_401),
.A2(n_293),
.B(n_286),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_418),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_428),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_429),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_455),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_442),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_418),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_414),
.A2(n_309),
.B1(n_285),
.B2(n_260),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_444),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_R g538 ( 
.A(n_409),
.B(n_451),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_407),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_470),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_455),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_419),
.B(n_293),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_370),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_402),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_454),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_421),
.B(n_370),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_456),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_458),
.B(n_392),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_404),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_R g553 ( 
.A(n_462),
.B(n_203),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_404),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_463),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_430),
.B(n_291),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_466),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_471),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_421),
.B(n_294),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_410),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_410),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_472),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_424),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_478),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_503),
.B(n_426),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_498),
.B(n_484),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_571),
.B(n_430),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_508),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_546),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_439),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_511),
.B(n_412),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_499),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_486),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_426),
.Y(n_586)
);

INVx8_ASAP7_75t_L g587 ( 
.A(n_559),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_529),
.B(n_431),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_551),
.B(n_488),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_499),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_501),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_570),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_507),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_570),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_559),
.B(n_396),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_529),
.B(n_431),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_546),
.B(n_443),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_553),
.B(n_489),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_493),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_559),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_527),
.B(n_482),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_507),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_507),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_495),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_495),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_502),
.B(n_443),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_538),
.B(n_491),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_517),
.B(n_427),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_493),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_559),
.A2(n_465),
.B1(n_490),
.B2(n_412),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_506),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_528),
.B(n_427),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_504),
.B(n_445),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_506),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_504),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_531),
.B(n_434),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_519),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_519),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_539),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_539),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_559),
.A2(n_434),
.B1(n_446),
.B2(n_445),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_527),
.B(n_396),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_544),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_549),
.B(n_435),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_544),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_549),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_532),
.B(n_446),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_548),
.B(n_447),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_547),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_547),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_527),
.B(n_435),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_521),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_552),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_554),
.B(n_448),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_534),
.B(n_447),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_554),
.B(n_448),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_556),
.B(n_453),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_506),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_549),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_549),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_506),
.Y(n_648)
);

AND2x2_ASAP7_75t_SL g649 ( 
.A(n_548),
.B(n_265),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_536),
.A2(n_457),
.B1(n_464),
.B2(n_453),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_514),
.B(n_452),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_513),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_514),
.B(n_452),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_565),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_513),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_497),
.B(n_425),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_513),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_565),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_567),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_567),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_520),
.B(n_294),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_537),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_524),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_524),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_524),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_555),
.A2(n_477),
.B1(n_469),
.B2(n_312),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_533),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_521),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_543),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_497),
.B(n_469),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_560),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_513),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_520),
.B(n_457),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_562),
.B(n_477),
.Y(n_678)
);

NAND2x1p5_ASAP7_75t_L g679 ( 
.A(n_529),
.B(n_464),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_545),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_545),
.B(n_467),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_513),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_505),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_425),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_543),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_564),
.B(n_467),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_515),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_516),
.B(n_468),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_572),
.B(n_494),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_543),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_550),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_550),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_516),
.B(n_468),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_515),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_516),
.B(n_474),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_515),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_561),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_561),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_561),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_510),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_566),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_R g704 ( 
.A(n_496),
.B(n_437),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_515),
.Y(n_705)
);

AND2x2_ASAP7_75t_SL g706 ( 
.A(n_515),
.B(n_265),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_511),
.B(n_437),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_566),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_530),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_566),
.Y(n_710)
);

NOR2x1p5_ASAP7_75t_L g711 ( 
.A(n_500),
.B(n_299),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_540),
.A2(n_345),
.B1(n_313),
.B2(n_315),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_515),
.B(n_339),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_569),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_522),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_522),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_569),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_569),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_540),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_522),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_516),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_522),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_558),
.B(n_474),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_558),
.Y(n_724)
);

INVx4_ASAP7_75t_SL g725 ( 
.A(n_522),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_585),
.B(n_535),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_649),
.B(n_339),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_649),
.A2(n_536),
.B1(n_487),
.B2(n_475),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_719),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_680),
.B(n_479),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_602),
.B(n_479),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_614),
.B(n_480),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_651),
.B(n_480),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_573),
.A2(n_375),
.B1(n_343),
.B2(n_349),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_649),
.B(n_518),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_598),
.B(n_483),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_587),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_598),
.A2(n_459),
.B1(n_376),
.B2(n_361),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_651),
.B(n_483),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_603),
.B(n_341),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_655),
.B(n_598),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_603),
.B(n_341),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_603),
.B(n_598),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_613),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_655),
.B(n_485),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_578),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_677),
.B(n_485),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_576),
.A2(n_348),
.B1(n_376),
.B2(n_361),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_681),
.B(n_492),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_686),
.B(n_492),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_593),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_578),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_719),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_713),
.A2(n_359),
.B1(n_306),
.B2(n_321),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_576),
.A2(n_383),
.B1(n_358),
.B2(n_353),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_632),
.B(n_523),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_620),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_684),
.B(n_558),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_584),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_620),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_576),
.B(n_245),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_684),
.B(n_558),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_622),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_684),
.B(n_441),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_684),
.B(n_441),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_622),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_L g767 ( 
.A(n_576),
.B(n_245),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_591),
.B(n_509),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_580),
.B(n_336),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_626),
.A2(n_324),
.B1(n_318),
.B2(n_316),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_594),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_607),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_702),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_580),
.B(n_449),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_604),
.B(n_481),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_SL g777 ( 
.A1(n_633),
.A2(n_481),
.B1(n_350),
.B2(n_391),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_587),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_576),
.A2(n_587),
.B1(n_629),
.B2(n_674),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_629),
.B(n_359),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_607),
.Y(n_781)
);

NOR2x2_ASAP7_75t_L g782 ( 
.A(n_633),
.B(n_525),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_604),
.B(n_226),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_629),
.B(n_346),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_623),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_631),
.B(n_526),
.Y(n_786)
);

INVxp33_ASAP7_75t_L g787 ( 
.A(n_658),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_629),
.B(n_627),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_576),
.B(n_346),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_638),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_615),
.B(n_340),
.C(n_328),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_627),
.B(n_226),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_608),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_719),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_623),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_608),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_583),
.B(n_542),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_583),
.B(n_707),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_576),
.B(n_600),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_713),
.A2(n_200),
.B1(n_321),
.B2(n_306),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_575),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_719),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_631),
.B(n_568),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_713),
.A2(n_200),
.B1(n_306),
.B2(n_321),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_638),
.B(n_229),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_630),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_663),
.A2(n_200),
.B1(n_245),
.B2(n_283),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_631),
.B(n_357),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_630),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_637),
.B(n_229),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_672),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_674),
.B(n_353),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_624),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_594),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_674),
.B(n_260),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_633),
.B(n_289),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_587),
.A2(n_358),
.B1(n_383),
.B2(n_253),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_707),
.B(n_672),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_663),
.A2(n_245),
.B1(n_283),
.B2(n_253),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_597),
.B(n_255),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_624),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_683),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_SL g824 ( 
.A1(n_587),
.A2(n_292),
.B1(n_334),
.B2(n_388),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_663),
.A2(n_245),
.B1(n_283),
.B2(n_221),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_625),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_646),
.A2(n_365),
.B1(n_390),
.B2(n_363),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_636),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_674),
.B(n_590),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_646),
.B(n_289),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_647),
.B(n_292),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_636),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_591),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_597),
.B(n_273),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_SL g835 ( 
.A1(n_633),
.A2(n_337),
.B1(n_335),
.B2(n_342),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_601),
.B(n_367),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_633),
.B(n_372),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_668),
.B(n_377),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_645),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_647),
.A2(n_326),
.B1(n_221),
.B2(n_311),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_597),
.B(n_254),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_581),
.B(n_296),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_707),
.B(n_296),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_711),
.B(n_300),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_594),
.B(n_254),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_581),
.B(n_300),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_591),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_645),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_581),
.A2(n_234),
.B1(n_244),
.B2(n_243),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_581),
.B(n_305),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_581),
.B(n_305),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_581),
.A2(n_227),
.B1(n_237),
.B2(n_233),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_707),
.B(n_379),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_581),
.A2(n_222),
.B1(n_239),
.B2(n_220),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_SL g855 ( 
.A1(n_625),
.A2(n_344),
.B(n_320),
.C(n_327),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_711),
.B(n_320),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_611),
.B(n_386),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_653),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_594),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_653),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_690),
.B(n_330),
.C(n_323),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_661),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_586),
.B(n_327),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_661),
.Y(n_864)
);

NOR2x2_ASAP7_75t_L g865 ( 
.A(n_591),
.B(n_7),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_628),
.B(n_254),
.Y(n_866)
);

INVx8_ASAP7_75t_L g867 ( 
.A(n_663),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_709),
.B(n_334),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_709),
.B(n_610),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_706),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_706),
.A2(n_213),
.B1(n_210),
.B2(n_218),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_628),
.B(n_254),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_634),
.B(n_335),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_698),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_588),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_634),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_617),
.B(n_263),
.Y(n_877)
);

AND3x2_ASAP7_75t_L g878 ( 
.A(n_664),
.B(n_362),
.C(n_337),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_664),
.Y(n_879)
);

O2A1O1Ixp5_ASAP7_75t_L g880 ( 
.A1(n_662),
.A2(n_352),
.B(n_366),
.C(n_342),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_635),
.B(n_344),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_621),
.B(n_322),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_635),
.B(n_639),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_639),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_650),
.B(n_352),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_666),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_L g887 ( 
.A(n_712),
.B(n_371),
.C(n_355),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_654),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_654),
.B(n_355),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_656),
.B(n_362),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_664),
.B(n_366),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_656),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_664),
.B(n_371),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_660),
.B(n_380),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_875),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_744),
.Y(n_896)
);

BUFx4f_ASAP7_75t_L g897 ( 
.A(n_774),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_SL g898 ( 
.A(n_726),
.B(n_678),
.C(n_641),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_R g899 ( 
.A(n_802),
.B(n_675),
.Y(n_899)
);

AND3x1_ASAP7_75t_SL g900 ( 
.A(n_787),
.B(n_387),
.C(n_380),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_746),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_802),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_736),
.B(n_788),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_757),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_736),
.B(n_609),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_737),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_790),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_760),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_751),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_736),
.B(n_618),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_823),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_788),
.B(n_640),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_737),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_746),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_883),
.A2(n_660),
.B(n_577),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_819),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_833),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_799),
.B(n_776),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_798),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_727),
.A2(n_675),
.B1(n_663),
.B2(n_706),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_737),
.B(n_778),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_727),
.A2(n_675),
.B1(n_663),
.B2(n_643),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_763),
.Y(n_923)
);

AND2x2_ASAP7_75t_SL g924 ( 
.A(n_761),
.B(n_612),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_798),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_778),
.Y(n_926)
);

AND2x6_ASAP7_75t_L g927 ( 
.A(n_779),
.B(n_612),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_741),
.B(n_642),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_778),
.B(n_725),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_875),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_766),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_785),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_812),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_875),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_768),
.Y(n_935)
);

AND2x6_ASAP7_75t_L g936 ( 
.A(n_817),
.B(n_592),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_875),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_752),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_752),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_796),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_733),
.B(n_663),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_800),
.A2(n_577),
.B(n_574),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_R g943 ( 
.A(n_833),
.B(n_675),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_885),
.A2(n_606),
.B1(n_605),
.B2(n_595),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_869),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_829),
.A2(n_574),
.B1(n_579),
.B2(n_582),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_761),
.A2(n_767),
.B1(n_838),
.B2(n_738),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_767),
.A2(n_579),
.B1(n_582),
.B2(n_721),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_772),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_776),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_869),
.Y(n_951)
);

CKINVDCx16_ASAP7_75t_R g952 ( 
.A(n_847),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_743),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_869),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_867),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_729),
.B(n_589),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_743),
.A2(n_721),
.B1(n_724),
.B2(n_592),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_759),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_847),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_814),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_817),
.B(n_725),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_822),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_870),
.B(n_698),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_826),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_794),
.B(n_689),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_739),
.B(n_595),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_879),
.Y(n_967)
);

AND3x1_ASAP7_75t_SL g968 ( 
.A(n_787),
.B(n_388),
.C(n_387),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_806),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_729),
.B(n_619),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_SL g971 ( 
.A1(n_885),
.A2(n_283),
.B1(n_266),
.B2(n_679),
.Y(n_971)
);

NOR2x1_ASAP7_75t_L g972 ( 
.A(n_786),
.B(n_695),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_867),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_745),
.B(n_605),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_876),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_867),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_884),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_888),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_892),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_764),
.B(n_697),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_773),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_773),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_759),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_869),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_867),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_SL g986 ( 
.A(n_804),
.B(n_723),
.C(n_219),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_781),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_792),
.B(n_606),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_792),
.B(n_724),
.Y(n_989)
);

CKINVDCx14_ASAP7_75t_R g990 ( 
.A(n_735),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_811),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_817),
.B(n_725),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_769),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_756),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_837),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_781),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_811),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_769),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_765),
.B(n_652),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_772),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_728),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_731),
.B(n_665),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_874),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_793),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_886),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_772),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_891),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_782),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_886),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_793),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_797),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_797),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_806),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_807),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_753),
.B(n_589),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_870),
.A2(n_673),
.B1(n_671),
.B2(n_665),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_SL g1017 ( 
.A(n_734),
.B(n_225),
.C(n_205),
.Y(n_1017)
);

BUFx4f_ASAP7_75t_L g1018 ( 
.A(n_753),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_807),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_815),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_809),
.A2(n_657),
.B1(n_652),
.B2(n_720),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_810),
.Y(n_1022)
);

BUFx8_ASAP7_75t_L g1023 ( 
.A(n_891),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_810),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_828),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_795),
.B(n_725),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_732),
.B(n_667),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_828),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_874),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_815),
.Y(n_1030)
);

NOR2x1p5_ASAP7_75t_L g1031 ( 
.A(n_868),
.B(n_843),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_832),
.Y(n_1032)
);

BUFx4f_ASAP7_75t_L g1033 ( 
.A(n_795),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_803),
.B(n_589),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_816),
.A2(n_673),
.B1(n_671),
.B2(n_718),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_887),
.A2(n_283),
.B1(n_693),
.B2(n_718),
.C(n_717),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_832),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_839),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_747),
.B(n_667),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_839),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_848),
.Y(n_1041)
);

AND3x1_ASAP7_75t_SL g1042 ( 
.A(n_865),
.B(n_11),
.C(n_12),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_868),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_848),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_858),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_816),
.A2(n_692),
.B1(n_693),
.B2(n_717),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_836),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_893),
.A2(n_657),
.B1(n_652),
.B2(n_716),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_874),
.B(n_715),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_858),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_815),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_748),
.A2(n_669),
.B(n_692),
.C(n_716),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_893),
.B(n_599),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_791),
.B(n_657),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_L g1055 ( 
.A(n_775),
.B(n_715),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_843),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_860),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_860),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_R g1059 ( 
.A(n_803),
.B(n_619),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_862),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_862),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_859),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_864),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_864),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_859),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_859),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_783),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_853),
.B(n_619),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_749),
.B(n_669),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_750),
.B(n_599),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_835),
.A2(n_599),
.B1(n_679),
.B2(n_716),
.C(n_659),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_783),
.B(n_648),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_827),
.B(n_771),
.C(n_873),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_730),
.B(n_679),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_R g1075 ( 
.A(n_844),
.B(n_856),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_878),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_770),
.B(n_648),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_758),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_789),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_813),
.A2(n_694),
.B1(n_666),
.B2(n_714),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_844),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_762),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_780),
.B(n_784),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_881),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_919),
.B(n_830),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_899),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_921),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_895),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_947),
.A2(n_854),
.B1(n_852),
.B2(n_849),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1074),
.A2(n_846),
.B(n_842),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_918),
.B(n_991),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_921),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_929),
.B(n_740),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_912),
.A2(n_755),
.B1(n_754),
.B2(n_801),
.Y(n_1094)
);

NAND2x1_ASAP7_75t_L g1095 ( 
.A(n_913),
.B(n_648),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_942),
.A2(n_872),
.B(n_866),
.Y(n_1096)
);

AND3x4_ASAP7_75t_L g1097 ( 
.A(n_902),
.B(n_861),
.C(n_856),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_915),
.A2(n_872),
.B(n_866),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_907),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_971),
.A2(n_805),
.B1(n_856),
.B2(n_844),
.Y(n_1100)
);

BUFx2_ASAP7_75t_SL g1101 ( 
.A(n_902),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1047),
.A2(n_924),
.B1(n_903),
.B2(n_910),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1031),
.B(n_824),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_924),
.A2(n_871),
.B1(n_850),
.B2(n_851),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_956),
.A2(n_845),
.B(n_841),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_961),
.B(n_740),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_901),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_956),
.A2(n_845),
.B(n_841),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_911),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1070),
.A2(n_834),
.B(n_821),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1039),
.A2(n_834),
.B(n_821),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1069),
.A2(n_742),
.B(n_831),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1015),
.A2(n_880),
.B(n_889),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_941),
.A2(n_863),
.B(n_890),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1015),
.A2(n_894),
.B(n_742),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_901),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_682),
.B(n_705),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1027),
.A2(n_682),
.B(n_705),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_997),
.B(n_877),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_1001),
.A2(n_999),
.B(n_1075),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_928),
.A2(n_840),
.B(n_825),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1052),
.A2(n_946),
.B(n_999),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_963),
.A2(n_687),
.B(n_688),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_994),
.A2(n_818),
.B1(n_782),
.B2(n_882),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_963),
.A2(n_687),
.B(n_688),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_966),
.A2(n_720),
.B(n_682),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_929),
.B(n_659),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_897),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_896),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_950),
.B(n_857),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1067),
.B(n_777),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_914),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1073),
.A2(n_808),
.B(n_820),
.C(n_855),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_980),
.B(n_670),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_925),
.B(n_685),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1084),
.B(n_685),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_974),
.A2(n_988),
.B(n_989),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1056),
.B(n_691),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1052),
.A2(n_705),
.B(n_720),
.Y(n_1139)
);

AND2x2_ASAP7_75t_SL g1140 ( 
.A(n_945),
.B(n_865),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_913),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1056),
.B(n_691),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1049),
.A2(n_688),
.B(n_694),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_905),
.A2(n_588),
.B1(n_722),
.B2(n_616),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_957),
.A2(n_1082),
.B(n_1078),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_SL g1146 ( 
.A1(n_920),
.A2(n_703),
.B(n_714),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1043),
.B(n_699),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_976),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_904),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1034),
.A2(n_855),
.B(n_722),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_908),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_SL g1152 ( 
.A1(n_1029),
.A2(n_699),
.B(n_700),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_969),
.B(n_700),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_969),
.B(n_701),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1007),
.B(n_701),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1034),
.A2(n_676),
.B(n_616),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1013),
.B(n_703),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1013),
.B(n_708),
.Y(n_1158)
);

BUFx4_ASAP7_75t_SL g1159 ( 
.A(n_967),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_1029),
.A2(n_708),
.B(n_710),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1043),
.B(n_1072),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1010),
.A2(n_710),
.B(n_722),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_914),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1072),
.B(n_588),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1010),
.A2(n_722),
.B(n_696),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1034),
.A2(n_722),
.B(n_696),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_976),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_923),
.B(n_588),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1073),
.A2(n_266),
.B(n_267),
.C(n_254),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1053),
.B(n_588),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1019),
.A2(n_696),
.B(n_676),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1071),
.A2(n_696),
.B(n_676),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_895),
.Y(n_1173)
);

O2A1O1Ixp5_ASAP7_75t_L g1174 ( 
.A1(n_1054),
.A2(n_1033),
.B(n_1018),
.C(n_1077),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_948),
.A2(n_596),
.B(n_240),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1019),
.A2(n_696),
.B(n_676),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1024),
.A2(n_676),
.B(n_644),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_931),
.B(n_616),
.Y(n_1178)
);

OA22x2_ASAP7_75t_L g1179 ( 
.A1(n_1008),
.A2(n_382),
.B1(n_251),
.B2(n_250),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1077),
.A2(n_596),
.B(n_246),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_916),
.B(n_522),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_1026),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_932),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_1017),
.A2(n_319),
.B(n_261),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_909),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_940),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1024),
.A2(n_644),
.B(n_616),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1025),
.A2(n_644),
.B(n_616),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_960),
.B(n_962),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1025),
.A2(n_644),
.B(n_596),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_922),
.A2(n_1033),
.B1(n_1018),
.B2(n_971),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1028),
.A2(n_596),
.B(n_563),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_SL g1193 ( 
.A1(n_1051),
.A2(n_12),
.B(n_17),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_SL g1194 ( 
.A1(n_1023),
.A2(n_332),
.B1(n_264),
.B2(n_385),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1003),
.B(n_541),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_964),
.B(n_19),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1028),
.A2(n_563),
.B(n_541),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_975),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_899),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_933),
.B(n_541),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1045),
.A2(n_563),
.B(n_541),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1051),
.A2(n_1062),
.B(n_1020),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1017),
.A2(n_381),
.B(n_271),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1020),
.A2(n_314),
.B(n_276),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_961),
.B(n_541),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1054),
.A2(n_1021),
.B(n_1048),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1045),
.A2(n_563),
.B(n_541),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_897),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_977),
.A2(n_338),
.B1(n_384),
.B2(n_378),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1020),
.A2(n_308),
.B(n_373),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1036),
.A2(n_267),
.B(n_563),
.C(n_360),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_952),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_992),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1035),
.A2(n_304),
.B(n_364),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_992),
.B(n_563),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_978),
.B(n_21),
.Y(n_1216)
);

BUFx8_ASAP7_75t_SL g1217 ( 
.A(n_917),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_979),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1035),
.A2(n_1046),
.B(n_1083),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_933),
.B(n_26),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1061),
.A2(n_267),
.B(n_121),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_981),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_953),
.B(n_26),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_982),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1023),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_984),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_987),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_935),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1061),
.A2(n_267),
.B(n_124),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1081),
.B(n_117),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_953),
.B(n_28),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_996),
.A2(n_267),
.B(n_351),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_986),
.A2(n_354),
.B(n_347),
.C(n_310),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1055),
.A2(n_111),
.B(n_189),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1003),
.B(n_298),
.Y(n_1235)
);

OA22x2_ASAP7_75t_L g1236 ( 
.A1(n_951),
.A2(n_954),
.B1(n_1076),
.B2(n_1044),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1046),
.A2(n_295),
.B(n_284),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_938),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1081),
.B(n_29),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1081),
.B(n_29),
.Y(n_1240)
);

NAND2x1_ASAP7_75t_L g1241 ( 
.A(n_906),
.B(n_108),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1081),
.B(n_30),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_943),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_955),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_938),
.A2(n_1009),
.B(n_939),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1088),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1230),
.B(n_973),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1161),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1092),
.Y(n_1249)
);

INVx4_ASAP7_75t_SL g1250 ( 
.A(n_1230),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1162),
.A2(n_1009),
.B(n_939),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1129),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1099),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1109),
.B(n_995),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1169),
.A2(n_1022),
.B(n_1014),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1245),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1087),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1245),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1107),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1100),
.A2(n_990),
.B1(n_936),
.B2(n_1079),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1169),
.B(n_986),
.C(n_898),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1149),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1182),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1102),
.B(n_1219),
.Y(n_1264)
);

CKINVDCx16_ASAP7_75t_R g1265 ( 
.A(n_1128),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1100),
.A2(n_1103),
.B1(n_990),
.B2(n_1155),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1151),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1089),
.A2(n_898),
.B(n_972),
.C(n_1006),
.Y(n_1268)
);

O2A1O1Ixp5_ASAP7_75t_L g1269 ( 
.A1(n_1122),
.A2(n_959),
.B(n_926),
.C(n_906),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1183),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1228),
.B(n_995),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1088),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1110),
.A2(n_965),
.B(n_927),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1107),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1130),
.A2(n_1000),
.B(n_1006),
.C(n_949),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1146),
.A2(n_1041),
.B(n_1037),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1137),
.A2(n_1172),
.B(n_1206),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1221),
.A2(n_1057),
.B(n_1011),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1213),
.B(n_959),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1221),
.A2(n_1229),
.B(n_1162),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1230),
.B(n_973),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1085),
.B(n_1155),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1087),
.A2(n_944),
.B1(n_1062),
.B2(n_1066),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1165),
.A2(n_1005),
.B(n_1004),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1185),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1159),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1091),
.B(n_943),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1116),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1147),
.B(n_1228),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1165),
.A2(n_1005),
.B(n_1012),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1150),
.A2(n_1032),
.B(n_1038),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1186),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1191),
.A2(n_1042),
.B(n_900),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1174),
.A2(n_927),
.B(n_1016),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1198),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1097),
.B(n_1076),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1097),
.B(n_1003),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1171),
.A2(n_1063),
.B(n_1050),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1243),
.B(n_936),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1119),
.B(n_936),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1094),
.A2(n_936),
.B1(n_927),
.B2(n_968),
.Y(n_1302)
);

CKINVDCx6p67_ASAP7_75t_R g1303 ( 
.A(n_1128),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1176),
.A2(n_1058),
.B(n_1064),
.Y(n_1304)
);

AOI221xp5_ASAP7_75t_L g1305 ( 
.A1(n_1124),
.A2(n_1121),
.B1(n_1120),
.B2(n_1131),
.C(n_1104),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1176),
.A2(n_1060),
.B(n_1080),
.Y(n_1306)
);

INVx8_ASAP7_75t_L g1307 ( 
.A(n_1205),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1177),
.A2(n_1080),
.B(n_1079),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1090),
.A2(n_1068),
.B(n_1040),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1229),
.A2(n_958),
.B(n_998),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1114),
.A2(n_1232),
.B(n_1170),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1170),
.A2(n_1068),
.B(n_983),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1177),
.A2(n_1016),
.B(n_993),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1112),
.A2(n_927),
.B(n_949),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1098),
.A2(n_944),
.B(n_927),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1220),
.A2(n_1042),
.B1(n_985),
.B2(n_900),
.Y(n_1316)
);

AOI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1214),
.A2(n_968),
.B1(n_970),
.B2(n_1059),
.C(n_1000),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1135),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1208),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1208),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1098),
.A2(n_256),
.B(n_279),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1182),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1187),
.A2(n_1030),
.B(n_926),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1218),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1182),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1217),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1211),
.A2(n_970),
.B(n_1059),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1187),
.A2(n_1188),
.B(n_1197),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1106),
.A2(n_1140),
.B1(n_936),
.B2(n_1212),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1217),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1211),
.A2(n_1066),
.B(n_1065),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1181),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1189),
.B(n_1003),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1132),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1133),
.A2(n_1030),
.B(n_955),
.C(n_1062),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1179),
.A2(n_1236),
.B1(n_1140),
.B2(n_1237),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1139),
.A2(n_985),
.B(n_1065),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1222),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1213),
.B(n_955),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1145),
.A2(n_1066),
.B(n_1065),
.Y(n_1340)
);

BUFx8_ASAP7_75t_L g1341 ( 
.A(n_1225),
.Y(n_1341)
);

AOI222xp33_ASAP7_75t_L g1342 ( 
.A1(n_1196),
.A2(n_955),
.B1(n_1065),
.B2(n_1062),
.C1(n_1020),
.C2(n_1066),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1132),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1153),
.B(n_937),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1086),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1163),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1188),
.A2(n_937),
.B(n_934),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1154),
.B(n_937),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1213),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1163),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1106),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1086),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1238),
.Y(n_1353)
);

OA21x2_ASAP7_75t_L g1354 ( 
.A1(n_1096),
.A2(n_937),
.B(n_934),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1087),
.B(n_934),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1111),
.A2(n_934),
.B(n_930),
.Y(n_1356)
);

CKINVDCx12_ASAP7_75t_R g1357 ( 
.A(n_1200),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1106),
.B(n_895),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1224),
.Y(n_1359)
);

BUFx2_ASAP7_75t_SL g1360 ( 
.A(n_1088),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1238),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1157),
.B(n_930),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1201),
.A2(n_930),
.B(n_895),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1158),
.B(n_930),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1096),
.A2(n_100),
.B(n_183),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1227),
.B(n_30),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1180),
.B(n_34),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1133),
.A2(n_38),
.B(n_39),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1199),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1088),
.B(n_112),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1199),
.B(n_44),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1173),
.B(n_110),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1101),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_SL g1374 ( 
.A1(n_1156),
.A2(n_46),
.B(n_47),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1207),
.A2(n_133),
.B(n_171),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1113),
.A2(n_126),
.B(n_167),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1115),
.A2(n_47),
.B(n_50),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1223),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1136),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1144),
.A2(n_52),
.A3(n_53),
.B(n_59),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1209),
.A2(n_52),
.B1(n_53),
.B2(n_63),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1134),
.B(n_63),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1190),
.A2(n_139),
.B(n_159),
.Y(n_1383)
);

CKINVDCx6p67_ASAP7_75t_R g1384 ( 
.A(n_1226),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1115),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1113),
.A2(n_1105),
.B(n_1108),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1190),
.A2(n_136),
.B(n_158),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1138),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1194),
.A2(n_1179),
.B1(n_1242),
.B2(n_1240),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1192),
.A2(n_135),
.B(n_155),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1231),
.A2(n_1126),
.B(n_1117),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1166),
.A2(n_106),
.B(n_154),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_L g1393 ( 
.A(n_1148),
.B(n_94),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1192),
.A2(n_1143),
.B(n_1108),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1141),
.A2(n_67),
.B1(n_70),
.B2(n_79),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1142),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1143),
.A2(n_84),
.B(n_146),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1216),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1105),
.A2(n_150),
.B(n_151),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1236),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1202),
.A2(n_67),
.B(n_186),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1205),
.B(n_1215),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1141),
.A2(n_1168),
.B1(n_1178),
.B2(n_1093),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1234),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1239),
.B(n_1184),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1093),
.A2(n_1226),
.B1(n_1164),
.B2(n_1167),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1118),
.A2(n_1123),
.B(n_1125),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1203),
.A2(n_1235),
.B1(n_1205),
.B2(n_1215),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1215),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1173),
.Y(n_1410)
);

AND2x2_ASAP7_75t_SL g1411 ( 
.A(n_1141),
.B(n_1173),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1173),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1127),
.B(n_1235),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1266),
.A2(n_1193),
.B1(n_1175),
.B2(n_1148),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1368),
.A2(n_1167),
.B1(n_1233),
.B2(n_1244),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1250),
.B(n_1402),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1305),
.A2(n_1204),
.B1(n_1210),
.B2(n_1244),
.Y(n_1417)
);

AOI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1293),
.A2(n_1233),
.B1(n_1152),
.B2(n_1160),
.C(n_1195),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1252),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1405),
.A2(n_1241),
.B(n_1195),
.C(n_1095),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1249),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1289),
.B(n_1127),
.Y(n_1422)
);

NAND2x1p5_ASAP7_75t_L g1423 ( 
.A(n_1257),
.B(n_1249),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1366),
.B(n_1282),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1366),
.B(n_1351),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1404),
.A2(n_1335),
.A3(n_1258),
.B(n_1256),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1264),
.A2(n_1260),
.B1(n_1336),
.B2(n_1400),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1264),
.A2(n_1302),
.B1(n_1261),
.B2(n_1381),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1247),
.B(n_1281),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1330),
.Y(n_1430)
);

O2A1O1Ixp5_ASAP7_75t_SL g1431 ( 
.A1(n_1378),
.A2(n_1367),
.B(n_1398),
.C(n_1385),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1262),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1330),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1338),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1257),
.B(n_1411),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1351),
.B(n_1265),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1268),
.A2(n_1389),
.B(n_1367),
.C(n_1335),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1373),
.A2(n_1369),
.B1(n_1371),
.B2(n_1377),
.C(n_1294),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1355),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1359),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1315),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1267),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1382),
.B(n_1248),
.Y(n_1443)
);

AND2x2_ASAP7_75t_SL g1444 ( 
.A(n_1411),
.B(n_1298),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1297),
.A2(n_1271),
.B1(n_1286),
.B2(n_1329),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1382),
.B(n_1402),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1270),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1277),
.A2(n_1391),
.B(n_1328),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1292),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1388),
.B(n_1396),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1314),
.A2(n_1273),
.B(n_1340),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_SL g1452 ( 
.A(n_1247),
.B(n_1281),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1318),
.A2(n_1379),
.B1(n_1332),
.B2(n_1301),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1402),
.B(n_1285),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1345),
.B(n_1352),
.Y(n_1455)
);

AO21x2_ASAP7_75t_L g1456 ( 
.A1(n_1404),
.A2(n_1309),
.B(n_1291),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1257),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1247),
.B(n_1281),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1295),
.B(n_1324),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1379),
.A2(n_1317),
.B1(n_1316),
.B2(n_1250),
.Y(n_1460)
);

INVx8_ASAP7_75t_L g1461 ( 
.A(n_1307),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1259),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1259),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1345),
.B(n_1352),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1341),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1274),
.Y(n_1466)
);

INVx6_ASAP7_75t_L g1467 ( 
.A(n_1257),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1247),
.A2(n_1281),
.B1(n_1287),
.B2(n_1395),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1253),
.A2(n_1254),
.B(n_1406),
.C(n_1319),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1303),
.Y(n_1470)
);

CKINVDCx16_ASAP7_75t_R g1471 ( 
.A(n_1326),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1250),
.B(n_1358),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1250),
.A2(n_1409),
.B1(n_1408),
.B2(n_1358),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1288),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1320),
.B(n_1303),
.Y(n_1475)
);

BUFx10_ASAP7_75t_L g1476 ( 
.A(n_1279),
.Y(n_1476)
);

NOR3xp33_ASAP7_75t_SL g1477 ( 
.A(n_1275),
.B(n_1300),
.C(n_1403),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1307),
.B(n_1413),
.Y(n_1478)
);

OAI22x1_ASAP7_75t_L g1479 ( 
.A1(n_1358),
.A2(n_1413),
.B1(n_1372),
.B2(n_1370),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1320),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1257),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1355),
.B(n_1279),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1344),
.B(n_1333),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1340),
.A2(n_1337),
.B(n_1407),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1283),
.A2(n_1349),
.B1(n_1279),
.B2(n_1307),
.Y(n_1485)
);

CKINVDCx6p67_ASAP7_75t_R g1486 ( 
.A(n_1384),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1349),
.B(n_1263),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1341),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1246),
.Y(n_1489)
);

NAND2xp33_ASAP7_75t_R g1490 ( 
.A(n_1315),
.B(n_1321),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1296),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1334),
.Y(n_1492)
);

AOI21xp33_ASAP7_75t_L g1493 ( 
.A1(n_1255),
.A2(n_1327),
.B(n_1315),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1307),
.B(n_1344),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1327),
.A2(n_1374),
.B1(n_1255),
.B2(n_1372),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1341),
.Y(n_1496)
);

CKINVDCx6p67_ASAP7_75t_R g1497 ( 
.A(n_1357),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1263),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1357),
.A2(n_1342),
.B1(n_1322),
.B2(n_1325),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1246),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1360),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1348),
.B(n_1362),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1322),
.B(n_1325),
.Y(n_1503)
);

INVx5_ASAP7_75t_L g1504 ( 
.A(n_1246),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_L g1505 ( 
.A(n_1246),
.B(n_1272),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1385),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1343),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1346),
.A2(n_1353),
.B1(n_1350),
.B2(n_1361),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1339),
.A2(n_1327),
.B1(n_1255),
.B2(n_1393),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1346),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1364),
.A2(n_1372),
.B1(n_1370),
.B2(n_1339),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_1360),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1246),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1350),
.B(n_1361),
.Y(n_1514)
);

AO31x2_ASAP7_75t_L g1515 ( 
.A1(n_1256),
.A2(n_1258),
.A3(n_1353),
.B(n_1410),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1370),
.A2(n_1376),
.B1(n_1412),
.B2(n_1272),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1337),
.B(n_1313),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1380),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1291),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1407),
.A2(n_1269),
.B(n_1376),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1272),
.B(n_1312),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1272),
.B(n_1312),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1380),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1339),
.B(n_1412),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1380),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1272),
.B(n_1312),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1380),
.B(n_1412),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1309),
.B(n_1356),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1356),
.B(n_1347),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1291),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1407),
.A2(n_1376),
.B(n_1363),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1299),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1321),
.A2(n_1365),
.B1(n_1380),
.B2(n_1374),
.Y(n_1533)
);

INVx8_ASAP7_75t_L g1534 ( 
.A(n_1401),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1354),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1321),
.A2(n_1365),
.B1(n_1386),
.B2(n_1392),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1386),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1304),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1394),
.A2(n_1306),
.B(n_1308),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_SL g1540 ( 
.A(n_1311),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1311),
.B(n_1309),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1331),
.B(n_1354),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1399),
.B(n_1323),
.Y(n_1543)
);

O2A1O1Ixp33_ASAP7_75t_SL g1544 ( 
.A1(n_1331),
.A2(n_1390),
.B(n_1387),
.C(n_1383),
.Y(n_1544)
);

INVx4_ASAP7_75t_SL g1545 ( 
.A(n_1383),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1276),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1276),
.A2(n_1365),
.B1(n_1313),
.B2(n_1399),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1304),
.B(n_1354),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1284),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1276),
.A2(n_1310),
.B1(n_1278),
.B2(n_1306),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1386),
.B(n_1284),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1290),
.B(n_1251),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1251),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1387),
.B(n_1397),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1390),
.A2(n_1397),
.B(n_1375),
.C(n_1278),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1278),
.B(n_1310),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1310),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1280),
.A2(n_1277),
.B(n_767),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1375),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1280),
.B(n_1282),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1280),
.A2(n_726),
.B1(n_1047),
.B2(n_649),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1293),
.A2(n_726),
.B1(n_1047),
.B2(n_649),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1250),
.B(n_1402),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1266),
.A2(n_1001),
.B1(n_649),
.B2(n_728),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1385),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1564),
.A2(n_1562),
.B1(n_1438),
.B2(n_1428),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1561),
.A2(n_1438),
.B1(n_1415),
.B2(n_1428),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1427),
.A2(n_1415),
.B1(n_1424),
.B2(n_1443),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1533),
.A2(n_1444),
.B1(n_1441),
.B2(n_1485),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_L g1571 ( 
.A1(n_1437),
.A2(n_1523),
.B(n_1518),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1425),
.B(n_1436),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1431),
.A2(n_1477),
.B(n_1420),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1558),
.A2(n_1516),
.B(n_1544),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1422),
.B(n_1455),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1445),
.A2(n_1460),
.B1(n_1485),
.B2(n_1468),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1414),
.A2(n_1468),
.B1(n_1469),
.B2(n_1421),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1419),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1515),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1483),
.B(n_1459),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1525),
.A2(n_1449),
.B1(n_1440),
.B2(n_1434),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1432),
.A2(n_1442),
.B1(n_1447),
.B2(n_1527),
.C(n_1493),
.Y(n_1582)
);

OAI211xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1418),
.A2(n_1477),
.B(n_1421),
.C(n_1450),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1493),
.A2(n_1450),
.B1(n_1414),
.B2(n_1453),
.C(n_1536),
.Y(n_1584)
);

AOI211xp5_ASAP7_75t_L g1585 ( 
.A1(n_1516),
.A2(n_1451),
.B(n_1536),
.C(n_1560),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1486),
.A2(n_1470),
.B1(n_1458),
.B2(n_1429),
.Y(n_1586)
);

AOI222xp33_ASAP7_75t_L g1587 ( 
.A1(n_1473),
.A2(n_1441),
.B1(n_1483),
.B2(n_1502),
.C1(n_1479),
.C2(n_1463),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1462),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1466),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1464),
.B(n_1475),
.Y(n_1590)
);

OAI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1495),
.A2(n_1418),
.B(n_1558),
.C(n_1470),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1497),
.A2(n_1458),
.B1(n_1429),
.B2(n_1495),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1474),
.Y(n_1593)
);

AO21x1_ASAP7_75t_L g1594 ( 
.A1(n_1490),
.A2(n_1511),
.B(n_1451),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1507),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1429),
.A2(n_1458),
.B1(n_1563),
.B2(n_1416),
.Y(n_1596)
);

OAI211xp5_ASAP7_75t_L g1597 ( 
.A1(n_1417),
.A2(n_1520),
.B(n_1509),
.C(n_1555),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1465),
.A2(n_1496),
.B1(n_1512),
.B2(n_1488),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1416),
.A2(n_1563),
.B1(n_1472),
.B2(n_1478),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1472),
.A2(n_1478),
.B1(n_1540),
.B2(n_1494),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1452),
.A2(n_1540),
.B1(n_1534),
.B2(n_1511),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1502),
.A2(n_1554),
.B1(n_1530),
.B2(n_1519),
.C(n_1541),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1499),
.A2(n_1471),
.B1(n_1435),
.B2(n_1423),
.Y(n_1603)
);

OAI21xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1498),
.A2(n_1501),
.B(n_1481),
.Y(n_1604)
);

AOI222xp33_ASAP7_75t_L g1605 ( 
.A1(n_1545),
.A2(n_1519),
.B1(n_1530),
.B2(n_1514),
.C1(n_1534),
.C2(n_1508),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1534),
.A2(n_1559),
.B1(n_1461),
.B2(n_1435),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1480),
.A2(n_1484),
.B1(n_1501),
.B2(n_1505),
.C(n_1551),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1423),
.A2(n_1482),
.B1(n_1487),
.B2(n_1503),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1461),
.A2(n_1546),
.B1(n_1457),
.B2(n_1467),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1461),
.A2(n_1491),
.B1(n_1492),
.B2(n_1510),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1439),
.A2(n_1467),
.B1(n_1457),
.B2(n_1481),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1500),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1546),
.A2(n_1457),
.B1(n_1522),
.B2(n_1521),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1430),
.A2(n_1524),
.B1(n_1526),
.B2(n_1433),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1506),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1433),
.Y(n_1616)
);

OAI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1547),
.A2(n_1504),
.B1(n_1517),
.B2(n_1565),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1524),
.A2(n_1545),
.B1(n_1528),
.B2(n_1456),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1528),
.A2(n_1537),
.B1(n_1557),
.B2(n_1565),
.C(n_1506),
.Y(n_1619)
);

OAI222xp33_ASAP7_75t_L g1620 ( 
.A1(n_1535),
.A2(n_1542),
.B1(n_1517),
.B2(n_1550),
.C1(n_1556),
.C2(n_1504),
.Y(n_1620)
);

A2O1A1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1484),
.A2(n_1542),
.B(n_1535),
.C(n_1556),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1448),
.A2(n_1543),
.B(n_1552),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1476),
.B(n_1489),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1537),
.A2(n_1549),
.B1(n_1548),
.B2(n_1529),
.C(n_1553),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1476),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1504),
.B(n_1513),
.Y(n_1626)
);

OR2x6_ASAP7_75t_SL g1627 ( 
.A(n_1538),
.B(n_1532),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1500),
.A2(n_1513),
.B1(n_1448),
.B2(n_1517),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1539),
.A2(n_1562),
.B1(n_726),
.B2(n_1438),
.C(n_1293),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1545),
.Y(n_1630)
);

AOI21xp33_ASAP7_75t_L g1631 ( 
.A1(n_1426),
.A2(n_1438),
.B(n_1405),
.Y(n_1631)
);

AOI222xp33_ASAP7_75t_L g1632 ( 
.A1(n_1426),
.A2(n_649),
.B1(n_536),
.B2(n_1564),
.C1(n_728),
.C2(n_1368),
.Y(n_1632)
);

AOI222xp33_ASAP7_75t_L g1633 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_536),
.B2(n_728),
.C1(n_1368),
.C2(n_1293),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1562),
.A2(n_1293),
.B(n_585),
.C(n_1561),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1637)
);

OR2x2_ASAP7_75t_SL g1638 ( 
.A(n_1471),
.B(n_1265),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1561),
.B2(n_1438),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1264),
.B2(n_1302),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1642)
);

AOI222xp33_ASAP7_75t_L g1643 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_536),
.B2(n_728),
.C1(n_1368),
.C2(n_1293),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_L g1644 ( 
.A1(n_1562),
.A2(n_1293),
.B(n_585),
.C(n_1561),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1430),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1419),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1047),
.B2(n_649),
.Y(n_1647)
);

OA21x2_ASAP7_75t_L g1648 ( 
.A1(n_1520),
.A2(n_1531),
.B(n_1493),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1561),
.B2(n_1438),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1264),
.B2(n_1302),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1489),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1424),
.B(n_1443),
.Y(n_1655)
);

NAND2x1_ASAP7_75t_L g1656 ( 
.A(n_1429),
.B(n_1458),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1419),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1562),
.A2(n_947),
.B(n_1368),
.C(n_1437),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1438),
.A2(n_649),
.B1(n_1368),
.B2(n_1428),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1454),
.B(n_1446),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1562),
.A2(n_1293),
.B(n_1561),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1264),
.B2(n_1302),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1419),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1562),
.B(n_1305),
.C(n_1437),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1438),
.A2(n_887),
.B1(n_503),
.B2(n_838),
.C(n_585),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1419),
.Y(n_1668)
);

BUFx4f_ASAP7_75t_SL g1669 ( 
.A(n_1486),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1419),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1471),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1561),
.B(n_1264),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1424),
.B(n_1443),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1558),
.A2(n_1277),
.B(n_1368),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1562),
.A2(n_947),
.B(n_1368),
.C(n_1437),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1561),
.B2(n_1438),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1562),
.A2(n_1293),
.B(n_1561),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1562),
.A2(n_1293),
.B1(n_1561),
.B2(n_1438),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1562),
.B(n_1293),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1430),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1564),
.A2(n_649),
.B1(n_1266),
.B2(n_1100),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1588),
.Y(n_1685)
);

INVxp67_ASAP7_75t_R g1686 ( 
.A(n_1586),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1589),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1568),
.B(n_1636),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1593),
.Y(n_1689)
);

INVx5_ASAP7_75t_L g1690 ( 
.A(n_1630),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1655),
.B(n_1580),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1579),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1615),
.B(n_1674),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1579),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1639),
.B(n_1651),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1595),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1633),
.A2(n_1643),
.B1(n_1661),
.B2(n_1632),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1578),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1627),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1646),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1673),
.B(n_1658),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1648),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1594),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1602),
.B(n_1619),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1654),
.B(n_1662),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1585),
.B(n_1665),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1668),
.B(n_1671),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1656),
.B(n_1675),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1590),
.B(n_1621),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1621),
.B(n_1624),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1604),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1571),
.B(n_1567),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1628),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1631),
.B(n_1582),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1566),
.A2(n_1683),
.B1(n_1637),
.B2(n_1642),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1570),
.B(n_1622),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1618),
.B(n_1648),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1618),
.B(n_1648),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1581),
.B(n_1577),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1607),
.B(n_1584),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1597),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1574),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1614),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1566),
.A2(n_1647),
.B1(n_1681),
.B2(n_1660),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1612),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1613),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1681),
.B(n_1576),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1653),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1640),
.B(n_1680),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1666),
.B(n_1629),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1650),
.B(n_1678),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1617),
.B(n_1638),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1605),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1600),
.B(n_1591),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1573),
.A2(n_1620),
.B(n_1679),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1612),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1592),
.B(n_1663),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1641),
.B(n_1664),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1653),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1711),
.B(n_1653),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1725),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_R g1742 ( 
.A(n_1728),
.B(n_1672),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1692),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1711),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1690),
.B(n_1653),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1569),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1700),
.Y(n_1747)
);

AOI222xp33_ASAP7_75t_L g1748 ( 
.A1(n_1730),
.A2(n_1667),
.B1(n_1569),
.B2(n_1635),
.C1(n_1644),
.C2(n_1676),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1697),
.A2(n_1683),
.B1(n_1634),
.B2(n_1637),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1730),
.A2(n_1660),
.B1(n_1676),
.B2(n_1583),
.C(n_1649),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1685),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1691),
.B(n_1608),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1685),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1693),
.B(n_1701),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1739),
.B(n_1616),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1687),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1724),
.A2(n_1603),
.B1(n_1652),
.B2(n_1641),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1709),
.B(n_1601),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1739),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1694),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1687),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1689),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1697),
.A2(n_1738),
.B1(n_1729),
.B2(n_1724),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1709),
.B(n_1623),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1715),
.A2(n_1642),
.B1(n_1677),
.B2(n_1670),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1706),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1725),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1706),
.Y(n_1769)
);

NAND3xp33_ASAP7_75t_L g1770 ( 
.A(n_1721),
.B(n_1664),
.C(n_1652),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1690),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1696),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1721),
.B(n_1587),
.C(n_1606),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1684),
.B(n_1596),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_R g1775 ( 
.A(n_1728),
.B(n_1645),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1715),
.A2(n_1733),
.B1(n_1712),
.B2(n_1677),
.Y(n_1776)
);

OAI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1729),
.A2(n_1634),
.B(n_1670),
.C(n_1659),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1684),
.B(n_1599),
.Y(n_1778)
);

AO21x2_ASAP7_75t_L g1779 ( 
.A1(n_1714),
.A2(n_1611),
.B(n_1626),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1688),
.B(n_1599),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1735),
.A2(n_1649),
.B1(n_1659),
.B2(n_1657),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1708),
.B(n_1625),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1696),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1738),
.A2(n_1657),
.B1(n_1609),
.B2(n_1598),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1736),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1731),
.A2(n_1669),
.B1(n_1610),
.B2(n_1682),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1720),
.B(n_1669),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1722),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1693),
.B(n_1701),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1712),
.A2(n_1704),
.B1(n_1703),
.B2(n_1714),
.C(n_1737),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1744),
.B(n_1716),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1788),
.B(n_1703),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1778),
.B(n_1702),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_SL g1794 ( 
.A(n_1745),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1747),
.B(n_1750),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1778),
.B(n_1716),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1780),
.B(n_1717),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1747),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1780),
.B(n_1702),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1750),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1770),
.A2(n_1704),
.B(n_1710),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1779),
.B(n_1710),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1774),
.B(n_1717),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1779),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1743),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1774),
.B(n_1718),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1755),
.B(n_1699),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1767),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1752),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1752),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1755),
.B(n_1699),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1779),
.B(n_1754),
.Y(n_1812)
);

BUFx12f_ASAP7_75t_L g1813 ( 
.A(n_1740),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1765),
.B(n_1718),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1765),
.B(n_1713),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1754),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1789),
.B(n_1713),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1757),
.B(n_1720),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1769),
.B(n_1705),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1762),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1782),
.B(n_1705),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1782),
.B(n_1688),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1782),
.B(n_1695),
.Y(n_1823)
);

NOR2xp67_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1732),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1763),
.B(n_1707),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1782),
.B(n_1695),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1742),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1771),
.B(n_1708),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1782),
.B(n_1702),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1772),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1789),
.B(n_1732),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1761),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1792),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1830),
.Y(n_1834)
);

NOR2x1_ASAP7_75t_L g1835 ( 
.A(n_1827),
.B(n_1740),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1830),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1809),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1818),
.B(n_1772),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1809),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1791),
.B(n_1740),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1791),
.B(n_1745),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1791),
.B(n_1745),
.Y(n_1843)
);

AOI21xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1827),
.A2(n_1787),
.B(n_1764),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1818),
.B(n_1746),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1794),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1809),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1796),
.B(n_1783),
.Y(n_1848)
);

NOR3x1_ASAP7_75t_L g1849 ( 
.A(n_1827),
.B(n_1770),
.C(n_1790),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1805),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1810),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_1783),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1817),
.B(n_1746),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1817),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1815),
.B(n_1745),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1817),
.B(n_1753),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1810),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1832),
.Y(n_1858)
);

NAND2x1p5_ASAP7_75t_L g1859 ( 
.A(n_1824),
.B(n_1690),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1815),
.B(n_1741),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1810),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1796),
.B(n_1707),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1815),
.B(n_1768),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1821),
.B(n_1785),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1816),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1821),
.B(n_1760),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1802),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1805),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1816),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1831),
.B(n_1753),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1816),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1832),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1820),
.Y(n_1873)
);

OAI21xp33_ASAP7_75t_L g1874 ( 
.A1(n_1801),
.A2(n_1748),
.B(n_1731),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1798),
.B(n_1698),
.Y(n_1875)
);

NOR2x1_ASAP7_75t_SL g1876 ( 
.A(n_1856),
.B(n_1813),
.Y(n_1876)
);

AOI31xp67_ASAP7_75t_SL g1877 ( 
.A1(n_1844),
.A2(n_1802),
.A3(n_1792),
.B(n_1801),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1837),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1853),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1842),
.Y(n_1880)
);

OR2x4_ASAP7_75t_L g1881 ( 
.A(n_1853),
.B(n_1807),
.Y(n_1881)
);

NOR3xp33_ASAP7_75t_SL g1882 ( 
.A(n_1874),
.B(n_1760),
.C(n_1786),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1837),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1845),
.B(n_1831),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1842),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1874),
.B(n_1808),
.Y(n_1886)
);

NAND4xp25_ASAP7_75t_L g1887 ( 
.A(n_1849),
.B(n_1751),
.C(n_1758),
.D(n_1773),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1845),
.B(n_1831),
.Y(n_1888)
);

NOR2x1_ASAP7_75t_L g1889 ( 
.A(n_1835),
.B(n_1807),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1835),
.B(n_1846),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1840),
.B(n_1821),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1839),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1846),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1839),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1870),
.A2(n_1781),
.B1(n_1749),
.B2(n_1733),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1862),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1862),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1840),
.B(n_1841),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1844),
.B(n_1807),
.Y(n_1899)
);

OAI33xp33_ASAP7_75t_L g1900 ( 
.A1(n_1867),
.A2(n_1812),
.A3(n_1804),
.B1(n_1811),
.B2(n_1795),
.B3(n_1800),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1833),
.B(n_1808),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1846),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1856),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1841),
.B(n_1822),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1846),
.B(n_1824),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1866),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1847),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1843),
.B(n_1824),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1833),
.B(n_1819),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1847),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1854),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1870),
.B(n_1819),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1843),
.B(n_1822),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1855),
.B(n_1822),
.Y(n_1914)
);

NOR4xp25_ASAP7_75t_L g1915 ( 
.A(n_1849),
.B(n_1804),
.C(n_1727),
.D(n_1812),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1842),
.Y(n_1916)
);

AOI211xp5_ASAP7_75t_SL g1917 ( 
.A1(n_1834),
.A2(n_1811),
.B(n_1829),
.C(n_1784),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1851),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1866),
.B(n_1811),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1851),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1903),
.B(n_1848),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1879),
.B(n_1848),
.Y(n_1922)
);

O2A1O1Ixp33_ASAP7_75t_SL g1923 ( 
.A1(n_1917),
.A2(n_1852),
.B(n_1838),
.C(n_1723),
.Y(n_1923)
);

NAND2x1p5_ASAP7_75t_L g1924 ( 
.A(n_1889),
.B(n_1728),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1911),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1878),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1915),
.B(n_1836),
.C(n_1834),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1887),
.A2(n_1735),
.B1(n_1766),
.B2(n_1719),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1878),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1899),
.B(n_1852),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1886),
.A2(n_1877),
.B1(n_1727),
.B2(n_1876),
.Y(n_1931)
);

OAI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1881),
.A2(n_1737),
.B1(n_1719),
.B2(n_1735),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1883),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1883),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1906),
.B(n_1838),
.Y(n_1935)
);

NAND2xp33_ASAP7_75t_L g1936 ( 
.A(n_1882),
.B(n_1775),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1892),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1884),
.B(n_1836),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1892),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1894),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1894),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1906),
.B(n_1813),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1907),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1900),
.A2(n_1881),
.B(n_1877),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1919),
.B(n_1813),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1896),
.B(n_1797),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1895),
.A2(n_1735),
.B1(n_1777),
.B2(n_1776),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1907),
.Y(n_1948)
);

O2A1O1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1901),
.A2(n_1735),
.B(n_1734),
.C(n_1797),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1884),
.B(n_1825),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1910),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1910),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1897),
.B(n_1797),
.Y(n_1953)
);

AOI321xp33_ASAP7_75t_L g1954 ( 
.A1(n_1881),
.A2(n_1734),
.A3(n_1759),
.B1(n_1806),
.B2(n_1803),
.C(n_1726),
.Y(n_1954)
);

AOI21xp33_ASAP7_75t_L g1955 ( 
.A1(n_1893),
.A2(n_1850),
.B(n_1872),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1893),
.B(n_1865),
.C(n_1857),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1918),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1926),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1929),
.Y(n_1959)
);

OAI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1944),
.A2(n_1888),
.B1(n_1723),
.B2(n_1686),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1933),
.Y(n_1961)
);

INVxp67_ASAP7_75t_L g1962 ( 
.A(n_1942),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1931),
.B(n_1876),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1931),
.B(n_1890),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1944),
.B(n_1954),
.Y(n_1965)
);

NAND2xp33_ASAP7_75t_SL g1966 ( 
.A(n_1925),
.B(n_1902),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1923),
.A2(n_1905),
.B(n_1890),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1945),
.B(n_1902),
.Y(n_1968)
);

OAI21xp33_ASAP7_75t_L g1969 ( 
.A1(n_1930),
.A2(n_1909),
.B(n_1890),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1949),
.A2(n_1885),
.B1(n_1916),
.B2(n_1880),
.C(n_1918),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1950),
.B(n_1898),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1938),
.Y(n_1972)
);

OAI211xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1949),
.A2(n_1912),
.B(n_1920),
.C(n_1888),
.Y(n_1973)
);

AOI211xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1932),
.A2(n_1955),
.B(n_1936),
.C(n_1935),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1934),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1922),
.Y(n_1976)
);

OAI32xp33_ASAP7_75t_L g1977 ( 
.A1(n_1927),
.A2(n_1859),
.A3(n_1920),
.B1(n_1916),
.B2(n_1880),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1937),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1939),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1940),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_L g1981 ( 
.A(n_1956),
.B(n_1908),
.Y(n_1981)
);

INVxp67_ASAP7_75t_SL g1982 ( 
.A(n_1924),
.Y(n_1982)
);

OAI321xp33_ASAP7_75t_L g1983 ( 
.A1(n_1947),
.A2(n_1726),
.A3(n_1859),
.B1(n_1723),
.B2(n_1885),
.C(n_1759),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1928),
.B(n_1898),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1971),
.B(n_1963),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1965),
.A2(n_1924),
.B(n_1957),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1972),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1958),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1964),
.A2(n_1921),
.B(n_1952),
.Y(n_1989)
);

NOR2x1_ASAP7_75t_L g1990 ( 
.A(n_1973),
.B(n_1941),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1968),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1958),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1972),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1976),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1976),
.B(n_1953),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1966),
.Y(n_1996)
);

NAND2xp33_ASAP7_75t_R g1997 ( 
.A(n_1963),
.B(n_1908),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1961),
.Y(n_1998)
);

XNOR2x1_ASAP7_75t_L g1999 ( 
.A(n_1960),
.B(n_1803),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1971),
.B(n_1914),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1961),
.Y(n_2001)
);

XOR2xp5_ASAP7_75t_L g2002 ( 
.A(n_1984),
.B(n_1946),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1981),
.B(n_1914),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1975),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1991),
.B(n_1962),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1987),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_2004),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_2004),
.Y(n_2008)
);

AOI211x1_ASAP7_75t_L g2009 ( 
.A1(n_1989),
.A2(n_1977),
.B(n_1967),
.C(n_1969),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2004),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1994),
.Y(n_2011)
);

AOI211xp5_ASAP7_75t_SL g2012 ( 
.A1(n_1986),
.A2(n_1983),
.B(n_1970),
.C(n_1982),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1985),
.B(n_1904),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1985),
.B(n_1966),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1996),
.A2(n_1977),
.B(n_1974),
.Y(n_2015)
);

AOI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1996),
.A2(n_1975),
.B(n_1979),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_2015),
.A2(n_2002),
.B1(n_1990),
.B2(n_1997),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_2012),
.A2(n_1990),
.B(n_1986),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_2009),
.B(n_1995),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2007),
.Y(n_2020)
);

O2A1O1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_2016),
.A2(n_1993),
.B(n_1994),
.C(n_2001),
.Y(n_2021)
);

AOI221x1_ASAP7_75t_L g2022 ( 
.A1(n_2016),
.A2(n_2011),
.B1(n_2006),
.B2(n_2005),
.C(n_2010),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2013),
.B(n_2000),
.Y(n_2023)
);

AOI222xp33_ASAP7_75t_L g2024 ( 
.A1(n_2008),
.A2(n_1993),
.B1(n_1988),
.B2(n_2001),
.C1(n_1992),
.C2(n_1998),
.Y(n_2024)
);

AOI211x1_ASAP7_75t_L g2025 ( 
.A1(n_2014),
.A2(n_2003),
.B(n_2000),
.C(n_1959),
.Y(n_2025)
);

OAI211xp5_ASAP7_75t_SL g2026 ( 
.A1(n_2015),
.A2(n_1988),
.B(n_1992),
.C(n_1998),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_2009),
.B(n_2003),
.C(n_1995),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_SL g2028 ( 
.A1(n_2018),
.A2(n_1999),
.B1(n_2002),
.B2(n_1980),
.Y(n_2028)
);

NAND2xp33_ASAP7_75t_SL g2029 ( 
.A(n_2023),
.B(n_1978),
.Y(n_2029)
);

NOR2xp67_ASAP7_75t_L g2030 ( 
.A(n_2027),
.B(n_1943),
.Y(n_2030)
);

OAI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_2017),
.A2(n_1999),
.B1(n_1948),
.B2(n_1951),
.C(n_1859),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_SL g2032 ( 
.A1(n_2026),
.A2(n_1908),
.B(n_1756),
.C(n_1913),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2025),
.B(n_1904),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_2019),
.B(n_2021),
.Y(n_2034)
);

OAI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_2020),
.A2(n_1913),
.B1(n_1871),
.B2(n_1869),
.Y(n_2035)
);

NOR4xp25_ASAP7_75t_L g2036 ( 
.A(n_2034),
.B(n_2022),
.C(n_2024),
.D(n_1891),
.Y(n_2036)
);

NOR2xp67_ASAP7_75t_L g2037 ( 
.A(n_2031),
.B(n_1891),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_2030),
.A2(n_2029),
.B(n_2028),
.Y(n_2038)
);

NAND3x1_ASAP7_75t_L g2039 ( 
.A(n_2033),
.B(n_1855),
.C(n_1860),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_2035),
.Y(n_2040)
);

NAND4xp75_ASAP7_75t_L g2041 ( 
.A(n_2032),
.B(n_1803),
.C(n_1806),
.D(n_1829),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2029),
.Y(n_2042)
);

AND4x1_ASAP7_75t_L g2043 ( 
.A(n_2036),
.B(n_1860),
.C(n_1863),
.D(n_1864),
.Y(n_2043)
);

NAND3x1_ASAP7_75t_L g2044 ( 
.A(n_2038),
.B(n_1863),
.C(n_1864),
.Y(n_2044)
);

NOR4xp25_ASAP7_75t_L g2045 ( 
.A(n_2042),
.B(n_1873),
.C(n_1861),
.D(n_1865),
.Y(n_2045)
);

NOR3xp33_ASAP7_75t_SL g2046 ( 
.A(n_2041),
.B(n_2040),
.C(n_2039),
.Y(n_2046)
);

AND4x1_ASAP7_75t_L g2047 ( 
.A(n_2037),
.B(n_1829),
.C(n_1823),
.D(n_1826),
.Y(n_2047)
);

OAI211xp5_ASAP7_75t_SL g2048 ( 
.A1(n_2038),
.A2(n_1871),
.B(n_1873),
.C(n_1857),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_2044),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2046),
.B(n_2043),
.Y(n_2050)
);

CKINVDCx20_ASAP7_75t_R g2051 ( 
.A(n_2048),
.Y(n_2051)
);

NAND4xp25_ASAP7_75t_L g2052 ( 
.A(n_2047),
.B(n_1739),
.C(n_1828),
.D(n_1829),
.Y(n_2052)
);

AOI22x1_ASAP7_75t_L g2053 ( 
.A1(n_2049),
.A2(n_2045),
.B1(n_1869),
.B2(n_1861),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2053),
.B(n_2050),
.Y(n_2054)
);

NOR2xp67_ASAP7_75t_L g2055 ( 
.A(n_2054),
.B(n_2052),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_2054),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2056),
.A2(n_2051),
.B1(n_1858),
.B2(n_1872),
.Y(n_2057)
);

XNOR2xp5_ASAP7_75t_L g2058 ( 
.A(n_2055),
.B(n_1806),
.Y(n_2058)
);

BUFx2_ASAP7_75t_L g2059 ( 
.A(n_2058),
.Y(n_2059)
);

AOI21xp33_ASAP7_75t_SL g2060 ( 
.A1(n_2057),
.A2(n_1872),
.B(n_1868),
.Y(n_2060)
);

AOI322xp5_ASAP7_75t_L g2061 ( 
.A1(n_2059),
.A2(n_1868),
.A3(n_1850),
.B1(n_1858),
.B2(n_1814),
.C1(n_1799),
.C2(n_1793),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_2061),
.A2(n_2060),
.B1(n_1850),
.B2(n_1858),
.Y(n_2062)
);

AOI211xp5_ASAP7_75t_L g2063 ( 
.A1(n_2062),
.A2(n_1728),
.B(n_1875),
.C(n_1793),
.Y(n_2063)
);


endmodule