module real_jpeg_14946_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_33),
.B1(n_49),
.B2(n_51),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_4),
.B(n_26),
.C(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_4),
.B(n_44),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_24),
.C(n_30),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_4),
.B(n_51),
.C(n_59),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_52),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_49),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_56),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_253)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_250),
.Y(n_11)
);

OAI21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_237),
.B(n_249),
.Y(n_12)
);

AOI21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_205),
.B(n_234),
.Y(n_13)
);

AO21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_103),
.B(n_204),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_85),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_16),
.B(n_85),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_66),
.C(n_77),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_17),
.B(n_66),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_46),
.B2(n_65),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_18),
.A2(n_19),
.B1(n_79),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_18),
.A2(n_19),
.B1(n_117),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_34),
.B2(n_45),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_20),
.A2(n_21),
.B1(n_57),
.B2(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_121),
.C(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_20),
.A2(n_21),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_34),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_21),
.A2(n_97),
.B(n_101),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_21),
.B(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_21),
.B(n_113),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_21),
.A2(n_113),
.B(n_150),
.C(n_155),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_32),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_22),
.A2(n_29),
.B1(n_32),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_22),
.A2(n_29),
.B1(n_217),
.B2(n_230),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_22),
.A2(n_29),
.B(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_29),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_23)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

OA22x2_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_43),
.Y(n_44)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_26),
.B(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_30),
.A2(n_31),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_30),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_33),
.B(n_75),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_33),
.B(n_54),
.Y(n_181)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_34),
.A2(n_45),
.B1(n_67),
.B2(n_68),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_34),
.A2(n_45),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_34),
.A2(n_45),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_34),
.A2(n_45),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_34),
.A2(n_45),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_34),
.B(n_214),
.C(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_34),
.B(n_226),
.C(n_232),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_35),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_37),
.B(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_40),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

AOI211xp5_ASAP7_75t_SL g137 ( 
.A1(n_45),
.A2(n_57),
.B(n_84),
.C(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_45),
.A2(n_67),
.B(n_91),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_45),
.B(n_213),
.C(n_229),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_78),
.B(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_47),
.A2(n_57),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_53),
.B1(n_54),
.B2(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_49),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_57),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_57),
.A2(n_80),
.B1(n_113),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_113),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_57),
.A2(n_113),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_57),
.A2(n_113),
.B1(n_167),
.B2(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_57),
.B(n_121),
.C(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_57),
.B(n_157),
.C(n_161),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_64),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_62),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_58),
.B(n_62),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_76),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_71),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_83),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_83),
.B(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_102),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_90),
.B(n_95),
.C(n_102),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_100),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_101),
.A2(n_209),
.B1(n_210),
.B2(n_219),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_101),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_123),
.B(n_203),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_107),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.C(n_115),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_201)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_115),
.A2(n_116),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_122),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_122),
.B1(n_132),
.B2(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_152),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_121),
.A2(n_122),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_121),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_121),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_122),
.B(n_183),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_144),
.B(n_197),
.C(n_202),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_131),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_126),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_127),
.A2(n_128),
.B1(n_150),
.B2(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_136),
.B(n_140),
.C(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_191),
.B(n_196),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_163),
.B(n_190),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_186),
.B(n_189),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_175),
.B(n_185),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_195),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_222),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_221),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_221),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_220),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_219),
.C(n_220),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_214),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_233),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_232),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_248),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_238),
.B(n_248),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_243),
.C(n_244),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_252),
.B(n_254),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule