module fake_jpeg_18942_n_325 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_0),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_45),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_21),
.B(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_34),
.B1(n_44),
.B2(n_24),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_61),
.B(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_56),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_33),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_35),
.C(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_24),
.B1(n_41),
.B2(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_60),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_39),
.B(n_41),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_41),
.B1(n_45),
.B2(n_34),
.Y(n_76)
);

BUFx24_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_36),
.C(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_36),
.C(n_29),
.Y(n_80)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_46),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_67),
.B1(n_49),
.B2(n_29),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_34),
.B1(n_24),
.B2(n_50),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_73),
.B(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_59),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_104),
.B(n_11),
.Y(n_143)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_105),
.B(n_110),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_62),
.C(n_63),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_82),
.C(n_52),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_119),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_43),
.C(n_59),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_115),
.B(n_13),
.C(n_15),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_72),
.B1(n_51),
.B2(n_76),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_127),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_72),
.B1(n_62),
.B2(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_79),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_70),
.B1(n_73),
.B2(n_71),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_67),
.B1(n_50),
.B2(n_24),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_129),
.B1(n_97),
.B2(n_83),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_90),
.B(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_95),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_31),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_30),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_30),
.B1(n_31),
.B2(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_92),
.B1(n_94),
.B2(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_81),
.Y(n_133)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_138),
.B1(n_152),
.B2(n_104),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_108),
.B1(n_104),
.B2(n_110),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_150),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_86),
.B1(n_29),
.B2(n_93),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_141),
.A2(n_163),
.B1(n_11),
.B2(n_23),
.Y(n_195)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_161),
.B(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_151),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_82),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_121),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_54),
.B1(n_30),
.B2(n_28),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_155),
.B1(n_164),
.B2(n_12),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_136),
.C(n_118),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_82),
.B(n_20),
.C(n_12),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_28),
.B1(n_12),
.B2(n_19),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_21),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_157),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_156),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_28),
.B1(n_56),
.B2(n_19),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_52),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_52),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_108),
.A2(n_28),
.B1(n_20),
.B2(n_21),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_52),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_165),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_103),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_155),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_179),
.C(n_162),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_103),
.B(n_104),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_184),
.B(n_186),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_102),
.C(n_128),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_187),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_101),
.B1(n_20),
.B2(n_12),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_191),
.B1(n_152),
.B2(n_23),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_101),
.B(n_20),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_140),
.A2(n_19),
.B(n_23),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_13),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_13),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_134),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_134),
.A2(n_19),
.B1(n_56),
.B2(n_22),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_164),
.B1(n_142),
.B2(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_156),
.B1(n_11),
.B2(n_22),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_200),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_208),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_131),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_217),
.B(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_170),
.B(n_131),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_158),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_159),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_130),
.C(n_148),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_168),
.B1(n_177),
.B2(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

AO22x1_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_143),
.B1(n_160),
.B2(n_151),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_195),
.B1(n_166),
.B2(n_174),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_166),
.B1(n_178),
.B2(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_237),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_185),
.B(n_173),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_179),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_180),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_189),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_206),
.C(n_218),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_185),
.B1(n_188),
.B2(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_241),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_186),
.B(n_188),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_204),
.B(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_205),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_206),
.B1(n_218),
.B2(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_239),
.B(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_13),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_233),
.B(n_219),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_261),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_259),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_25),
.C(n_17),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.C(n_226),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_231),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_253),
.A3(n_252),
.B1(n_247),
.B2(n_254),
.C1(n_240),
.C2(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_272),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_221),
.B(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_224),
.C(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_25),
.C(n_17),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_276),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_25),
.C(n_17),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_17),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_279),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_250),
.B(n_259),
.Y(n_279)
);

OAI221xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_255),
.B1(n_249),
.B2(n_18),
.C(n_13),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_281),
.B(n_286),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_15),
.B(n_10),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_275),
.A2(n_25),
.B1(n_8),
.B2(n_9),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_266),
.Y(n_294)
);

AO221x1_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_15),
.B1(n_17),
.B2(n_14),
.C(n_25),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_1),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_267),
.A2(n_6),
.B(n_10),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_277),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_264),
.C(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_272),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_17),
.C(n_14),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_9),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.C(n_2),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_1),
.C(n_2),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_304),
.A2(n_303),
.B1(n_6),
.B2(n_8),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_283),
.B1(n_288),
.B2(n_6),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_311),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_312),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_6),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_306),
.B(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_307),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_304),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_316),
.C(n_315),
.Y(n_320)
);

A2O1A1O1Ixp25_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_8),
.B(n_4),
.C(n_5),
.D(n_3),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_8),
.C(n_4),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_3),
.C(n_4),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_5),
.B(n_3),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_4),
.B(n_5),
.Y(n_325)
);


endmodule