module fake_aes_7905_n_688 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_688);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_688;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_84;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_72), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_73), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_40), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_53), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_70), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_35), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_76), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_59), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_46), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_32), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_11), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_34), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_61), .Y(n_91) );
CKINVDCx14_ASAP7_75t_R g92 ( .A(n_54), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_71), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_13), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_39), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_29), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_31), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_22), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_16), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_63), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_20), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_14), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_8), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_56), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_22), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_69), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_48), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_60), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_26), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_12), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_18), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_20), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_49), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_44), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_24), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_25), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_43), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_97), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_122), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_102), .B(n_0), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_111), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_114), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_80), .B(n_1), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_115), .B(n_1), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_78), .B(n_2), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_80), .B(n_2), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_111), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_89), .B(n_3), .Y(n_145) );
NOR2xp33_ASAP7_75t_SL g146 ( .A(n_79), .B(n_75), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_89), .B(n_3), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_92), .B(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_77), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_77), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_94), .B(n_4), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_94), .B(n_5), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_100), .B(n_5), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_91), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_91), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_96), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_100), .B(n_6), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_96), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_101), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
XOR2x2_ASAP7_75t_L g168 ( .A(n_129), .B(n_99), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_130), .B(n_81), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
OAI22xp33_ASAP7_75t_SL g171 ( .A1(n_140), .A2(n_118), .B1(n_95), .B2(n_108), .Y(n_171) );
AO22x2_ASAP7_75t_L g172 ( .A1(n_156), .A2(n_118), .B1(n_95), .B2(n_124), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_130), .B(n_93), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_131), .B(n_106), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_131), .B(n_106), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_149), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_129), .B(n_117), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_149), .B(n_117), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_128), .B(n_81), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_150), .B(n_103), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_150), .B(n_105), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_156), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_131), .B(n_104), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_151), .B(n_105), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_131), .B(n_108), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_151), .B(n_109), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_127), .Y(n_201) );
INVxp67_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_153), .B(n_109), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_131), .B(n_113), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_138), .B(n_113), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_127), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_153), .B(n_104), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_154), .B(n_116), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_127), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_138), .B(n_124), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_132), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_154), .B(n_82), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_156), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
INVx8_ASAP7_75t_L g222 ( .A(n_138), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_142), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_142), .Y(n_224) );
AO22x2_ASAP7_75t_L g225 ( .A1(n_156), .A2(n_121), .B1(n_119), .B2(n_112), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_158), .B(n_107), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_158), .B(n_121), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_139), .Y(n_229) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_164), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_222), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_222), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_222), .B(n_164), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
AND3x2_ASAP7_75t_SL g236 ( .A(n_172), .B(n_167), .C(n_157), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_227), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_222), .B(n_164), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_190), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_172), .A2(n_164), .B1(n_85), .B2(n_110), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g241 ( .A1(n_191), .A2(n_123), .B1(n_141), .B2(n_137), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_176), .B(n_164), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_172), .A2(n_98), .B1(n_166), .B2(n_165), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_174), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_169), .B(n_159), .Y(n_247) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_163), .B(n_166), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_170), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_211), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_211), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_173), .B(n_159), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_186), .B(n_161), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_176), .B(n_137), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_191), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_178), .Y(n_256) );
INVx3_ASAP7_75t_SL g257 ( .A(n_168), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_174), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_172), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_227), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_202), .B(n_141), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_183), .B(n_160), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_225), .B(n_145), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_174), .Y(n_264) );
NOR3xp33_ASAP7_75t_L g265 ( .A(n_171), .B(n_145), .C(n_152), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_174), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_225), .A2(n_161), .B1(n_165), .B2(n_162), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_175), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_182), .Y(n_270) );
BUFx4f_ASAP7_75t_L g271 ( .A(n_214), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_170), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_217), .B(n_226), .Y(n_273) );
INVx5_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_194), .Y(n_275) );
BUFx12f_ASAP7_75t_L g276 ( .A(n_175), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_194), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_182), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_192), .B(n_162), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_225), .A2(n_163), .B1(n_160), .B2(n_152), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_212), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_168), .B(n_147), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_196), .B(n_198), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_212), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_220), .A2(n_147), .B1(n_163), .B2(n_146), .Y(n_287) );
AOI211xp5_ASAP7_75t_L g288 ( .A1(n_171), .A2(n_167), .B(n_157), .C(n_125), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_175), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_230), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_185), .B(n_163), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_183), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_203), .B(n_167), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_194), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_214), .B(n_157), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_201), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_201), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_262), .B(n_209), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_232), .B(n_230), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_262), .B(n_209), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_232), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_276), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_239), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g305 ( .A(n_232), .B(n_230), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_270), .B(n_193), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_262), .B(n_225), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_257), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_233), .B(n_195), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_259), .A2(n_214), .B1(n_195), .B2(n_197), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_232), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_254), .B(n_195), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_271), .A2(n_214), .B1(n_195), .B2(n_204), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_232), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g315 ( .A1(n_244), .A2(n_146), .B1(n_197), .B2(n_204), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_233), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_272), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_245), .B(n_197), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_254), .B(n_197), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_250), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_263), .A2(n_204), .B1(n_205), .B2(n_228), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_271), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_263), .Y(n_325) );
BUFx4f_ASAP7_75t_L g326 ( .A(n_234), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_259), .A2(n_205), .B1(n_204), .B2(n_208), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_248), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_234), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_257), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_272), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_273), .A2(n_253), .B(n_251), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_254), .B(n_205), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_292), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_260), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_260), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_250), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_290), .B(n_205), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_251), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_260), .B(n_206), .Y(n_340) );
NAND2x1_ASAP7_75t_SL g341 ( .A(n_240), .B(n_208), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_235), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_285), .B(n_206), .Y(n_343) );
OR2x6_ASAP7_75t_L g344 ( .A(n_263), .B(n_213), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_255), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_263), .A2(n_229), .B1(n_218), .B2(n_215), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_269), .A2(n_181), .B(n_177), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_278), .B(n_90), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_332), .A2(n_281), .B(n_267), .Y(n_349) );
NOR2x1_ASAP7_75t_SL g350 ( .A(n_344), .B(n_234), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_326), .A2(n_284), .B1(n_236), .B2(n_252), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_326), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_317), .A2(n_291), .B(n_293), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_329), .B(n_290), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_334), .B(n_284), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_323), .A2(n_241), .B1(n_265), .B2(n_242), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_323), .A2(n_288), .B(n_247), .C(n_242), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_326), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_345), .A2(n_261), .B1(n_234), .B2(n_238), .Y(n_359) );
OAI22xp5_ASAP7_75t_SL g360 ( .A1(n_330), .A2(n_236), .B1(n_261), .B2(n_238), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_315), .A2(n_242), .B1(n_238), .B2(n_261), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_343), .B(n_296), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_304), .A2(n_238), .B1(n_279), .B2(n_236), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_343), .B(n_246), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_322), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_329), .A2(n_290), .B1(n_297), .B2(n_295), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_344), .A2(n_266), .B1(n_258), .B2(n_264), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_301), .A2(n_136), .B1(n_126), .B2(n_133), .C(n_134), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_301), .B(n_296), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_317), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_SL g374 ( .A1(n_300), .A2(n_287), .B(n_297), .C(n_215), .Y(n_374) );
CKINVDCx14_ASAP7_75t_R g375 ( .A(n_330), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_344), .A2(n_268), .B1(n_289), .B2(n_280), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_298), .B(n_235), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_328), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_312), .B(n_235), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_371), .A2(n_348), .B1(n_306), .B2(n_364), .C(n_357), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_363), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_363), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_361), .A2(n_344), .B1(n_329), .B2(n_307), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_361), .A2(n_346), .B1(n_310), .B2(n_327), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_351), .A2(n_325), .B1(n_313), .B2(n_321), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_375), .Y(n_387) );
AOI33xp33_ASAP7_75t_L g388 ( .A1(n_359), .A2(n_126), .A3(n_125), .B1(n_143), .B2(n_136), .B3(n_133), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_379), .A2(n_347), .B(n_339), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_325), .B1(n_333), .B2(n_318), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_360), .A2(n_309), .B1(n_338), .B2(n_320), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_362), .B(n_340), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_356), .A2(n_299), .B1(n_318), .B2(n_308), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_144), .B(n_207), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_341), .B(n_303), .C(n_299), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_363), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_360), .A2(n_309), .B1(n_338), .B2(n_320), .Y(n_398) );
CKINVDCx11_ASAP7_75t_R g399 ( .A(n_376), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_355), .A2(n_309), .B1(n_338), .B2(n_320), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_355), .A2(n_341), .B1(n_324), .B2(n_308), .C(n_318), .Y(n_401) );
AOI222xp33_ASAP7_75t_L g402 ( .A1(n_365), .A2(n_339), .B1(n_337), .B2(n_324), .C1(n_269), .C2(n_282), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_370), .A2(n_305), .B1(n_316), .B2(n_336), .C(n_337), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_365), .A2(n_286), .B1(n_283), .B2(n_282), .C(n_229), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
BUFx4f_ASAP7_75t_SL g406 ( .A(n_376), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_349), .A2(n_286), .B1(n_283), .B2(n_218), .C(n_213), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_401), .A2(n_143), .B(n_134), .C(n_135), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_394), .B(n_352), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g411 ( .A1(n_396), .A2(n_370), .B(n_367), .C(n_352), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_392), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_373), .B(n_379), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_395), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_399), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_393), .B(n_362), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_386), .A2(n_372), .B1(n_349), .B2(n_369), .C(n_377), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_406), .A2(n_358), .B1(n_376), .B2(n_316), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_386), .A2(n_112), .B(n_119), .Y(n_420) );
OAI21x1_ASAP7_75t_L g421 ( .A1(n_389), .A2(n_379), .B(n_373), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_405), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_381), .A2(n_372), .B1(n_378), .B2(n_135), .C(n_374), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_385), .A2(n_378), .B1(n_135), .B2(n_380), .C(n_353), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_391), .A2(n_358), .B1(n_354), .B2(n_380), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_383), .B(n_382), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g428 ( .A1(n_405), .A2(n_144), .A3(n_181), .B1(n_177), .B2(n_180), .B3(n_188), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_383), .B(n_350), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_407), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_398), .A2(n_354), .B1(n_316), .B2(n_353), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_384), .A2(n_354), .B1(n_316), .B2(n_311), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_403), .A2(n_354), .B1(n_328), .B2(n_319), .Y(n_435) );
AOI221x1_ASAP7_75t_SL g436 ( .A1(n_390), .A2(n_144), .B1(n_148), .B2(n_8), .C(n_9), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_402), .A2(n_316), .B1(n_336), .B2(n_311), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_383), .B(n_368), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_402), .A2(n_311), .B1(n_302), .B2(n_319), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_382), .B(n_350), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_400), .A2(n_135), .B1(n_342), .B2(n_142), .C(n_335), .Y(n_441) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_382), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_404), .A2(n_302), .B1(n_331), .B2(n_335), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_417), .B(n_382), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_387), .B1(n_397), .B2(n_382), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_420), .A2(n_387), .B1(n_397), .B2(n_408), .Y(n_448) );
AND4x1_ASAP7_75t_L g449 ( .A(n_437), .B(n_418), .C(n_434), .D(n_388), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_412), .B(n_397), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_416), .B(n_397), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_422), .B(n_423), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_419), .B(n_397), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_422), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
OR2x2_ASAP7_75t_SL g456 ( .A(n_443), .B(n_395), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_423), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_429), .Y(n_458) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_443), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_436), .B(n_180), .C(n_184), .D(n_188), .Y(n_460) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_421), .A2(n_210), .B(n_207), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_429), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_429), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_431), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_425), .A2(n_305), .B1(n_335), .B2(n_342), .C(n_368), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_431), .B(n_368), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_426), .A2(n_368), .B1(n_328), .B2(n_305), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_440), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_433), .A2(n_331), .B1(n_314), .B2(n_328), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_432), .B(n_6), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_432), .B(n_7), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_424), .B(n_7), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
AOI21xp33_ASAP7_75t_SL g474 ( .A1(n_411), .A2(n_9), .B(n_10), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_414), .B(n_10), .Y(n_475) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_430), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_409), .A2(n_142), .B(n_84), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_413), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_441), .A2(n_314), .B1(n_328), .B2(n_342), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_440), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_439), .B(n_11), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_415), .B(n_87), .C(n_210), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_428), .A2(n_314), .B1(n_142), .B2(n_274), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_444), .A2(n_184), .B(n_200), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
OAI221xp5_ASAP7_75t_SL g490 ( .A1(n_438), .A2(n_12), .B1(n_13), .B2(n_14), .C(n_15), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_427), .B(n_17), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_427), .B(n_18), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_435), .A2(n_427), .B1(n_442), .B2(n_314), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_412), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_455), .B(n_19), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_468), .B(n_19), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_468), .B(n_21), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_483), .B(n_21), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_483), .B(n_23), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_445), .B(n_24), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_474), .A2(n_277), .B(n_274), .C(n_275), .Y(n_502) );
AOI31xp33_ASAP7_75t_L g503 ( .A1(n_474), .A2(n_25), .A3(n_27), .B(n_28), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_460), .B(n_207), .C(n_210), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_451), .B(n_30), .Y(n_505) );
NAND4xp25_ASAP7_75t_L g506 ( .A(n_490), .B(n_447), .C(n_448), .D(n_491), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_489), .B(n_216), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_446), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_489), .B(n_216), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_478), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_470), .B(n_216), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_445), .B(n_36), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_451), .B(n_37), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_485), .B(n_38), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_454), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_449), .B(n_41), .Y(n_517) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_461), .A2(n_221), .B(n_187), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_473), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_471), .B(n_189), .C(n_200), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_454), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_491), .B(n_42), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_470), .B(n_219), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_459), .B(n_45), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_492), .B(n_50), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_476), .B(n_51), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_475), .B(n_179), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_457), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_492), .B(n_52), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_457), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_464), .B(n_216), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_458), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_475), .A2(n_277), .B(n_274), .C(n_275), .Y(n_534) );
NAND4xp25_ASAP7_75t_L g535 ( .A(n_472), .B(n_189), .C(n_221), .D(n_223), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_467), .A2(n_274), .B1(n_224), .B2(n_178), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_473), .B(n_216), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_464), .Y(n_538) );
NOR2xp33_ASAP7_75t_R g539 ( .A(n_458), .B(n_55), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_453), .A2(n_294), .B(n_249), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_494), .B(n_224), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_477), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_494), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_466), .B(n_219), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_462), .B(n_57), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_462), .B(n_62), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_450), .B(n_219), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_463), .B(n_64), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_498), .B(n_463), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_506), .B(n_449), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_508), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_519), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_539), .B(n_481), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_495), .B(n_456), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_519), .B(n_456), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_533), .B(n_480), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_513), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_539), .B(n_480), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_516), .Y(n_561) );
OAI21xp33_ASAP7_75t_L g562 ( .A1(n_517), .A2(n_486), .B(n_493), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_501), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_544), .B(n_484), .Y(n_564) );
XNOR2xp5_ASAP7_75t_L g565 ( .A(n_522), .B(n_469), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_517), .B(n_465), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_533), .B(n_484), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_544), .B(n_461), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_521), .B(n_461), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_528), .B(n_482), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_496), .B(n_487), .C(n_488), .D(n_479), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_530), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_510), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_540), .B(n_223), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_515), .A2(n_219), .B1(n_224), .B2(n_178), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_538), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_540), .B(n_199), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_545), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_497), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_499), .B(n_65), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_540), .B(n_66), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_510), .B(n_179), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_512), .B(n_67), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_515), .A2(n_178), .B1(n_219), .B2(n_224), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_531), .B(n_68), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_503), .A2(n_274), .B(n_243), .C(n_237), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_543), .B(n_199), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_500), .B(n_256), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_542), .B(n_256), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_537), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_542), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_525), .B(n_256), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_256), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_507), .B(n_231), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_509), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_549), .B(n_231), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_555), .B(n_502), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_555), .A2(n_502), .B(n_534), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_560), .A2(n_524), .B1(n_550), .B2(n_548), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_553), .Y(n_602) );
XNOR2xp5_ASAP7_75t_L g603 ( .A(n_563), .B(n_514), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_552), .B(n_547), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_560), .B(n_526), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_586), .A2(n_534), .B(n_520), .C(n_504), .Y(n_607) );
NAND3x1_ASAP7_75t_SL g608 ( .A(n_583), .B(n_504), .C(n_520), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_561), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_572), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_557), .B(n_546), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_551), .B(n_558), .Y(n_612) );
AOI21x1_ASAP7_75t_L g613 ( .A1(n_590), .A2(n_511), .B(n_523), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_576), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_556), .B(n_536), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_578), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_556), .B(n_536), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_554), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_592), .B(n_518), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_552), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_592), .B(n_518), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_579), .B(n_505), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_573), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_573), .B(n_541), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_566), .B(n_535), .Y(n_626) );
XNOR2x2_ASAP7_75t_L g627 ( .A(n_566), .B(n_249), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_597), .B(n_294), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_586), .B(n_256), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_588), .B(n_237), .Y(n_630) );
NOR2xp33_ASAP7_75t_SL g631 ( .A(n_562), .B(n_237), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_593), .B(n_567), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_568), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_580), .B(n_243), .C(n_571), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_595), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_570), .B(n_243), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_569), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_567), .B(n_587), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_565), .A2(n_580), .B1(n_575), .B2(n_584), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_582), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_585), .A2(n_598), .B1(n_581), .B2(n_594), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_585), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_574), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_577), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_596), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_591), .Y(n_648) );
OA21x2_ASAP7_75t_L g649 ( .A1(n_589), .A2(n_569), .B(n_481), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_589), .Y(n_650) );
OAI21xp33_ASAP7_75t_SL g651 ( .A1(n_594), .A2(n_555), .B(n_560), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_563), .B(n_415), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_555), .B(n_560), .Y(n_653) );
AOI321xp33_ASAP7_75t_L g654 ( .A1(n_626), .A2(n_605), .A3(n_653), .B1(n_641), .B2(n_615), .C(n_617), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_620), .A2(n_603), .B1(n_607), .B2(n_652), .Y(n_655) );
AOI331xp33_ASAP7_75t_L g656 ( .A1(n_626), .A2(n_605), .A3(n_652), .B1(n_634), .B2(n_602), .B3(n_604), .C1(n_616), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_629), .A2(n_651), .B(n_599), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_629), .A2(n_651), .B(n_599), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_633), .Y(n_659) );
AOI211xp5_ASAP7_75t_SL g660 ( .A1(n_631), .A2(n_607), .B(n_600), .C(n_643), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_635), .A2(n_611), .B1(n_627), .B2(n_650), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_634), .B(n_639), .Y(n_662) );
AOI221x1_ASAP7_75t_L g663 ( .A1(n_635), .A2(n_618), .B1(n_621), .B2(n_639), .C(n_610), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_606), .A2(n_601), .B1(n_636), .B2(n_623), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_640), .A2(n_636), .B(n_606), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_624), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_636), .A2(n_650), .B1(n_613), .B2(n_648), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_655), .A2(n_611), .B1(n_627), .B2(n_647), .Y(n_668) );
INVxp67_ASAP7_75t_SL g669 ( .A(n_657), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_664), .B(n_608), .C(n_638), .Y(n_670) );
AOI211x1_ASAP7_75t_SL g671 ( .A1(n_658), .A2(n_608), .B(n_630), .C(n_646), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_664), .B(n_614), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_654), .Y(n_673) );
OAI22xp5_ASAP7_75t_SL g674 ( .A1(n_661), .A2(n_649), .B1(n_644), .B2(n_637), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g675 ( .A1(n_660), .A2(n_609), .B(n_647), .C(n_628), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_673), .A2(n_667), .B1(n_659), .B2(n_665), .C(n_662), .Y(n_676) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_669), .B(n_667), .C(n_656), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_672), .B(n_663), .C(n_666), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_668), .B(n_611), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_679), .Y(n_680) );
OAI222xp33_ASAP7_75t_L g681 ( .A1(n_677), .A2(n_675), .B1(n_671), .B2(n_674), .C1(n_670), .C2(n_632), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g682 ( .A1(n_676), .A2(n_645), .B(n_649), .C(n_622), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_681), .A2(n_678), .B(n_649), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_680), .A2(n_649), .B1(n_645), .B2(n_644), .C(n_642), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_683), .A2(n_682), .B1(n_622), .B2(n_619), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_685), .Y(n_686) );
AOI22x1_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_684), .B1(n_632), .B2(n_612), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_642), .B1(n_619), .B2(n_625), .C(n_646), .Y(n_688) );
endmodule