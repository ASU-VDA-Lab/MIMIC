module fake_jpeg_21612_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_22),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_25),
.B1(n_21),
.B2(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_21),
.B1(n_25),
.B2(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_25),
.B1(n_38),
.B2(n_30),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_70),
.B1(n_65),
.B2(n_27),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_39),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_71),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_16),
.B1(n_30),
.B2(n_17),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_33),
.B1(n_24),
.B2(n_17),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_76),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_74),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_79),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_33),
.B1(n_16),
.B2(n_30),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_91),
.B1(n_15),
.B2(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_109),
.B1(n_56),
.B2(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_20),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_20),
.B(n_18),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_18),
.B1(n_15),
.B2(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_83),
.Y(n_136)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_31),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_71),
.C(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_56),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_114),
.B(n_122),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_140),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_61),
.C(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_23),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_59),
.B1(n_79),
.B2(n_69),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_141),
.B1(n_0),
.B2(n_1),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_22),
.B(n_31),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_111),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_14),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_13),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_0),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_86),
.B1(n_96),
.B2(n_85),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_106),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_139),
.Y(n_151)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_56),
.B1(n_22),
.B2(n_14),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_99),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_125),
.C(n_122),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_100),
.B(n_101),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_150),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_93),
.B1(n_102),
.B2(n_112),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_164),
.B1(n_141),
.B2(n_165),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_148),
.A2(n_155),
.B(n_156),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_1),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_98),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_111),
.B(n_103),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_91),
.A3(n_85),
.B1(n_96),
.B2(n_109),
.C1(n_103),
.C2(n_31),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_3),
.B(n_4),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_162),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_86),
.C(n_22),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_94),
.B1(n_88),
.B2(n_95),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_169),
.B1(n_171),
.B2(n_128),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_95),
.B(n_88),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_4),
.B(n_5),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_0),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_12),
.B1(n_13),
.B2(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_180),
.B1(n_183),
.B2(n_194),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_142),
.Y(n_206)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_191),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_187),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_119),
.B(n_118),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_204),
.B(n_168),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_118),
.B(n_120),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_182),
.A2(n_198),
.B(n_146),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_140),
.B1(n_120),
.B2(n_2),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_184),
.A2(n_201),
.B1(n_203),
.B2(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_153),
.B(n_3),
.Y(n_195)
);

XOR2x2_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_144),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_5),
.C(n_6),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_195),
.C(n_169),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_167),
.B1(n_156),
.B2(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_5),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_144),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_7),
.B(n_8),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_172),
.B(n_7),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_188),
.C(n_175),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_203),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_224),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_160),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_228),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_143),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_159),
.B1(n_145),
.B2(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_225),
.B1(n_178),
.B2(n_201),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_204),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_145),
.B1(n_163),
.B2(n_170),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_148),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_245),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_224),
.B1(n_216),
.B2(n_189),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_237),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_199),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_197),
.C(n_146),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_244),
.C(n_183),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_182),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_189),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_197),
.C(n_176),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_213),
.B(n_228),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_223),
.B(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_244),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_250),
.B(n_238),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_231),
.A2(n_216),
.B1(n_207),
.B2(n_179),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_254),
.B1(n_247),
.B2(n_234),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_184),
.B1(n_193),
.B2(n_227),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_149),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_187),
.B(n_209),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_262),
.B(n_219),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_212),
.C(n_221),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_241),
.C(n_242),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_196),
.B(n_194),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_269),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_257),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_270),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_273),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_222),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_8),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_263),
.B1(n_251),
.B2(n_10),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_260),
.C(n_258),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_286),
.C(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_268),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_260),
.C(n_258),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_272),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_248),
.B1(n_262),
.B2(n_274),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_249),
.B(n_261),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_261),
.B(n_9),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_10),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_286),
.C(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_297),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_289),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.C(n_300),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_303),
.B(n_302),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_292),
.C(n_291),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_285),
.B(n_299),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_311),
.Y(n_312)
);


endmodule