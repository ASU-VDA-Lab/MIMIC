module fake_netlist_1_6665_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_SL g13 ( .A(n_9), .Y(n_13) );
INVx8_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
BUFx10_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
NAND2x1p5_ASAP7_75t_L g18 ( .A(n_16), .B(n_0), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_15), .B(n_1), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_19), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
INVx2_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
OAI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_13), .B1(n_17), .B2(n_14), .C(n_5), .Y(n_23) );
INVx3_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
OAI22xp5_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_6), .B1(n_11), .B2(n_12), .Y(n_26) );
endmodule