module fake_netlist_1_8658_n_949 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_191, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_949);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_949;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_918;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_881;
wire n_806;
wire n_539;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_948;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_912;
wire n_924;
wire n_841;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g200 ( .A(n_176), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_192), .B(n_191), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_188), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_110), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_3), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_98), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_73), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_100), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_127), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_43), .Y(n_210) );
INVxp67_ASAP7_75t_SL g211 ( .A(n_138), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
INVx1_ASAP7_75t_SL g213 ( .A(n_131), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_36), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_78), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_183), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_51), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_50), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_76), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_121), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_122), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_175), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_144), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_142), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_113), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_48), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_152), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_47), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_91), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_12), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_177), .Y(n_232) );
INVxp33_ASAP7_75t_L g233 ( .A(n_66), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_143), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_48), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_159), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_197), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_186), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_182), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_5), .Y(n_241) );
BUFx5_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_155), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_59), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_115), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_162), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_189), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_193), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_42), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_88), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_154), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_118), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g253 ( .A(n_111), .B(n_151), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_160), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_15), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_4), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_95), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_180), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_24), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_109), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_82), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_73), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_80), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_47), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_168), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_77), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_119), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_93), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_116), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_120), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_147), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_139), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_146), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_198), .Y(n_274) );
INVxp33_ASAP7_75t_L g275 ( .A(n_199), .Y(n_275) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_157), .B(n_148), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_59), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_114), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_87), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_105), .Y(n_280) );
INVxp33_ASAP7_75t_SL g281 ( .A(n_24), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_125), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_169), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_170), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_45), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_108), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_129), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_171), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_15), .Y(n_289) );
CKINVDCx16_ASAP7_75t_R g290 ( .A(n_51), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_117), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_46), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_134), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_174), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_167), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_2), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_28), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_123), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_153), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_82), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_22), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_164), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_173), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_156), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_172), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_150), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_94), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_68), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_13), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_140), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_106), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_136), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_5), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_36), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_50), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_149), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_230), .B(n_0), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_241), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_274), .B(n_0), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_242), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_231), .B(n_1), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_241), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_315), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_233), .B(n_1), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_231), .B(n_3), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_226), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_261), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_200), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_245), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_242), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_202), .Y(n_334) );
NOR2x1_ASAP7_75t_L g335 ( .A(n_206), .B(n_4), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_281), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_245), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_209), .Y(n_338) );
OAI22xp5_ASAP7_75t_SL g339 ( .A1(n_235), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g340 ( .A(n_242), .B(n_85), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_212), .Y(n_341) );
NOR2x1_ASAP7_75t_L g342 ( .A(n_216), .B(n_9), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_242), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_233), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_242), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_275), .B(n_9), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_247), .B(n_10), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_221), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_208), .A2(n_89), .B(n_86), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_242), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_255), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_344), .B(n_243), .Y(n_352) );
INVx4_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_344), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_351), .B(n_275), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_331), .B(n_222), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_324), .B(n_290), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
INVx5_ASAP7_75t_L g364 ( .A(n_332), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_346), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
NAND2xp33_ASAP7_75t_L g367 ( .A(n_346), .B(n_204), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_331), .B(n_203), .Y(n_368) );
INVx6_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
NAND3xp33_ASAP7_75t_L g370 ( .A(n_340), .B(n_224), .C(n_223), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_334), .B(n_255), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_329), .A2(n_297), .B1(n_281), .B2(n_240), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_325), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
NAND2xp33_ASAP7_75t_L g375 ( .A(n_338), .B(n_228), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_338), .B(n_237), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_341), .B(n_237), .Y(n_377) );
AND3x2_ASAP7_75t_L g378 ( .A(n_324), .B(n_286), .C(n_211), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_341), .B(n_262), .Y(n_380) );
NAND2xp33_ASAP7_75t_L g381 ( .A(n_348), .B(n_234), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_332), .Y(n_382) );
BUFx10_ASAP7_75t_L g383 ( .A(n_325), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_333), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_332), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_333), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_333), .Y(n_387) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_325), .B(n_208), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_348), .B(n_262), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_328), .B(n_251), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_317), .B(n_285), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_343), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_325), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_339), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_317), .A2(n_215), .B1(n_217), .B2(n_214), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_354), .B(n_319), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_365), .B(n_335), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_360), .B(n_319), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_354), .A2(n_240), .B1(n_252), .B2(n_225), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_365), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_392), .Y(n_404) );
O2A1O1Ixp5_ASAP7_75t_L g405 ( .A1(n_353), .A2(n_347), .B(n_330), .C(n_328), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_392), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_356), .B(n_285), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_371), .B(n_347), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_388), .A2(n_345), .B1(n_350), .B2(n_330), .Y(n_409) );
NOR2x1p5_ASAP7_75t_L g410 ( .A(n_360), .B(n_292), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_388), .A2(n_349), .B(n_345), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_252), .B1(n_295), .B2(n_225), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_352), .A2(n_299), .B1(n_295), .B2(n_339), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_369), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_380), .B(n_268), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_389), .B(n_268), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_368), .B(n_273), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_383), .B(n_350), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_359), .A2(n_349), .B(n_350), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_353), .B(n_273), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_373), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_383), .B(n_357), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_357), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_358), .B(n_318), .Y(n_426) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_357), .B(n_235), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_361), .B(n_232), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_362), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_372), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_396), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g434 ( .A1(n_367), .A2(n_322), .B(n_323), .C(n_318), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_361), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_397), .A2(n_314), .B1(n_336), .B2(n_308), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_395), .A2(n_342), .B1(n_335), .B2(n_323), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_376), .B(n_229), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_395), .A2(n_342), .B1(n_327), .B2(n_322), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_377), .B(n_327), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_390), .B(n_218), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_375), .B(n_264), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_359), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_381), .B(n_278), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_362), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_363), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_370), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_374), .B(n_283), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_379), .B(n_283), .Y(n_450) );
BUFx5_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_384), .B(n_284), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_384), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_386), .B(n_236), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_386), .A2(n_227), .B1(n_244), .B2(n_219), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_387), .B(n_238), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_387), .B(n_284), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_393), .B(n_296), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_393), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_394), .A2(n_256), .B1(n_259), .B2(n_249), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_394), .B(n_263), .Y(n_461) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_391), .B(n_349), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_382), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_364), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_364), .B(n_293), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_382), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_382), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_391), .A2(n_220), .B(n_304), .C(n_246), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_364), .B(n_293), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_366), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_366), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_366), .A2(n_277), .B1(n_289), .B2(n_266), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_366), .B(n_294), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_366), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_451), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_411), .A2(n_349), .B(n_201), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_409), .A2(n_301), .B1(n_309), .B2(n_300), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_404), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_409), .A2(n_313), .B1(n_257), .B2(n_258), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_451), .B(n_239), .Y(n_480) );
INVxp33_ASAP7_75t_SL g481 ( .A(n_401), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_400), .B(n_265), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_420), .A2(n_269), .B(n_267), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_427), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_408), .A2(n_271), .B(n_272), .C(n_270), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_403), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_407), .B(n_213), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_420), .A2(n_280), .B(n_279), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_414), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_399), .B(n_282), .Y(n_490) );
INVx3_ASAP7_75t_SL g491 ( .A(n_427), .Y(n_491) );
OR2x6_ASAP7_75t_SL g492 ( .A(n_433), .B(n_250), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_424), .A2(n_288), .B(n_287), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_399), .B(n_254), .Y(n_494) );
OAI21x1_ASAP7_75t_L g495 ( .A1(n_421), .A2(n_246), .B(n_220), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_424), .A2(n_298), .B(n_291), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_458), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_414), .Y(n_498) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_468), .A2(n_303), .B(n_302), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_410), .A2(n_306), .B1(n_310), .B2(n_305), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_451), .B(n_311), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_428), .A2(n_312), .B(n_276), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_435), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_405), .A2(n_253), .B(n_260), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_413), .B(n_10), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_461), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_442), .B(n_205), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_412), .B(n_11), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_428), .A2(n_316), .B(n_385), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_435), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_448), .A2(n_205), .B(n_207), .C(n_210), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_459), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_432), .B(n_210), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_440), .A2(n_385), .B(n_248), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_459), .B(n_245), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_422), .A2(n_385), .B(n_307), .Y(n_517) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_425), .B(n_307), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_439), .A2(n_337), .B1(n_12), .B2(n_13), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_415), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_417), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_438), .B(n_11), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_439), .B(n_14), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_442), .A2(n_16), .B(n_17), .C(n_18), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_426), .A2(n_337), .B(n_17), .C(n_18), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_443), .B(n_16), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_472), .A2(n_19), .B(n_20), .C(n_21), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_416), .A2(n_337), .B(n_90), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_452), .B(n_19), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_418), .A2(n_337), .B(n_92), .Y(n_530) );
INVx5_ASAP7_75t_L g531 ( .A(n_402), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_454), .A2(n_20), .B(n_21), .C(n_22), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_444), .B(n_23), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_454), .A2(n_23), .B(n_25), .C(n_26), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_436), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_449), .B(n_27), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_441), .B(n_29), .Y(n_537) );
AO22x1_ASAP7_75t_L g538 ( .A1(n_433), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_450), .A2(n_97), .B(n_96), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_447), .A2(n_30), .B(n_31), .C(n_32), .Y(n_540) );
O2A1O1Ixp5_ASAP7_75t_L g541 ( .A1(n_456), .A2(n_124), .B(n_196), .C(n_195), .Y(n_541) );
OAI22x1_ASAP7_75t_L g542 ( .A1(n_455), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_457), .A2(n_101), .B(n_99), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_419), .B(n_33), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_402), .Y(n_545) );
AOI22x1_ASAP7_75t_L g546 ( .A1(n_453), .A2(n_126), .B1(n_194), .B2(n_190), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_437), .B(n_34), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_445), .B(n_423), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_430), .A2(n_103), .B(n_102), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_460), .B(n_35), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_437), .B(n_35), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_464), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_429), .A2(n_446), .B(n_473), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_460), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_456), .B(n_37), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_465), .B(n_39), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_463), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_469), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_467), .B(n_40), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_471), .A2(n_128), .B(n_187), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_468), .A2(n_40), .B(n_41), .C(n_42), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g562 ( .A1(n_466), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g563 ( .A1(n_470), .A2(n_44), .B1(n_46), .B2(n_49), .C(n_52), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_474), .A2(n_133), .B(n_185), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_403), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_403), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_403), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_411), .A2(n_135), .B(n_184), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_411), .A2(n_132), .B(n_181), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_398), .B(n_53), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_400), .A2(n_54), .B(n_55), .C(n_56), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_411), .A2(n_137), .B(n_179), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_435), .Y(n_573) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_462), .A2(n_130), .B(n_178), .Y(n_574) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_513), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_491), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_576) );
INVx6_ASAP7_75t_SL g577 ( .A(n_526), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_486), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_508), .A2(n_500), .B1(n_497), .B2(n_535), .C(n_478), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_565), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_503), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_481), .B(n_57), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_566), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_492), .Y(n_585) );
BUFx2_ASAP7_75t_R g586 ( .A(n_484), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_545), .Y(n_587) );
BUFx12f_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_477), .B(n_58), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_487), .A2(n_60), .B(n_61), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_567), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_477), .A2(n_62), .B1(n_63), .B2(n_64), .C(n_65), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_554), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_504), .A2(n_145), .B(n_163), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_505), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_533), .Y(n_596) );
AO32x2_ASAP7_75t_L g597 ( .A1(n_479), .A2(n_67), .A3(n_69), .B1(n_70), .B2(n_71), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_475), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_538), .Y(n_599) );
AO31x2_ASAP7_75t_L g600 ( .A1(n_561), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_522), .A2(n_72), .B(n_74), .C(n_75), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_482), .B(n_72), .Y(n_602) );
NOR2xp33_ASAP7_75t_SL g603 ( .A(n_552), .B(n_74), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_548), .A2(n_75), .B(n_76), .C(n_77), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_531), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_562), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_490), .B(n_79), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_533), .Y(n_608) );
O2A1O1Ixp5_ASAP7_75t_L g609 ( .A1(n_504), .A2(n_536), .B(n_517), .C(n_529), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_570), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_552), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_545), .A2(n_80), .B1(n_81), .B2(n_83), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_503), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_501), .A2(n_84), .B1(n_104), .B2(n_107), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_550), .B(n_112), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_555), .Y(n_616) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_503), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_519), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_512), .B(n_531), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_494), .B(n_479), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_485), .B(n_551), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_SL g622 ( .A1(n_525), .A2(n_511), .B(n_559), .C(n_569), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_551), .A2(n_547), .B1(n_523), .B2(n_537), .Y(n_623) );
AO32x2_ASAP7_75t_L g624 ( .A1(n_558), .A2(n_499), .A3(n_542), .B1(n_524), .B2(n_527), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_531), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_507), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_540), .A2(n_532), .B(n_534), .C(n_514), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_557), .B(n_520), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_518), .A2(n_480), .B(n_515), .Y(n_629) );
AO31x2_ASAP7_75t_L g630 ( .A1(n_572), .A2(n_516), .A3(n_528), .B(n_530), .Y(n_630) );
AO31x2_ASAP7_75t_L g631 ( .A1(n_539), .A2(n_543), .A3(n_502), .B(n_549), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_521), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_563), .A2(n_496), .B1(n_493), .B2(n_483), .C(n_488), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_556), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_SL g635 ( .A1(n_560), .A2(n_509), .B(n_564), .C(n_573), .Y(n_635) );
INVx4_ASAP7_75t_L g636 ( .A(n_489), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_510), .Y(n_637) );
AO31x2_ASAP7_75t_L g638 ( .A1(n_499), .A2(n_546), .A3(n_541), .B(n_498), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_506), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_476), .A2(n_553), .B(n_411), .Y(n_640) );
BUFx3_ASAP7_75t_L g641 ( .A(n_491), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_476), .A2(n_411), .B(n_405), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_506), .B(n_406), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_506), .B(n_404), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_481), .A2(n_427), .B1(n_484), .B2(n_477), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_475), .Y(n_646) );
BUFx12f_ASAP7_75t_L g647 ( .A(n_478), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_506), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_497), .A2(n_406), .B1(n_431), .B2(n_413), .C(n_400), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_506), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_506), .B(n_406), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_476), .A2(n_553), .B(n_411), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_497), .A2(n_431), .B1(n_404), .B2(n_477), .C(n_354), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_485), .A2(n_571), .B(n_431), .C(n_404), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_548), .A2(n_544), .B(n_434), .C(n_571), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_478), .B(n_404), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_548), .A2(n_544), .B(n_434), .C(n_571), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_495), .A2(n_574), .B(n_462), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_548), .A2(n_544), .B(n_434), .C(n_571), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_481), .A2(n_412), .B1(n_401), .B2(n_427), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_491), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_506), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_491), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_545), .Y(n_664) );
AO32x2_ASAP7_75t_L g665 ( .A1(n_479), .A2(n_519), .A3(n_554), .B1(n_562), .B2(n_477), .Y(n_665) );
BUFx8_ASAP7_75t_SL g666 ( .A(n_478), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_478), .B(n_404), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_478), .Y(n_668) );
AOI22xp5_ASAP7_75t_SL g669 ( .A1(n_481), .A2(n_396), .B1(n_296), .B2(n_301), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_506), .B(n_404), .Y(n_670) );
INVx5_ASAP7_75t_L g671 ( .A(n_475), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_481), .B(n_431), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_506), .B(n_404), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_476), .A2(n_553), .B(n_411), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_476), .A2(n_553), .B(n_411), .Y(n_675) );
AO21x1_ASAP7_75t_L g676 ( .A1(n_568), .A2(n_572), .B(n_569), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_640), .A2(n_674), .B(n_652), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_649), .A2(n_653), .B1(n_580), .B2(n_672), .C(n_654), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_601), .B(n_657), .C(n_655), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_578), .B(n_639), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_628), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_675), .A2(n_635), .B(n_642), .Y(n_682) );
OR2x6_ASAP7_75t_L g683 ( .A(n_588), .B(n_641), .Y(n_683) );
NAND2x1p5_ASAP7_75t_L g684 ( .A(n_671), .B(n_619), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_647), .Y(n_685) );
INVxp33_ASAP7_75t_L g686 ( .A(n_666), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_620), .A2(n_659), .B(n_627), .C(n_621), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_622), .A2(n_629), .B(n_676), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_625), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_671), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_648), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_623), .A2(n_596), .B(n_608), .C(n_610), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_579), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_645), .B(n_671), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_618), .A2(n_589), .B1(n_575), .B2(n_602), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_590), .A2(n_583), .B(n_603), .Y(n_696) );
OR2x6_ASAP7_75t_L g697 ( .A(n_661), .B(n_663), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_609), .A2(n_634), .B(n_604), .C(n_633), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_650), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_581), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_662), .B(n_616), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g702 ( .A1(n_660), .A2(n_644), .B(n_673), .C(n_670), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_656), .B(n_667), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_584), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_592), .A2(n_595), .B(n_615), .C(n_626), .Y(n_705) );
AND2x6_ASAP7_75t_L g706 ( .A(n_619), .B(n_598), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_591), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_643), .B(n_651), .Y(n_708) );
AO22x1_ASAP7_75t_L g709 ( .A1(n_585), .A2(n_599), .B1(n_606), .B2(n_668), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_587), .A2(n_664), .B1(n_577), .B2(n_593), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g711 ( .A(n_605), .B(n_646), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_582), .Y(n_712) );
INVx4_ASAP7_75t_L g713 ( .A(n_582), .Y(n_713) );
AND2x4_ASAP7_75t_L g714 ( .A(n_611), .B(n_632), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_637), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_586), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_607), .A2(n_576), .B(n_612), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_669), .B(n_577), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_600), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_597), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_636), .B(n_600), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_624), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_665), .A2(n_624), .B1(n_613), .B2(n_617), .C(n_597), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_613), .B(n_631), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_631), .B(n_630), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_631), .A2(n_630), .B(n_638), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_628), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_672), .A2(n_481), .B1(n_645), .B2(n_620), .Y(n_728) );
AO21x1_ASAP7_75t_L g729 ( .A1(n_594), .A2(n_614), .B(n_601), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_645), .B(n_671), .Y(n_730) );
INVx1_ASAP7_75t_SL g731 ( .A(n_625), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_620), .A2(n_657), .B(n_659), .C(n_655), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_668), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_645), .A2(n_660), .B1(n_580), .B2(n_672), .C(n_649), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_596), .B(n_608), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_640), .A2(n_675), .B(n_674), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_620), .A2(n_657), .B(n_659), .C(n_655), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_656), .B(n_667), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_578), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_672), .A2(n_481), .B1(n_645), .B2(n_620), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_643), .B(n_404), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_672), .B(n_481), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_578), .Y(n_743) );
OA21x2_ASAP7_75t_L g744 ( .A1(n_658), .A2(n_495), .B(n_640), .Y(n_744) );
INVx4_ASAP7_75t_L g745 ( .A(n_641), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_578), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_640), .A2(n_675), .B(n_674), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_640), .A2(n_675), .B(n_674), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_671), .B(n_619), .Y(n_749) );
AOI222xp33_ASAP7_75t_L g750 ( .A1(n_672), .A2(n_339), .B1(n_481), .B2(n_653), .C1(n_396), .C2(n_606), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_596), .B(n_608), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g752 ( .A1(n_642), .A2(n_623), .B(n_674), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_640), .A2(n_675), .B(n_674), .Y(n_753) );
OR2x2_ASAP7_75t_L g754 ( .A(n_656), .B(n_667), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_672), .A2(n_481), .B1(n_645), .B2(n_620), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_578), .Y(n_756) );
OR2x6_ASAP7_75t_L g757 ( .A(n_588), .B(n_641), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_666), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_653), .B(n_404), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_640), .A2(n_675), .B(n_674), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_578), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_653), .B(n_404), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_653), .B(n_404), .Y(n_763) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_658), .A2(n_495), .B(n_640), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_628), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_653), .B(n_404), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_660), .A2(n_412), .B1(n_401), .B2(n_413), .Y(n_767) );
BUFx2_ASAP7_75t_L g768 ( .A(n_647), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_726), .A2(n_688), .B(n_682), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_681), .B(n_727), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_734), .A2(n_710), .B1(n_695), .B2(n_679), .Y(n_771) );
OA21x2_ASAP7_75t_L g772 ( .A1(n_677), .A2(n_747), .B(n_736), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g773 ( .A1(n_705), .A2(n_679), .B(n_692), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_765), .B(n_703), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_735), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_706), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_732), .B(n_737), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_702), .A2(n_678), .B1(n_750), .B2(n_728), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_698), .A2(n_687), .B(n_717), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_767), .A2(n_759), .B1(n_766), .B2(n_763), .C(n_762), .Y(n_780) );
AND2x4_ASAP7_75t_SL g781 ( .A(n_749), .B(n_690), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_751), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_749), .B(n_752), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_751), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_738), .B(n_754), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_693), .B(n_700), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_720), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_715), .B(n_704), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_707), .B(n_691), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_719), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_695), .B(n_708), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_699), .B(n_739), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_725), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_743), .B(n_746), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_725), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_721), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_756), .Y(n_797) );
OR2x6_ASAP7_75t_L g798 ( .A(n_694), .B(n_730), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_761), .Y(n_799) );
OA21x2_ASAP7_75t_L g800 ( .A1(n_748), .A2(n_753), .B(n_760), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_701), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_724), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_680), .Y(n_803) );
INVxp67_ASAP7_75t_L g804 ( .A(n_741), .Y(n_804) );
OAI211xp5_ASAP7_75t_L g805 ( .A1(n_750), .A2(n_755), .B(n_740), .C(n_696), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_684), .B(n_711), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_710), .B(n_733), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_706), .Y(n_808) );
INVxp67_ASAP7_75t_L g809 ( .A(n_718), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_742), .A2(n_717), .B1(n_696), .B2(n_729), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_722), .B(n_706), .Y(n_811) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_731), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_689), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_723), .Y(n_814) );
INVx3_ASAP7_75t_SL g815 ( .A(n_683), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_744), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_731), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_714), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_714), .B(n_709), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_713), .B(n_712), .Y(n_820) );
INVxp67_ASAP7_75t_L g821 ( .A(n_768), .Y(n_821) );
NOR2xp33_ASAP7_75t_SL g822 ( .A(n_758), .B(n_716), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_764), .B(n_716), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_697), .A2(n_683), .B1(n_757), .B2(n_685), .Y(n_824) );
BUFx3_ASAP7_75t_L g825 ( .A(n_697), .Y(n_825) );
CKINVDCx6p67_ASAP7_75t_R g826 ( .A(n_683), .Y(n_826) );
OR2x2_ASAP7_75t_L g827 ( .A(n_697), .B(n_745), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_802), .B(n_745), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_802), .B(n_757), .Y(n_829) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_816), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_787), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_793), .B(n_686), .Y(n_832) );
OR2x6_ASAP7_75t_L g833 ( .A(n_776), .B(n_808), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_795), .B(n_796), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_791), .B(n_795), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_783), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_778), .A2(n_771), .B1(n_780), .B2(n_777), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_783), .B(n_796), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_790), .Y(n_839) );
AND2x4_ASAP7_75t_L g840 ( .A(n_783), .B(n_811), .Y(n_840) );
INVx5_ASAP7_75t_SL g841 ( .A(n_826), .Y(n_841) );
INVx2_ASAP7_75t_SL g842 ( .A(n_781), .Y(n_842) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_825), .B(n_827), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_783), .B(n_786), .Y(n_844) );
AND2x4_ASAP7_75t_L g845 ( .A(n_811), .B(n_823), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_805), .B(n_821), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_804), .B(n_809), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_791), .B(n_785), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_786), .B(n_789), .Y(n_849) );
INVx1_ASAP7_75t_SL g850 ( .A(n_820), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_789), .B(n_792), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_792), .B(n_794), .Y(n_852) );
BUFx2_ASAP7_75t_L g853 ( .A(n_798), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_807), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_794), .B(n_788), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_775), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_788), .B(n_814), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_814), .B(n_777), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_782), .Y(n_859) );
INVx1_ASAP7_75t_SL g860 ( .A(n_820), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_797), .B(n_799), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_834), .B(n_801), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_834), .B(n_801), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_831), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_848), .B(n_800), .Y(n_865) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_839), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_854), .B(n_800), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_854), .B(n_800), .Y(n_868) );
OR2x2_ASAP7_75t_L g869 ( .A(n_835), .B(n_800), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_845), .B(n_769), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_845), .B(n_769), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_844), .B(n_769), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g873 ( .A(n_846), .B(n_773), .C(n_779), .Y(n_873) );
INVx1_ASAP7_75t_SL g874 ( .A(n_850), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_844), .B(n_769), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_838), .B(n_772), .Y(n_876) );
INVx1_ASAP7_75t_SL g877 ( .A(n_850), .Y(n_877) );
INVx2_ASAP7_75t_SL g878 ( .A(n_843), .Y(n_878) );
NOR2xp67_ASAP7_75t_L g879 ( .A(n_828), .B(n_827), .Y(n_879) );
BUFx2_ASAP7_75t_L g880 ( .A(n_843), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_856), .B(n_784), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_856), .B(n_803), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_873), .A2(n_837), .B1(n_858), .B2(n_810), .C(n_832), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_872), .B(n_836), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_872), .B(n_840), .Y(n_885) );
INVx1_ASAP7_75t_SL g886 ( .A(n_874), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_864), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_864), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_862), .B(n_851), .Y(n_889) );
NOR3xp33_ASAP7_75t_L g890 ( .A(n_873), .B(n_819), .C(n_832), .Y(n_890) );
NOR2x1_ASAP7_75t_L g891 ( .A(n_879), .B(n_828), .Y(n_891) );
AND2x4_ASAP7_75t_L g892 ( .A(n_870), .B(n_871), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_875), .B(n_852), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_862), .B(n_852), .Y(n_894) );
AND2x4_ASAP7_75t_L g895 ( .A(n_870), .B(n_853), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_863), .B(n_822), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_866), .A2(n_830), .B(n_842), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_865), .B(n_860), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_875), .B(n_855), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_882), .B(n_849), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_865), .B(n_859), .Y(n_901) );
INVx3_ASAP7_75t_L g902 ( .A(n_892), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_887), .Y(n_903) );
OAI21xp33_ASAP7_75t_L g904 ( .A1(n_891), .A2(n_877), .B(n_847), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_893), .B(n_869), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_888), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_892), .B(n_870), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_892), .B(n_871), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_899), .B(n_861), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_899), .B(n_861), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_888), .Y(n_911) );
OR2x2_ASAP7_75t_L g912 ( .A(n_898), .B(n_869), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_898), .B(n_869), .Y(n_913) );
OAI32xp33_ASAP7_75t_L g914 ( .A1(n_890), .A2(n_829), .A3(n_817), .B1(n_812), .B2(n_881), .Y(n_914) );
INVxp67_ASAP7_75t_L g915 ( .A(n_896), .Y(n_915) );
NOR2xp67_ASAP7_75t_L g916 ( .A(n_897), .B(n_878), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_885), .B(n_876), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_912), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_912), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_904), .A2(n_883), .B1(n_895), .B2(n_884), .Y(n_920) );
HB1xp67_ASAP7_75t_L g921 ( .A(n_913), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_914), .A2(n_878), .B(n_901), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_913), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_914), .A2(n_901), .B(n_880), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_905), .B(n_886), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_903), .Y(n_926) );
INVxp67_ASAP7_75t_L g927 ( .A(n_915), .Y(n_927) );
INVxp67_ASAP7_75t_L g928 ( .A(n_927), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_920), .A2(n_902), .B1(n_916), .B2(n_908), .Y(n_929) );
O2A1O1Ixp33_ASAP7_75t_L g930 ( .A1(n_921), .A2(n_815), .B(n_818), .C(n_813), .Y(n_930) );
OAI21xp5_ASAP7_75t_L g931 ( .A1(n_922), .A2(n_824), .B(n_907), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_918), .A2(n_919), .B1(n_923), .B2(n_921), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_926), .Y(n_933) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_924), .A2(n_900), .B1(n_813), .B2(n_894), .C(n_889), .Y(n_934) );
AOI21xp33_ASAP7_75t_L g935 ( .A1(n_925), .A2(n_868), .B(n_867), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_928), .Y(n_936) );
INVxp67_ASAP7_75t_L g937 ( .A(n_931), .Y(n_937) );
AOI221xp5_ASAP7_75t_L g938 ( .A1(n_934), .A2(n_909), .B1(n_910), .B2(n_911), .C(n_906), .Y(n_938) );
NOR3xp33_ASAP7_75t_L g939 ( .A(n_936), .B(n_930), .C(n_929), .Y(n_939) );
AOI211xp5_ASAP7_75t_L g940 ( .A1(n_937), .A2(n_935), .B(n_932), .C(n_933), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_940), .B(n_938), .Y(n_941) );
NAND3x1_ASAP7_75t_L g942 ( .A(n_939), .B(n_841), .C(n_806), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_941), .Y(n_943) );
XNOR2xp5_ASAP7_75t_L g944 ( .A(n_943), .B(n_942), .Y(n_944) );
OAI22xp5_ASAP7_75t_SL g945 ( .A1(n_944), .A2(n_833), .B1(n_798), .B2(n_774), .Y(n_945) );
AO21x2_ASAP7_75t_L g946 ( .A1(n_945), .A2(n_799), .B(n_797), .Y(n_946) );
AND2x4_ASAP7_75t_SL g947 ( .A(n_946), .B(n_770), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_947), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g949 ( .A1(n_948), .A2(n_917), .B1(n_857), .B2(n_895), .Y(n_949) );
endmodule