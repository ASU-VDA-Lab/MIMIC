module fake_jpeg_30394_n_527 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_7),
.B(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_22),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_94),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_85),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_8),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_87),
.Y(n_170)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_90),
.Y(n_163)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_17),
.B(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_8),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_6),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_102),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_105),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_26),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_52),
.B(n_41),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_133),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_67),
.B(n_35),
.Y(n_133)
);

NAND2x1_ASAP7_75t_SL g186 ( 
.A(n_136),
.B(n_35),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_94),
.B(n_38),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_42),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_69),
.B1(n_95),
.B2(n_64),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_157),
.B1(n_168),
.B2(n_51),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_39),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_54),
.B(n_29),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_46),
.B(n_25),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_154),
.A2(n_31),
.B(n_26),
.C(n_45),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_51),
.B1(n_49),
.B2(n_52),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_70),
.B(n_37),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_162),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_106),
.A2(n_51),
.B1(n_46),
.B2(n_48),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_159),
.A2(n_160),
.B1(n_43),
.B2(n_25),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_58),
.A2(n_37),
.B1(n_50),
.B2(n_48),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_57),
.B(n_38),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_24),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_59),
.A2(n_24),
.B1(n_50),
.B2(n_29),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_68),
.B(n_22),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_124),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_176),
.Y(n_225)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_187),
.Y(n_232)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_119),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_42),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_192),
.Y(n_233)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_191),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_122),
.B(n_34),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_118),
.B(n_34),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_194),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_126),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_204),
.Y(n_229)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_198),
.Y(n_239)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_124),
.A2(n_68),
.B1(n_71),
.B2(n_82),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_200),
.B1(n_210),
.B2(n_217),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_202),
.Y(n_247)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_205),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_110),
.B(n_33),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_207),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_33),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_131),
.B(n_41),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_209),
.Y(n_262)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_133),
.A2(n_45),
.B(n_90),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_157),
.Y(n_240)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_224),
.Y(n_261)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_135),
.A2(n_84),
.B1(n_80),
.B2(n_79),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_112),
.B1(n_150),
.B2(n_137),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_253)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

INVx5_ASAP7_75t_SL g221 ( 
.A(n_121),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_154),
.A2(n_71),
.B(n_45),
.C(n_74),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_164),
.B1(n_153),
.B2(n_149),
.Y(n_254)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_174),
.B(n_133),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_248),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_134),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_240),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_235),
.B1(n_249),
.B2(n_252),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_141),
.B1(n_164),
.B2(n_153),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_177),
.B(n_128),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_242),
.B(n_250),
.Y(n_280)
);

NAND2x1p5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_144),
.Y(n_243)
);

NOR2x1p5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_221),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_31),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_112),
.B1(n_150),
.B2(n_140),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_188),
.B(n_43),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_178),
.B(n_166),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_116),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_199),
.A2(n_77),
.B1(n_73),
.B2(n_76),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_183),
.A2(n_66),
.B1(n_151),
.B2(n_147),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_139),
.B1(n_201),
.B2(n_195),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_216),
.B1(n_173),
.B2(n_185),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_214),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_279),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_271),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_229),
.A2(n_186),
.B1(n_113),
.B2(n_170),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_278),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_125),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_268),
.C(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_230),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_277),
.B(n_286),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_232),
.B(n_202),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_189),
.B(n_179),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_258),
.B(n_263),
.Y(n_302)
);

INVx3_ASAP7_75t_SL g283 ( 
.A(n_228),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_283),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_198),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_289),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_231),
.A2(n_142),
.B(n_172),
.C(n_45),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_243),
.B(n_258),
.C(n_231),
.Y(n_301)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_291),
.B1(n_260),
.B2(n_200),
.Y(n_317)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_294),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_229),
.A2(n_140),
.B1(n_147),
.B2(n_151),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_297),
.B1(n_227),
.B2(n_261),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_229),
.A2(n_139),
.B1(n_134),
.B2(n_170),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_253),
.B1(n_237),
.B2(n_254),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_232),
.B(n_121),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_296),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_243),
.A2(n_224),
.B1(n_209),
.B2(n_210),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_248),
.A3(n_237),
.B1(n_231),
.B2(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_299),
.A2(n_304),
.B1(n_308),
.B2(n_319),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_301),
.B(n_285),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_286),
.B1(n_290),
.B2(n_272),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_240),
.Y(n_306)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_259),
.B(n_254),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_314),
.B(n_321),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_273),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_251),
.C(n_259),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_327),
.C(n_311),
.Y(n_337)
);

AOI22x1_ASAP7_75t_SL g314 ( 
.A1(n_278),
.A2(n_254),
.B1(n_252),
.B2(n_242),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_317),
.A2(n_324),
.B1(n_292),
.B2(n_283),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_270),
.A2(n_254),
.B1(n_233),
.B2(n_230),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_291),
.A2(n_262),
.B1(n_264),
.B2(n_256),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_270),
.A2(n_233),
.B1(n_260),
.B2(n_264),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_328),
.B1(n_281),
.B2(n_285),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_274),
.A2(n_277),
.B1(n_279),
.B2(n_293),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_257),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_265),
.A2(n_250),
.B1(n_262),
.B2(n_244),
.Y(n_328)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_354),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_282),
.B(n_268),
.C(n_296),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_331),
.A2(n_307),
.B(n_298),
.Y(n_374)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_300),
.Y(n_334)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_353),
.Y(n_362)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_343),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_339),
.A2(n_299),
.B1(n_308),
.B2(n_344),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_266),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_340),
.B(n_349),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_303),
.B1(n_297),
.B2(n_321),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_356),
.B1(n_322),
.B2(n_306),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_347),
.Y(n_364)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_316),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_316),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_284),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_352),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_325),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_327),
.C(n_300),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_280),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_303),
.A2(n_269),
.B1(n_295),
.B2(n_280),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_257),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_238),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_319),
.A2(n_269),
.B1(n_283),
.B2(n_288),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_246),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_361),
.B(n_374),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_365),
.C(n_368),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_351),
.B(n_313),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_363),
.B(n_383),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_320),
.C(n_302),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_355),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_307),
.C(n_320),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_307),
.B(n_328),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_369),
.A2(n_345),
.B(n_333),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_350),
.Y(n_370)
);

INVx13_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_377),
.B1(n_378),
.B2(n_384),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_331),
.B(n_306),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_341),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_329),
.A2(n_318),
.B1(n_323),
.B2(n_288),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_335),
.Y(n_379)
);

INVx13_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_389),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_381),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_336),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_386),
.B(n_379),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_356),
.A2(n_289),
.B1(n_275),
.B2(n_238),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_339),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_246),
.C(n_245),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_191),
.C(n_203),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_246),
.B1(n_228),
.B2(n_236),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_400),
.B1(n_410),
.B2(n_412),
.Y(n_427)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_397),
.B(n_401),
.Y(n_426)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_396),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_358),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_355),
.B1(n_346),
.B2(n_347),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_381),
.Y(n_402)
);

INVx11_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_341),
.Y(n_406)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_217),
.Y(n_436)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_361),
.B(n_343),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_408),
.A2(n_414),
.B1(n_375),
.B2(n_376),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_380),
.A2(n_338),
.B1(n_352),
.B2(n_330),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_411),
.A2(n_413),
.B1(n_129),
.B2(n_10),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_385),
.B(n_236),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_360),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_376),
.B(n_236),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_416),
.B(n_418),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_364),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_368),
.B(n_245),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_362),
.C(n_365),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_422),
.C(n_424),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_421),
.B(n_433),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_388),
.C(n_364),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_410),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_377),
.C(n_374),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_378),
.C(n_372),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_429),
.C(n_391),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_372),
.C(n_373),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_371),
.Y(n_433)
);

FAx1_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_384),
.CI(n_373),
.CON(n_434),
.SN(n_434)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_438),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_366),
.C(n_387),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_435),
.B(n_436),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_409),
.A2(n_182),
.B1(n_129),
.B2(n_116),
.Y(n_438)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_439),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_165),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_440),
.B(n_395),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_447),
.Y(n_466)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_455),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_397),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_437),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_454),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_450),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_452),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_426),
.A2(n_402),
.B(n_399),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_453),
.Y(n_465)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_395),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_459),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_396),
.C(n_411),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_458),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_426),
.A2(n_402),
.B(n_414),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_397),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_460),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_392),
.B1(n_406),
.B2(n_441),
.Y(n_461)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_446),
.A2(n_392),
.B(n_430),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_462),
.A2(n_416),
.B(n_460),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_445),
.A2(n_427),
.B1(n_393),
.B2(n_430),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_474),
.B1(n_475),
.B2(n_438),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_457),
.A2(n_406),
.B1(n_425),
.B2(n_424),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_477),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_455),
.A2(n_393),
.B1(n_440),
.B2(n_428),
.Y(n_474)
);

OAI321xp33_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_405),
.A3(n_404),
.B1(n_413),
.B2(n_415),
.C(n_434),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_458),
.A2(n_421),
.B1(n_429),
.B2(n_434),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_477),
.B(n_449),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_484),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_471),
.B(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_456),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_447),
.C(n_443),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_483),
.C(n_485),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_423),
.C(n_449),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_451),
.C(n_435),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_486),
.A2(n_467),
.B1(n_468),
.B2(n_464),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_408),
.C(n_415),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_487),
.B(n_488),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_404),
.C(n_165),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_463),
.A2(n_465),
.B(n_470),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_489),
.B(n_492),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_45),
.C(n_1),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_0),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_SL g492 ( 
.A(n_462),
.B(n_9),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_493),
.B(n_494),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_490),
.A2(n_474),
.B1(n_10),
.B2(n_11),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_482),
.A2(n_5),
.B1(n_14),
.B2(n_13),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_493),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_478),
.A2(n_15),
.B1(n_10),
.B2(n_5),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_498),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_488),
.Y(n_501)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_501),
.A2(n_491),
.B(n_1),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_15),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_0),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_506),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_483),
.C(n_485),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_496),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_504),
.B(n_0),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_499),
.C(n_501),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_500),
.A2(n_4),
.B(n_1),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_511),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_517),
.C(n_509),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_499),
.B(n_503),
.Y(n_516)
);

NAND2x1_ASAP7_75t_SL g518 ( 
.A(n_516),
.B(n_512),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_518),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_513),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_519),
.A2(n_520),
.B1(n_516),
.B2(n_515),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_522),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_0),
.B(n_2),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_524),
.A2(n_2),
.B(n_3),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_4),
.B(n_2),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_3),
.B(n_402),
.Y(n_527)
);


endmodule