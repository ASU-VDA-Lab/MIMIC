module fake_jpeg_8577_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_57),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_23),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_62),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_58),
.B1(n_23),
.B2(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_SL g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_31),
.B1(n_33),
.B2(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_39),
.C(n_38),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_76),
.C(n_78),
.Y(n_107)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_33),
.B1(n_17),
.B2(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_98),
.B1(n_54),
.B2(n_47),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_21),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_28),
.B1(n_27),
.B2(n_19),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_88),
.B1(n_95),
.B2(n_68),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_22),
.C(n_18),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_0),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_35),
.B1(n_30),
.B2(n_11),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_30),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_61),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_18),
.B1(n_35),
.B2(n_25),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_112),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_113),
.B1(n_100),
.B2(n_93),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_109),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_67),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_47),
.B1(n_18),
.B2(n_56),
.Y(n_113)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_78),
.B(n_1),
.Y(n_145)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_0),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_127),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_100),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_82),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_150),
.C(n_159),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_126),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_75),
.B1(n_83),
.B2(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_129),
.B1(n_120),
.B2(n_116),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_154),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_92),
.B1(n_101),
.B2(n_102),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_139),
.B1(n_114),
.B2(n_106),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_146),
.Y(n_179)
);

AND2x4_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_78),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_145),
.B(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_80),
.C(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_80),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_25),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_77),
.C(n_25),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_0),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_1),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_164),
.B1(n_142),
.B2(n_162),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_128),
.B1(n_116),
.B2(n_121),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_173),
.C(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_169),
.B(n_171),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_119),
.B1(n_115),
.B2(n_113),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_172),
.B1(n_143),
.B2(n_144),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_146),
.B1(n_149),
.B2(n_154),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_124),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_175),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_133),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_115),
.B(n_106),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_182),
.B1(n_193),
.B2(n_152),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_180),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_109),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_129),
.B1(n_121),
.B2(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_143),
.B1(n_161),
.B2(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_109),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_131),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_117),
.B1(n_109),
.B2(n_4),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_200),
.A2(n_206),
.B(n_210),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_162),
.B1(n_138),
.B2(n_160),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_212),
.B1(n_215),
.B2(n_221),
.Y(n_232)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_205),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_204),
.B(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_143),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_173),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_222),
.B1(n_193),
.B2(n_195),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_143),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_214),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_163),
.A2(n_170),
.B1(n_171),
.B2(n_194),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_167),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_133),
.B(n_148),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_218),
.B(n_176),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_214),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_143),
.B1(n_137),
.B2(n_158),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_159),
.B1(n_109),
.B2(n_117),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_190),
.C(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_224),
.C(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_190),
.C(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_230),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_234),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_237),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_206),
.B1(n_210),
.B2(n_197),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_180),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_191),
.B1(n_178),
.B2(n_181),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_238),
.B1(n_197),
.B2(n_205),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_174),
.B1(n_186),
.B2(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_186),
.C(n_183),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_248)
);

OAI322xp33_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_187),
.A3(n_168),
.B1(n_12),
.B2(n_13),
.C1(n_16),
.C2(n_8),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_213),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_168),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_117),
.C(n_3),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_204),
.C(n_222),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_258),
.C(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_204),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_202),
.B1(n_243),
.B2(n_11),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g256 ( 
.A(n_239),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_210),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_242),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_206),
.C(n_218),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_208),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_15),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_235),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_240),
.C(n_231),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_237),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_245),
.B1(n_249),
.B2(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_13),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_248),
.B1(n_250),
.B2(n_16),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_2),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_261),
.C(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_280),
.B(n_277),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_274),
.B(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_4),
.C(n_5),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_285),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

OAI311xp33_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_7),
.A3(n_286),
.B1(n_273),
.C1(n_281),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_7),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);


endmodule