module real_jpeg_33004_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_0),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_0),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_1),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_1),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_1),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_1),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_1),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_2),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_2),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_2),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_2),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_2),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_2),
.B(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_6),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_7),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_7),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_7),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_7),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_7),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_7),
.B(n_137),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_9),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_9),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_9),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_9),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_10),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_11),
.B(n_77),
.Y(n_76)
);

NAND2x1_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_12),
.Y(n_138)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_13),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_14),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_14),
.B(n_105),
.Y(n_104)
);

NAND2x1_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_127),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_14),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_14),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_15),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_15),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_15),
.B(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_191),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_188),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_164),
.B(n_167),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_21),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_21),
.A2(n_111),
.B1(n_165),
.B2(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.C(n_94),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_22),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.C(n_53),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_23),
.A2(n_24),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_25),
.B(n_32),
.C(n_37),
.Y(n_131)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_29),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_29),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_43),
.A2(n_44),
.B1(n_53),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_45),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_45),
.B(n_156),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_46),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_47),
.Y(n_269)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_47),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_48),
.A2(n_49),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_52),
.Y(n_271)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_53),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.C(n_64),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_54),
.B(n_64),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_59),
.B(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_60),
.B(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_94),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_79),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_76),
.C(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_90),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_81),
.A2(n_82),
.B1(n_90),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_84),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_85),
.B(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_90),
.Y(n_171)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_109),
.B2(n_110),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_96),
.Y(n_304)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_108),
.C(n_109),
.Y(n_163)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_104),
.Y(n_108)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_142),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_132),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_125),
.C(n_131),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.C(n_122),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_115),
.B(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_124),
.Y(n_235)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_126),
.B(n_129),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_152),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_156),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_156),
.A2(n_241),
.B1(n_243),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_190),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_184),
.C(n_186),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_184),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_172),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_174),
.A2(n_175),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_221),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_219),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_219),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.C(n_216),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.C(n_213),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.C(n_208),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_206),
.B(n_209),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_247),
.B(n_331),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_227),
.B(n_229),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.C(n_244),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_230),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_232),
.B(n_244),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_240),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_325),
.B(n_330),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_285),
.B(n_324),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_275),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_250),
.B(n_275),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_266),
.C(n_272),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_251),
.A2(n_252),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_259),
.B2(n_262),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_262),
.C(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_266),
.A2(n_272),
.B1(n_273),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

NAND2x1_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_270),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_280),
.C(n_327),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

AOI21x1_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_317),
.B(n_323),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_305),
.B(n_316),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_296),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_288),
.B(n_296),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_293),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx4f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_300),
.C(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_311),
.B(n_315),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_328),
.Y(n_330)
);


endmodule