module fake_jpeg_1471_n_395 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_23),
.B1(n_39),
.B2(n_38),
.Y(n_92)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_51),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_52),
.B(n_60),
.Y(n_123)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_1),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_1),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_64),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_2),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_68),
.Y(n_100)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_75),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_19),
.B(n_4),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_79),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_81),
.Y(n_109)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_80),
.A2(n_21),
.B(n_30),
.Y(n_132)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_23),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_84),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_88),
.B(n_116),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_97),
.B1(n_101),
.B2(n_129),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_41),
.B1(n_28),
.B2(n_19),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_21),
.C(n_39),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_46),
.C(n_77),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_41),
.B1(n_28),
.B2(n_38),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_28),
.B1(n_39),
.B2(n_25),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_112),
.B1(n_54),
.B2(n_63),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_110),
.B1(n_126),
.B2(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_48),
.A2(n_21),
.B1(n_38),
.B2(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_52),
.B(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_111),
.B(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_44),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_42),
.B(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_21),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_35),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_57),
.B(n_25),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_59),
.B(n_25),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_53),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_21),
.B1(n_27),
.B2(n_22),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_61),
.B(n_29),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_30),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_27),
.B1(n_29),
.B2(n_21),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_49),
.A2(n_27),
.B1(n_21),
.B2(n_32),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_5),
.Y(n_175)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_165),
.C(n_120),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_148),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_139),
.A2(n_146),
.B1(n_154),
.B2(n_162),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_30),
.B(n_71),
.C(n_47),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_147),
.B(n_161),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_75),
.B1(n_73),
.B2(n_50),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_141),
.A2(n_180),
.B1(n_102),
.B2(n_105),
.Y(n_204)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_126),
.B1(n_100),
.B2(n_103),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_144),
.A2(n_149),
.B1(n_169),
.B2(n_182),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_83),
.A2(n_79),
.B1(n_81),
.B2(n_32),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_30),
.B(n_32),
.C(n_24),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_88),
.B(n_83),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_150),
.A2(n_175),
.B(n_96),
.Y(n_211)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_5),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_163),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_87),
.A2(n_32),
.B1(n_24),
.B2(n_17),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

AO22x2_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_32),
.B1(n_24),
.B2(n_17),
.Y(n_156)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_167),
.C(n_5),
.Y(n_203)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_26),
.B(n_32),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_86),
.A2(n_32),
.B1(n_24),
.B2(n_17),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_94),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_98),
.B(n_24),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_168),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_24),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_87),
.A2(n_24),
.B1(n_17),
.B2(n_26),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_171),
.B1(n_182),
.B2(n_105),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_17),
.B1(n_26),
.B2(n_7),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_174),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_85),
.B(n_91),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_181),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_108),
.A2(n_17),
.B1(n_26),
.B2(n_7),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_112),
.A2(n_17),
.B1(n_6),
.B2(n_9),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_190),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_187),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_92),
.B(n_107),
.C(n_90),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_189),
.A2(n_156),
.B(n_172),
.C(n_181),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_107),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_201),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_211),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_158),
.A2(n_90),
.B1(n_82),
.B2(n_102),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_198),
.A2(n_204),
.B1(n_212),
.B2(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_102),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_135),
.B(n_93),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_214),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_139),
.B1(n_146),
.B2(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_96),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_220),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_118),
.C(n_92),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_161),
.C(n_159),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_138),
.A2(n_128),
.B1(n_95),
.B2(n_92),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_148),
.B(n_118),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_134),
.B(n_128),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g224 ( 
.A(n_167),
.B(n_95),
.C(n_9),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_151),
.Y(n_250)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_136),
.A2(n_6),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_246),
.C(n_259),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_190),
.B1(n_199),
.B2(n_212),
.Y(n_228)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_228),
.A2(n_251),
.B(n_260),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_141),
.B1(n_170),
.B2(n_154),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_238),
.A2(n_255),
.B1(n_191),
.B2(n_195),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_200),
.B1(n_204),
.B2(n_201),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_261),
.B1(n_219),
.B2(n_202),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_205),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_156),
.B1(n_140),
.B2(n_147),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_177),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_205),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_250),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_199),
.A2(n_156),
.B1(n_166),
.B2(n_160),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_163),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_256),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_198),
.B(n_225),
.C(n_197),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_156),
.B1(n_178),
.B2(n_143),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_193),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_211),
.A2(n_179),
.B(n_133),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_188),
.B(n_218),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_194),
.B(n_155),
.C(n_142),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_200),
.A2(n_168),
.B1(n_164),
.B2(n_11),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_264),
.A2(n_269),
.B(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_202),
.C(n_183),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_273),
.C(n_247),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_266),
.A2(n_232),
.B1(n_238),
.B2(n_255),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_206),
.B1(n_192),
.B2(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_267),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_213),
.Y(n_270)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_282),
.C(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_197),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_272),
.B(n_275),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_223),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_231),
.B(n_223),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_231),
.B(n_215),
.CI(n_186),
.CON(n_279),
.SN(n_279)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_293),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_242),
.A2(n_218),
.A3(n_187),
.B1(n_185),
.B2(n_208),
.C1(n_188),
.C2(n_195),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_281),
.B(n_283),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_208),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_191),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_228),
.B1(n_251),
.B2(n_232),
.Y(n_295)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_243),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_295),
.A2(n_302),
.B1(n_307),
.B2(n_310),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_291),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_297),
.B(n_315),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_227),
.C(n_258),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_235),
.C(n_233),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_235),
.C(n_233),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_242),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_286),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_259),
.C(n_257),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_305),
.C(n_312),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_248),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_280),
.A2(n_244),
.B1(n_256),
.B2(n_252),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_280),
.A2(n_244),
.B1(n_254),
.B2(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_248),
.C(n_237),
.Y(n_312)
);

OA21x2_ASAP7_75t_SL g314 ( 
.A1(n_263),
.A2(n_10),
.B(n_12),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_276),
.Y(n_327)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_14),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_318),
.C(n_277),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_10),
.C(n_13),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_310),
.B1(n_295),
.B2(n_280),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_269),
.B1(n_278),
.B2(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_271),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_327),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_332),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_264),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_330),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_305),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_301),
.B(n_279),
.CI(n_277),
.CON(n_334),
.SN(n_334)
);

AOI321xp33_ASAP7_75t_L g343 ( 
.A1(n_334),
.A2(n_299),
.A3(n_303),
.B1(n_313),
.B2(n_319),
.C(n_306),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_317),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_288),
.B(n_274),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_269),
.B(n_312),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_279),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_339),
.C(n_267),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_290),
.C(n_274),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_SL g341 ( 
.A(n_320),
.B(n_316),
.C(n_313),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_348),
.Y(n_362)
);

OAI31xp33_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_355),
.A3(n_336),
.B(n_344),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_344),
.A2(n_352),
.B(n_351),
.Y(n_367)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_331),
.Y(n_345)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

AOI321xp33_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_330),
.A3(n_338),
.B1(n_334),
.B2(n_321),
.C(n_329),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_336),
.B(n_349),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_351),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_280),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_353),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_278),
.C(n_280),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_332),
.C(n_335),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_354),
.A2(n_337),
.B1(n_333),
.B2(n_321),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g355 ( 
.A(n_322),
.B(n_269),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_328),
.B(n_326),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_349),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_357),
.A2(n_359),
.B1(n_363),
.B2(n_365),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_323),
.B1(n_339),
.B2(n_334),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_367),
.B(n_355),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_357),
.B(n_367),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_368),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.Y(n_370)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_356),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_350),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_376),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_372),
.A2(n_355),
.B1(n_368),
.B2(n_369),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_343),
.B(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_347),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_378),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_377),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_383),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_358),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_384),
.B(n_370),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_387),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_381),
.A2(n_374),
.B(n_376),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_358),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_379),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_386),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_389),
.A2(n_379),
.B(n_380),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_390),
.B(n_391),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_392),
.B(n_393),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_394),
.Y(n_395)
);


endmodule