module real_aes_5743_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_287;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_666;
wire n_320;
wire n_537;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_932;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_0), .A2(n_68), .B1(n_384), .B2(n_385), .Y(n_383) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_1), .Y(n_677) );
AND2x4_ASAP7_75t_L g687 ( .A(n_1), .B(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g695 ( .A(n_1), .B(n_240), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_2), .A2(n_37), .B1(n_711), .B2(n_712), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_3), .A2(n_72), .B1(n_469), .B2(n_472), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_4), .A2(n_101), .B1(n_446), .B2(n_450), .Y(n_609) );
INVx1_ASAP7_75t_L g519 ( .A(n_5), .Y(n_519) );
XOR2x2_ASAP7_75t_SL g503 ( .A(n_6), .B(n_504), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_7), .A2(n_151), .B1(n_444), .B2(n_447), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_8), .A2(n_109), .B1(n_701), .B2(n_702), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_9), .A2(n_86), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_10), .A2(n_225), .B1(n_435), .B2(n_436), .Y(n_575) );
INVx1_ASAP7_75t_L g935 ( .A(n_11), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_12), .A2(n_24), .B1(n_382), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_13), .A2(n_210), .B1(n_438), .B2(n_439), .Y(n_574) );
INVx1_ASAP7_75t_L g515 ( .A(n_14), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_15), .A2(n_246), .B1(n_446), .B2(n_447), .Y(n_897) );
INVx1_ASAP7_75t_L g649 ( .A(n_16), .Y(n_649) );
AO22x1_ASAP7_75t_L g584 ( .A1(n_17), .A2(n_137), .B1(n_452), .B2(n_453), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_18), .A2(n_135), .B1(n_474), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_19), .A2(n_46), .B1(n_376), .B2(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_20), .A2(n_172), .B1(n_328), .B2(n_335), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_21), .A2(n_184), .B1(n_352), .B2(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g640 ( .A(n_22), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_23), .A2(n_58), .B1(n_435), .B2(n_439), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_25), .A2(n_99), .B1(n_432), .B2(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g692 ( .A(n_26), .Y(n_692) );
INVx1_ASAP7_75t_L g526 ( .A(n_27), .Y(n_526) );
INVx1_ASAP7_75t_L g560 ( .A(n_28), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_29), .A2(n_103), .B1(n_707), .B2(n_709), .Y(n_724) );
INVx1_ASAP7_75t_L g908 ( .A(n_29), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_29), .A2(n_915), .B1(n_917), .B2(n_942), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_30), .A2(n_432), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g280 ( .A(n_31), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_31), .B(n_185), .Y(n_297) );
INVxp67_ASAP7_75t_L g316 ( .A(n_31), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_32), .A2(n_169), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_33), .A2(n_128), .B1(n_432), .B2(n_436), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_34), .A2(n_227), .B1(n_694), .B2(n_696), .Y(n_693) );
AO22x1_ASAP7_75t_L g582 ( .A1(n_35), .A2(n_131), .B1(n_446), .B2(n_450), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_36), .A2(n_64), .B1(n_432), .B2(n_433), .C(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_38), .B(n_265), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_39), .A2(n_234), .B1(n_306), .B2(n_308), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_40), .A2(n_238), .B1(n_335), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_41), .A2(n_219), .B1(n_354), .B2(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_42), .A2(n_114), .B1(n_391), .B2(n_392), .Y(n_390) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_43), .A2(n_593), .B(n_610), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_43), .B(n_594), .C(n_600), .D(n_607), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_44), .A2(n_67), .B1(n_260), .B2(n_283), .C(n_289), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_45), .A2(n_216), .B1(n_319), .B2(n_321), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_47), .A2(n_83), .B1(n_435), .B2(n_436), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_48), .A2(n_167), .B1(n_596), .B2(n_597), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_49), .A2(n_118), .B1(n_701), .B2(n_702), .Y(n_700) );
OAI22x1_ASAP7_75t_L g462 ( .A1(n_50), .A2(n_463), .B1(n_499), .B2(n_500), .Y(n_462) );
INVx1_ASAP7_75t_L g500 ( .A(n_50), .Y(n_500) );
NAND2xp33_ASAP7_75t_L g652 ( .A(n_51), .B(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_52), .A2(n_223), .B1(n_375), .B2(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_53), .A2(n_142), .B1(n_381), .B2(n_385), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_54), .B(n_433), .Y(n_573) );
INVx1_ASAP7_75t_L g556 ( .A(n_55), .Y(n_556) );
INVx2_ASAP7_75t_L g675 ( .A(n_56), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_57), .A2(n_205), .B1(n_485), .B2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g686 ( .A(n_59), .Y(n_686) );
AND2x4_ASAP7_75t_L g691 ( .A(n_59), .B(n_675), .Y(n_691) );
INVx1_ASAP7_75t_SL g708 ( .A(n_59), .Y(n_708) );
INVx1_ASAP7_75t_L g939 ( .A(n_60), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_61), .A2(n_62), .B1(n_340), .B2(n_342), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_63), .A2(n_191), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_65), .A2(n_102), .B1(n_438), .B2(n_903), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_66), .B(n_363), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_69), .A2(n_143), .B1(n_407), .B2(n_484), .Y(n_608) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_70), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_71), .A2(n_138), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_73), .A2(n_168), .B1(n_435), .B2(n_436), .Y(n_606) );
INVx1_ASAP7_75t_L g666 ( .A(n_74), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_75), .A2(n_181), .B1(n_438), .B2(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_76), .A2(n_88), .B1(n_489), .B2(n_491), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_77), .A2(n_144), .B1(n_711), .B2(n_712), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_78), .A2(n_163), .B1(n_438), .B2(n_439), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_79), .A2(n_87), .B1(n_373), .B2(n_558), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_80), .A2(n_230), .B1(n_447), .B2(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_81), .A2(n_182), .B1(n_637), .B2(n_638), .C(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_82), .A2(n_200), .B1(n_328), .B2(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g743 ( .A(n_84), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_85), .B(n_439), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_89), .A2(n_243), .B1(n_707), .B2(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g929 ( .A(n_90), .Y(n_929) );
AO22x1_ASAP7_75t_L g366 ( .A1(n_91), .A2(n_179), .B1(n_367), .B2(n_368), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_92), .A2(n_115), .B1(n_449), .B2(n_450), .Y(n_898) );
INVx1_ASAP7_75t_L g269 ( .A(n_93), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_93), .B(n_183), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_94), .A2(n_100), .B1(n_707), .B2(n_709), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_95), .A2(n_175), .B1(n_452), .B2(n_453), .Y(n_922) );
INVx1_ASAP7_75t_L g603 ( .A(n_96), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_97), .A2(n_201), .B1(n_345), .B2(n_382), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_98), .A2(n_212), .B1(n_370), .B2(n_372), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_104), .A2(n_226), .B1(n_483), .B2(n_485), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_105), .A2(n_176), .B1(n_340), .B2(n_342), .Y(n_510) );
INVx1_ASAP7_75t_L g578 ( .A(n_106), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_107), .B(n_420), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_108), .B(n_413), .Y(n_565) );
XOR2x2_ASAP7_75t_L g357 ( .A(n_109), .B(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_110), .A2(n_166), .B1(n_443), .B2(n_449), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_111), .A2(n_162), .B1(n_340), .B2(n_342), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_112), .A2(n_235), .B1(n_446), .B2(n_447), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_113), .A2(n_206), .B1(n_382), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_116), .A2(n_188), .B1(n_696), .B2(n_711), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_117), .A2(n_180), .B1(n_352), .B2(n_512), .Y(n_511) );
INVxp33_ASAP7_75t_SL g748 ( .A(n_119), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_120), .A2(n_149), .B1(n_684), .B2(n_704), .Y(n_703) );
XOR2xp5_ASAP7_75t_L g917 ( .A(n_121), .B(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_122), .A2(n_214), .B1(n_617), .B2(n_619), .Y(n_616) );
AO22x1_ASAP7_75t_L g583 ( .A1(n_123), .A2(n_237), .B1(n_443), .B2(n_449), .Y(n_583) );
INVx1_ASAP7_75t_L g524 ( .A(n_124), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_125), .A2(n_211), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_126), .A2(n_193), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_127), .A2(n_189), .B1(n_446), .B2(n_450), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_129), .A2(n_207), .B1(n_345), .B2(n_348), .Y(n_344) );
INVx1_ASAP7_75t_L g937 ( .A(n_130), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_132), .A2(n_361), .B(n_366), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_133), .A2(n_155), .B1(n_340), .B2(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g424 ( .A(n_134), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_136), .A2(n_147), .B1(n_386), .B2(n_405), .Y(n_404) );
AOI22x1_ASAP7_75t_L g612 ( .A1(n_139), .A2(n_613), .B1(n_614), .B2(n_641), .Y(n_612) );
INVx1_ASAP7_75t_L g641 ( .A(n_139), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_140), .A2(n_156), .B1(n_444), .B2(n_447), .Y(n_659) );
INVx1_ASAP7_75t_L g746 ( .A(n_141), .Y(n_746) );
CKINVDCx14_ASAP7_75t_R g427 ( .A(n_144), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_145), .A2(n_217), .B1(n_443), .B2(n_444), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_146), .A2(n_154), .B1(n_342), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_148), .A2(n_187), .B1(n_352), .B2(n_546), .Y(n_545) );
XNOR2x2_ASAP7_75t_L g570 ( .A(n_150), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_152), .B(n_368), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g374 ( .A1(n_153), .A2(n_178), .B1(n_375), .B2(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g933 ( .A(n_157), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_158), .A2(n_213), .B1(n_421), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_159), .A2(n_221), .B1(n_446), .B2(n_450), .Y(n_926) );
OA22x2_ASAP7_75t_L g263 ( .A1(n_160), .A2(n_185), .B1(n_264), .B2(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g304 ( .A(n_160), .Y(n_304) );
INVx1_ASAP7_75t_L g522 ( .A(n_161), .Y(n_522) );
AOI21xp5_ASAP7_75t_SL g931 ( .A1(n_164), .A2(n_432), .B(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_165), .A2(n_248), .B1(n_328), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_170), .A2(n_239), .B1(n_684), .B2(n_704), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_171), .A2(n_186), .B1(n_412), .B2(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g906 ( .A(n_173), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_174), .A2(n_228), .B1(n_494), .B2(n_496), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_177), .A2(n_215), .B1(n_380), .B2(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g282 ( .A(n_183), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_183), .B(n_301), .Y(n_300) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_185), .A2(n_202), .B(n_317), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_188), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_190), .A2(n_198), .B1(n_452), .B2(n_453), .Y(n_662) );
INVx1_ASAP7_75t_L g689 ( .A(n_192), .Y(n_689) );
INVx1_ASAP7_75t_L g563 ( .A(n_194), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_195), .A2(n_208), .B1(n_707), .B2(n_709), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_196), .A2(n_220), .B1(n_444), .B2(n_447), .Y(n_923) );
INVx1_ASAP7_75t_L g552 ( .A(n_197), .Y(n_552) );
INVx1_ASAP7_75t_SL g566 ( .A(n_199), .Y(n_566) );
INVx1_ASAP7_75t_L g271 ( .A(n_202), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_202), .B(n_231), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_203), .A2(n_245), .B1(n_443), .B2(n_449), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_204), .A2(n_229), .B1(n_452), .B2(n_453), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_209), .A2(n_242), .B1(n_474), .B2(n_475), .C(n_477), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_218), .A2(n_233), .B1(n_352), .B2(n_354), .Y(n_409) );
AOI21xp33_ASAP7_75t_SL g664 ( .A1(n_222), .A2(n_432), .B(n_665), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_224), .A2(n_260), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_231), .B(n_275), .Y(n_274) );
AOI21xp33_ASAP7_75t_L g904 ( .A1(n_232), .A2(n_435), .B(n_905), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_236), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g688 ( .A(n_240), .Y(n_688) );
INVxp33_ASAP7_75t_L g742 ( .A(n_241), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_244), .Y(n_290) );
INVx1_ASAP7_75t_L g478 ( .A(n_247), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_532), .B(n_669), .C(n_678), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_250), .A2(n_532), .B(n_670), .Y(n_669) );
XOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_396), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_357), .B1(n_394), .B2(n_395), .Y(n_252) );
INVx2_ASAP7_75t_L g395 ( .A(n_253), .Y(n_395) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
XNOR2x1_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_326), .Y(n_257) );
NAND3xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_305), .C(n_318), .Y(n_258) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g376 ( .A(n_261), .Y(n_376) );
INVx1_ASAP7_75t_L g518 ( .A(n_261), .Y(n_518) );
BUFx3_ASAP7_75t_L g637 ( .A(n_261), .Y(n_637) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_272), .Y(n_261) );
AND2x4_ASAP7_75t_L g320 ( .A(n_262), .B(n_287), .Y(n_320) );
AND2x2_ASAP7_75t_L g432 ( .A(n_262), .B(n_287), .Y(n_432) );
AND2x4_ASAP7_75t_L g435 ( .A(n_262), .B(n_272), .Y(n_435) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
AND2x2_ASAP7_75t_L g286 ( .A(n_263), .B(n_267), .Y(n_286) );
AND2x2_ASAP7_75t_L g314 ( .A(n_263), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g331 ( .A(n_263), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_264), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp33_ASAP7_75t_L g268 ( .A(n_265), .B(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
INVx1_ASAP7_75t_L g317 ( .A(n_265), .Y(n_317) );
AND2x4_ASAP7_75t_L g330 ( .A(n_266), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_269), .B(n_304), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_271), .A2(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g307 ( .A(n_272), .B(n_286), .Y(n_307) );
AND2x4_ASAP7_75t_L g341 ( .A(n_272), .B(n_330), .Y(n_341) );
AND2x4_ASAP7_75t_L g438 ( .A(n_272), .B(n_286), .Y(n_438) );
AND2x4_ASAP7_75t_L g452 ( .A(n_272), .B(n_330), .Y(n_452) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
INVx2_ASAP7_75t_L g288 ( .A(n_273), .Y(n_288) );
AND2x2_ASAP7_75t_L g311 ( .A(n_273), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g332 ( .A(n_273), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g338 ( .A(n_273), .B(n_334), .Y(n_338) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_276), .B(n_300), .C(n_302), .Y(n_299) );
AND2x4_ASAP7_75t_L g287 ( .A(n_277), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g334 ( .A(n_278), .Y(n_334) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g528 ( .A(n_284), .Y(n_528) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g365 ( .A(n_285), .Y(n_365) );
BUFx3_ASAP7_75t_L g420 ( .A(n_285), .Y(n_420) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x4_ASAP7_75t_L g346 ( .A(n_286), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_286), .B(n_332), .Y(n_353) );
AND2x2_ASAP7_75t_L g433 ( .A(n_286), .B(n_287), .Y(n_433) );
AND2x4_ASAP7_75t_L g446 ( .A(n_286), .B(n_332), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_286), .B(n_337), .Y(n_447) );
AND2x2_ASAP7_75t_L g495 ( .A(n_286), .B(n_332), .Y(n_495) );
AND2x4_ASAP7_75t_L g323 ( .A(n_287), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g343 ( .A(n_287), .B(n_330), .Y(n_343) );
AND2x4_ASAP7_75t_L g436 ( .A(n_287), .B(n_324), .Y(n_436) );
AND2x4_ASAP7_75t_L g453 ( .A(n_287), .B(n_330), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_291), .B(n_666), .Y(n_665) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_SL g368 ( .A(n_292), .Y(n_368) );
INVx1_ASAP7_75t_L g554 ( .A(n_292), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_292), .B(n_933), .Y(n_932) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g423 ( .A(n_293), .Y(n_423) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_296), .B(n_299), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_295), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_296), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_301), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g324 ( .A(n_302), .B(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g377 ( .A(n_306), .Y(n_377) );
INVx2_ASAP7_75t_L g520 ( .A(n_306), .Y(n_520) );
BUFx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_307), .Y(n_412) );
INVx2_ASAP7_75t_L g634 ( .A(n_307), .Y(n_634) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g367 ( .A(n_309), .Y(n_367) );
INVx4_ASAP7_75t_L g413 ( .A(n_309), .Y(n_413) );
INVx3_ASAP7_75t_L g474 ( .A(n_309), .Y(n_474) );
INVx5_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_310), .Y(n_530) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
AND2x4_ASAP7_75t_L g439 ( .A(n_311), .B(n_314), .Y(n_439) );
AND2x2_ASAP7_75t_L g903 ( .A(n_311), .B(n_314), .Y(n_903) );
INVx2_ASAP7_75t_L g523 ( .A(n_319), .Y(n_523) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_320), .Y(n_371) );
INVx2_ASAP7_75t_L g418 ( .A(n_320), .Y(n_418) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_320), .Y(n_471) );
INVx2_ASAP7_75t_L g559 ( .A(n_320), .Y(n_559) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g472 ( .A(n_322), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_322), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_521) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_323), .Y(n_373) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_323), .Y(n_415) );
AND2x4_ASAP7_75t_L g350 ( .A(n_324), .B(n_337), .Y(n_350) );
AND2x4_ASAP7_75t_L g356 ( .A(n_324), .B(n_332), .Y(n_356) );
AND2x4_ASAP7_75t_L g444 ( .A(n_324), .B(n_337), .Y(n_444) );
AND2x4_ASAP7_75t_L g450 ( .A(n_324), .B(n_332), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g326 ( .A(n_327), .B(n_339), .C(n_344), .D(n_351), .Y(n_326) );
BUFx2_ASAP7_75t_SL g391 ( .A(n_328), .Y(n_391) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx12f_ASAP7_75t_L g484 ( .A(n_329), .Y(n_484) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_329), .Y(n_542) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AND2x4_ASAP7_75t_L g336 ( .A(n_330), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g443 ( .A(n_330), .B(n_347), .Y(n_443) );
AND2x4_ASAP7_75t_L g449 ( .A(n_330), .B(n_332), .Y(n_449) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_336), .Y(n_407) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_336), .Y(n_487) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_336), .Y(n_507) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g347 ( .A(n_338), .Y(n_347) );
BUFx12f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g490 ( .A(n_341), .Y(n_490) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_341), .Y(n_544) );
BUFx2_ASAP7_75t_SL g491 ( .A(n_342), .Y(n_491) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx5_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
BUFx3_ASAP7_75t_L g597 ( .A(n_343), .Y(n_597) );
INVx1_ASAP7_75t_L g622 ( .A(n_343), .Y(n_622) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_346), .Y(n_509) );
BUFx3_ASAP7_75t_L g629 ( .A(n_346), .Y(n_629) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx5_ASAP7_75t_L g405 ( .A(n_349), .Y(n_405) );
INVx3_ASAP7_75t_L g599 ( .A(n_349), .Y(n_599) );
INVx6_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
BUFx3_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx8_ASAP7_75t_L g627 ( .A(n_353), .Y(n_627) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
INVx1_ASAP7_75t_L g497 ( .A(n_355), .Y(n_497) );
INVx4_ASAP7_75t_L g512 ( .A(n_355), .Y(n_512) );
INVx4_ASAP7_75t_L g546 ( .A(n_355), .Y(n_546) );
INVx8_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
NOR2x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_378), .Y(n_358) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_369), .C(n_374), .Y(n_359) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g476 ( .A(n_364), .Y(n_476) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx4_ASAP7_75t_L g561 ( .A(n_373), .Y(n_561) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND4xp25_ASAP7_75t_SL g378 ( .A(n_379), .B(n_383), .C(n_387), .D(n_390), .Y(n_378) );
BUFx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
XNOR2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_460), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_425), .B1(n_457), .B2(n_459), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g458 ( .A(n_399), .Y(n_458) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XOR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_424), .Y(n_401) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_410), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .C(n_408), .D(n_409), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .C(n_416), .D(n_419), .Y(n_410) );
BUFx3_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
INVx3_ASAP7_75t_L g564 ( .A(n_412), .Y(n_564) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g638 ( .A(n_420), .Y(n_638) );
INVx4_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_422), .B(n_578), .Y(n_577) );
INVx4_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g479 ( .A(n_423), .Y(n_479) );
INVx2_ASAP7_75t_L g459 ( .A(n_425), .Y(n_459) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI21x1_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_454), .Y(n_426) );
NAND3xp33_ASAP7_75t_SL g454 ( .A(n_427), .B(n_455), .C(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_441), .Y(n_429) );
INVx1_ASAP7_75t_L g456 ( .A(n_430), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .C(n_437), .D(n_440), .Y(n_430) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_433), .Y(n_653) );
INVx2_ASAP7_75t_L g930 ( .A(n_433), .Y(n_930) );
INVx2_ASAP7_75t_L g936 ( .A(n_435), .Y(n_936) );
INVx2_ASAP7_75t_L g656 ( .A(n_436), .Y(n_656) );
INVx1_ASAP7_75t_L g940 ( .A(n_438), .Y(n_940) );
INVxp67_ASAP7_75t_L g455 ( .A(n_441), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .C(n_448), .D(n_451), .Y(n_441) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_501), .B1(n_502), .B2(n_531), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g531 ( .A(n_462), .Y(n_531) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_480), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_464), .B(n_480), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_479), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_479), .B(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_479), .B(n_906), .Y(n_905) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_488), .Y(n_481) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx12f_ASAP7_75t_L g624 ( .A(n_484), .Y(n_624) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g596 ( .A(n_490), .Y(n_596) );
INVx2_ASAP7_75t_L g618 ( .A(n_490), .Y(n_618) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .Y(n_492) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
AND4x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .C(n_510), .D(n_511), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_521), .C(n_525), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_519), .B2(n_520), .Y(n_514) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_587), .B1(n_667), .B2(n_668), .Y(n_532) );
INVx1_ASAP7_75t_L g667 ( .A(n_533), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_567), .B1(n_585), .B2(n_586), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g585 ( .A(n_537), .Y(n_585) );
XOR2x1_ASAP7_75t_L g537 ( .A(n_538), .B(n_566), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .Y(n_538) );
AND4x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .C(n_543), .D(n_545), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_555), .C(n_562), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_560), .B2(n_561), .Y(n_555) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_565), .Y(n_562) );
INVx2_ASAP7_75t_L g586 ( .A(n_567), .Y(n_586) );
BUFx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_579), .Y(n_571) );
AND4x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .C(n_575), .D(n_576), .Y(n_572) );
NOR4xp25_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .C(n_583), .D(n_584), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g668 ( .A(n_587), .Y(n_668) );
XOR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_646), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_611), .B1(n_642), .B2(n_644), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g645 ( .A(n_590), .Y(n_645) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND3x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_600), .C(n_607), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g643 ( .A(n_612), .Y(n_643) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND4xp75_ASAP7_75t_L g614 ( .A(n_615), .B(n_625), .C(n_630), .D(n_636), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_623), .Y(n_615) );
BUFx4f_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx3_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
XNOR2x1_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_658), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .C(n_657), .Y(n_651) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_656), .A2(n_935), .B1(n_936), .B2(n_937), .Y(n_934) );
NAND4xp25_ASAP7_75t_SL g658 ( .A(n_659), .B(n_660), .C(n_661), .D(n_664), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
BUFx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .C(n_677), .Y(n_672) );
AND2x2_ASAP7_75t_L g911 ( .A(n_673), .B(n_912), .Y(n_911) );
AND2x2_ASAP7_75t_L g916 ( .A(n_673), .B(n_913), .Y(n_916) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OA21x2_ASAP7_75t_L g943 ( .A1(n_674), .A2(n_708), .B(n_944), .Y(n_943) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g685 ( .A(n_675), .B(n_686), .Y(n_685) );
AND3x4_ASAP7_75t_L g707 ( .A(n_675), .B(n_687), .C(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_676), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_677), .Y(n_913) );
OAI221xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_889), .B1(n_890), .B2(n_909), .C(n_914), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_697), .B(n_776), .C(n_885), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI221xp5_ASAP7_75t_SL g806 ( .A1(n_681), .A2(n_805), .B1(n_807), .B2(n_808), .C(n_809), .Y(n_806) );
INVx1_ASAP7_75t_L g849 ( .A(n_681), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_681), .B(n_781), .Y(n_861) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_682), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_689), .B1(n_690), .B2(n_692), .C(n_693), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_683), .A2(n_690), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
AND2x4_ASAP7_75t_L g694 ( .A(n_685), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g701 ( .A(n_685), .B(n_695), .Y(n_701) );
AND2x2_ASAP7_75t_L g711 ( .A(n_685), .B(n_695), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_687), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g704 ( .A(n_687), .B(n_691), .Y(n_704) );
AND2x4_ASAP7_75t_L g709 ( .A(n_687), .B(n_691), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_687), .Y(n_944) );
BUFx2_ASAP7_75t_L g889 ( .A(n_690), .Y(n_889) );
AND2x4_ASAP7_75t_L g696 ( .A(n_691), .B(n_695), .Y(n_696) );
AND2x2_ASAP7_75t_L g702 ( .A(n_691), .B(n_695), .Y(n_702) );
AND2x2_ASAP7_75t_L g712 ( .A(n_691), .B(n_695), .Y(n_712) );
INVx3_ASAP7_75t_L g745 ( .A(n_694), .Y(n_745) );
INVx2_ASAP7_75t_L g747 ( .A(n_696), .Y(n_747) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_713), .B(n_726), .C(n_766), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_698), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g769 ( .A(n_698), .Y(n_769) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_705), .Y(n_698) );
INVx1_ASAP7_75t_L g782 ( .A(n_699), .Y(n_782) );
INVx1_ASAP7_75t_L g794 ( .A(n_699), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
AND2x2_ASAP7_75t_L g739 ( .A(n_705), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g775 ( .A(n_705), .B(n_740), .Y(n_775) );
INVx2_ASAP7_75t_L g801 ( .A(n_705), .Y(n_801) );
OR2x2_ASAP7_75t_L g809 ( .A(n_705), .B(n_794), .Y(n_809) );
AND2x2_ASAP7_75t_L g818 ( .A(n_705), .B(n_794), .Y(n_818) );
OR2x2_ASAP7_75t_L g822 ( .A(n_705), .B(n_754), .Y(n_822) );
AND2x2_ASAP7_75t_L g848 ( .A(n_705), .B(n_793), .Y(n_848) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_705), .Y(n_856) );
AND2x2_ASAP7_75t_L g860 ( .A(n_705), .B(n_754), .Y(n_860) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .Y(n_705) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI31xp33_ASAP7_75t_L g766 ( .A1(n_714), .A2(n_735), .A3(n_767), .B(n_773), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_714), .A2(n_771), .B1(n_775), .B2(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_719), .Y(n_714) );
AND2x2_ASAP7_75t_L g796 ( .A(n_715), .B(n_728), .Y(n_796) );
AND2x2_ASAP7_75t_L g819 ( .A(n_715), .B(n_772), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_715), .B(n_723), .Y(n_826) );
AND2x2_ASAP7_75t_L g881 ( .A(n_715), .B(n_734), .Y(n_881) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g727 ( .A(n_716), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g737 ( .A(n_716), .Y(n_737) );
AND2x2_ASAP7_75t_L g771 ( .A(n_716), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_716), .B(n_723), .Y(n_805) );
OR2x2_ASAP7_75t_L g811 ( .A(n_716), .B(n_733), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_716), .A2(n_817), .B1(n_819), .B2(n_820), .C(n_823), .Y(n_816) );
OR2x2_ASAP7_75t_L g824 ( .A(n_716), .B(n_758), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_716), .B(n_813), .Y(n_853) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_719), .B(n_785), .Y(n_807) );
AND2x2_ASAP7_75t_L g846 ( .A(n_719), .B(n_736), .Y(n_846) );
INVx1_ASAP7_75t_L g858 ( .A(n_719), .Y(n_858) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .Y(n_719) );
OR2x2_ASAP7_75t_L g733 ( .A(n_720), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g738 ( .A(n_720), .B(n_734), .Y(n_738) );
OR2x2_ASAP7_75t_L g758 ( .A(n_720), .B(n_723), .Y(n_758) );
INVx1_ASAP7_75t_L g772 ( .A(n_720), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_720), .A2(n_779), .B1(n_789), .B2(n_792), .C(n_795), .Y(n_778) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g734 ( .A(n_723), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_723), .A2(n_855), .B1(n_857), .B2(n_859), .Y(n_854) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_735), .B(n_739), .C(n_749), .Y(n_726) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .Y(n_728) );
AND2x2_ASAP7_75t_L g751 ( .A(n_729), .B(n_740), .Y(n_751) );
AND2x2_ASAP7_75t_L g770 ( .A(n_729), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g774 ( .A(n_729), .Y(n_774) );
INVx2_ASAP7_75t_L g785 ( .A(n_729), .Y(n_785) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_729), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g803 ( .A(n_729), .B(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g813 ( .A(n_729), .B(n_738), .Y(n_813) );
INVx2_ASAP7_75t_L g833 ( .A(n_729), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_729), .B(n_782), .Y(n_882) );
INVx4_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g765 ( .A(n_730), .B(n_736), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_730), .B(n_754), .Y(n_791) );
AND2x2_ASAP7_75t_L g829 ( .A(n_730), .B(n_740), .Y(n_829) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx3_ASAP7_75t_SL g842 ( .A(n_733), .Y(n_842) );
NAND2xp67_ASAP7_75t_L g878 ( .A(n_735), .B(n_785), .Y(n_878) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
AND2x4_ASAP7_75t_L g756 ( .A(n_736), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g764 ( .A(n_738), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_738), .B(n_828), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_738), .A2(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_739), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g808 ( .A(n_739), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_739), .A2(n_804), .B1(n_820), .B2(n_877), .C(n_879), .Y(n_876) );
INVx2_ASAP7_75t_L g754 ( .A(n_740), .Y(n_754) );
INVx1_ASAP7_75t_L g761 ( .A(n_740), .Y(n_761) );
AND2x2_ASAP7_75t_L g817 ( .A(n_740), .B(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B(n_755), .C(n_759), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_751), .B(n_781), .Y(n_825) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g815 ( .A(n_754), .B(n_782), .Y(n_815) );
INVx2_ASAP7_75t_L g831 ( .A(n_754), .Y(n_831) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_756), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_758), .B(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_760), .B(n_792), .Y(n_872) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_761), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_763), .B(n_808), .Y(n_884) );
OR2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g841 ( .A(n_765), .Y(n_841) );
INVxp33_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
O2A1O1Ixp33_ASAP7_75t_L g883 ( .A1(n_770), .A2(n_821), .B(n_846), .C(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_774), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g788 ( .A(n_775), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_775), .A2(n_824), .B1(n_825), .B2(n_826), .C(n_827), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_775), .A2(n_803), .B1(n_809), .B2(n_880), .Y(n_879) );
NAND5xp2_ASAP7_75t_L g776 ( .A(n_777), .B(n_850), .C(n_870), .D(n_876), .E(n_883), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_797), .B(n_835), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .B1(n_786), .B2(n_788), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g820 ( .A(n_781), .B(n_821), .Y(n_820) );
AOI21xp33_ASAP7_75t_L g885 ( .A1(n_781), .A2(n_886), .B(n_888), .Y(n_885) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
BUFx3_ASAP7_75t_L g867 ( .A(n_782), .Y(n_867) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_786), .B(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_786), .B(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_787), .B(n_845), .Y(n_844) );
OAI21xp33_ASAP7_75t_SL g851 ( .A1(n_787), .A2(n_852), .B(n_853), .Y(n_851) );
AND2x2_ASAP7_75t_L g866 ( .A(n_788), .B(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g888 ( .A(n_796), .Y(n_888) );
NAND3xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_816), .C(n_830), .Y(n_797) );
AOI211xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .B(n_806), .C(n_810), .Y(n_798) );
CKINVDCx14_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
CKINVDCx14_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
AND2x2_ASAP7_75t_L g828 ( .A(n_801), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AOI21xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B(n_814), .Y(n_810) );
INVx1_ASAP7_75t_L g869 ( .A(n_811), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g862 ( .A1(n_812), .A2(n_863), .B(n_865), .C(n_868), .Y(n_862) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_817), .B(n_869), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_818), .A2(n_851), .B1(n_854), .B2(n_861), .C(n_862), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_819), .Y(n_852) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g834 ( .A(n_824), .Y(n_834) );
INVx1_ASAP7_75t_L g864 ( .A(n_826), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
INVx2_ASAP7_75t_L g843 ( .A(n_831), .Y(n_843) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g837 ( .A(n_833), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_838), .B(n_847), .C(n_849), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_837), .B(n_846), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_843), .B(n_844), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_843), .B(n_878), .Y(n_887) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
OAI211xp5_ASAP7_75t_L g870 ( .A1(n_860), .A2(n_871), .B(n_873), .C(n_875), .Y(n_870) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVxp67_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVxp33_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
XOR2x2_ASAP7_75t_L g893 ( .A(n_894), .B(n_908), .Y(n_893) );
NOR2xp67_ASAP7_75t_L g894 ( .A(n_895), .B(n_900), .Y(n_894) );
NAND4xp25_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .C(n_898), .D(n_899), .Y(n_895) );
NAND4xp25_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .C(n_904), .D(n_907), .Y(n_900) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVxp33_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_927), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_924), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .Y(n_924) );
NOR3xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_934), .C(n_938), .Y(n_927) );
OAI21xp33_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B(n_931), .Y(n_928) );
OAI21xp5_ASAP7_75t_SL g938 ( .A1(n_939), .A2(n_940), .B(n_941), .Y(n_938) );
BUFx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
endmodule