module fake_netlist_1_296_n_18 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_18);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
NAND2xp5_ASAP7_75t_L g8 ( .A(n_7), .B(n_4), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_5), .B(n_1), .Y(n_9) );
NOR2xp33_ASAP7_75t_L g10 ( .A(n_3), .B(n_7), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
AOI22xp5_ASAP7_75t_L g12 ( .A1(n_2), .A2(n_6), .B1(n_3), .B2(n_0), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
OAI22xp5_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_13), .B(n_8), .Y(n_15) );
NOR3xp33_ASAP7_75t_L g16 ( .A(n_15), .B(n_14), .C(n_9), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_16), .B(n_10), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_10), .B1(n_4), .B2(n_6), .Y(n_18) );
endmodule