module fake_aes_189_n_29 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVxp67_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
OAI22xp5_ASAP7_75t_SL g15 ( .A1(n_6), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_1), .B(n_9), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_0), .B(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_18), .B(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_21), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_25), .B(n_15), .C(n_14), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_20), .Y(n_27) );
AOI222xp33_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_5), .B1(n_7), .B2(n_8), .C1(n_10), .C2(n_13), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
endmodule