module fake_jpeg_24205_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_45),
.B1(n_21),
.B2(n_19),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_28),
.B1(n_32),
.B2(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_16),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_57),
.B(n_40),
.C(n_38),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_36),
.B1(n_37),
.B2(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_18),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_60),
.B(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_63),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_80),
.Y(n_95)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_24),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_87),
.B1(n_18),
.B2(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_84),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_19),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_36),
.B1(n_29),
.B2(n_20),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_40),
.A3(n_38),
.B1(n_49),
.B2(n_56),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_33),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_102),
.B1(n_103),
.B2(n_76),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_64),
.B1(n_61),
.B2(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_45),
.B1(n_40),
.B2(n_38),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_40),
.B(n_22),
.C(n_27),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_27),
.B(n_22),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_78),
.A3(n_59),
.B1(n_77),
.B2(n_80),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_42),
.B1(n_18),
.B2(n_46),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_18),
.B1(n_56),
.B2(n_31),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_18),
.B1(n_56),
.B2(n_17),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_17),
.B1(n_33),
.B2(n_26),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_118),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_112),
.B1(n_58),
.B2(n_107),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_86),
.B(n_74),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_130),
.B(n_133),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_67),
.C(n_84),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_132),
.C(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_135),
.Y(n_144)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_131),
.B1(n_134),
.B2(n_85),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_83),
.B1(n_81),
.B2(n_67),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_39),
.C(n_34),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_33),
.B(n_63),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_0),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_139),
.B(n_94),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_39),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_140),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_0),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_149),
.B(n_161),
.Y(n_194)
);

AO22x2_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_7),
.B(n_8),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_98),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_104),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_160),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_139),
.B1(n_118),
.B2(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_156),
.A2(n_173),
.B1(n_174),
.B2(n_9),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_114),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_135),
.C(n_129),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_88),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_115),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_0),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_113),
.B(n_25),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_108),
.C(n_93),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_170),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_69),
.Y(n_176)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_7),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_116),
.A2(n_85),
.B1(n_63),
.B2(n_88),
.Y(n_173)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_69),
.Y(n_177)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_183),
.B(n_191),
.Y(n_205)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_197),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_93),
.B1(n_113),
.B2(n_92),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_195),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_92),
.B1(n_26),
.B2(n_39),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_1),
.B(n_2),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_184),
.B(n_187),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_174),
.A2(n_34),
.B1(n_26),
.B2(n_3),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_144),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_34),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_161),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_203),
.B1(n_185),
.B2(n_188),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_158),
.C(n_150),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_217),
.C(n_221),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_176),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_186),
.B1(n_197),
.B2(n_189),
.Y(n_236)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_152),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_219),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_168),
.C(n_165),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_149),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_166),
.C(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_197),
.B(n_199),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_242),
.B(n_162),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_202),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_214),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_175),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_10),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_238),
.B1(n_212),
.B2(n_210),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_191),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_240),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_195),
.B1(n_164),
.B2(n_182),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_202),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_191),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.C(n_205),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_178),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_253),
.B1(n_249),
.B2(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_248),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_183),
.B(n_207),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_250),
.B1(n_256),
.B2(n_227),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_218),
.B1(n_213),
.B2(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_226),
.B1(n_245),
.B2(n_250),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_220),
.B(n_216),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_224),
.B1(n_196),
.B2(n_181),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_223),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_257),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_171),
.B(n_200),
.C(n_204),
.D(n_222),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_10),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_261),
.B(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_263),
.B1(n_269),
.B2(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_270),
.Y(n_272)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_231),
.B1(n_243),
.B2(n_254),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_252),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_229),
.C(n_12),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_280),
.B(n_14),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_275),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_11),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_11),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_265),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_13),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_267),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_276),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_275),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_11),
.B(n_12),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_284),
.B(n_286),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_14),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_13),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_14),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_15),
.C(n_285),
.Y(n_292)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_273),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_288),
.B(n_15),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_298),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_296),
.Y(n_301)
);


endmodule