module fake_jpeg_15568_n_396 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_47),
.B(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_62),
.Y(n_104)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_31),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_64),
.Y(n_107)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_16),
.B(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_28),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_68),
.B(n_89),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_22),
.B1(n_26),
.B2(n_38),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_70),
.A2(n_75),
.B1(n_77),
.B2(n_97),
.Y(n_140)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_34),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_22),
.B1(n_26),
.B2(n_38),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_115),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_37),
.B1(n_23),
.B2(n_24),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_88),
.B(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_37),
.B1(n_31),
.B2(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_17),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_19),
.B1(n_32),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_108),
.B1(n_59),
.B2(n_48),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_45),
.A2(n_25),
.B1(n_36),
.B2(n_35),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_105),
.B1(n_69),
.B2(n_81),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_37),
.B1(n_33),
.B2(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_55),
.A2(n_28),
.B1(n_33),
.B2(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_62),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_27),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_76),
.Y(n_134)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_125),
.Y(n_173)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_34),
.Y(n_121)
);

XNOR2x1_ASAP7_75t_SL g187 ( 
.A(n_121),
.B(n_83),
.Y(n_187)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_33),
.B1(n_24),
.B2(n_19),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_138),
.B1(n_27),
.B2(n_21),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_134),
.Y(n_176)
);

AO22x1_ASAP7_75t_SL g130 ( 
.A1(n_77),
.A2(n_59),
.B1(n_48),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_101),
.B1(n_109),
.B2(n_93),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_79),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_137),
.Y(n_193)
);

INVx6_ASAP7_75t_SL g137 ( 
.A(n_82),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_30),
.B1(n_21),
.B2(n_2),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_151),
.Y(n_204)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_63),
.C(n_39),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_155),
.C(n_4),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_14),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_29),
.Y(n_147)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_10),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_10),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_150),
.B(n_162),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_165),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_69),
.B(n_46),
.C(n_30),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_62),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_158),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_8),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_157),
.A2(n_159),
.B(n_13),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_40),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_70),
.B(n_7),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_80),
.B(n_9),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_84),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_9),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_166),
.B(n_167),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_91),
.B(n_5),
.Y(n_167)
);

INVx6_ASAP7_75t_SL g168 ( 
.A(n_79),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_171),
.Y(n_215)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_83),
.B(n_27),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_172),
.B(n_184),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_175),
.B1(n_211),
.B2(n_213),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_109),
.B1(n_117),
.B2(n_93),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_216),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_180),
.A2(n_161),
.B1(n_137),
.B2(n_143),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_126),
.A2(n_21),
.B(n_13),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_183),
.A2(n_208),
.B(n_198),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_123),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_149),
.A2(n_113),
.B1(n_87),
.B2(n_117),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_185),
.A2(n_186),
.B1(n_207),
.B2(n_212),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_126),
.A2(n_140),
.B1(n_130),
.B2(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_187),
.B(n_139),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_200),
.B1(n_168),
.B2(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_113),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_199),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_132),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_195),
.B(n_218),
.Y(n_235)
);

AO21x2_ASAP7_75t_L g196 ( 
.A1(n_130),
.A2(n_0),
.B(n_1),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_165),
.B(n_132),
.Y(n_239)
);

NAND2x1_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_0),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_198),
.A2(n_209),
.B(n_213),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_0),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_205),
.C(n_152),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_3),
.C(n_4),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_3),
.B1(n_10),
.B2(n_12),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_142),
.A2(n_159),
.B1(n_148),
.B2(n_153),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_131),
.A2(n_12),
.B1(n_13),
.B2(n_1),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_12),
.B1(n_13),
.B2(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_122),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_128),
.B(n_1),
.CI(n_121),
.CON(n_218),
.SN(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_258),
.B1(n_261),
.B2(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_223),
.B(n_225),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_218),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_125),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_259),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_244),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_120),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_256),
.C(n_205),
.Y(n_262)
);

CKINVDCx6p67_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_239),
.A2(n_231),
.B1(n_230),
.B2(n_220),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_254),
.B(n_208),
.Y(n_266)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_242),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_191),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_246),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_203),
.B(n_164),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_247),
.B(n_218),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_248),
.A2(n_202),
.B1(n_172),
.B2(n_184),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_139),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_250),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_188),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_252),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_196),
.A2(n_170),
.B1(n_145),
.B2(n_141),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_190),
.B1(n_179),
.B2(n_206),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_194),
.B(n_152),
.C(n_145),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_198),
.B(n_209),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_196),
.A2(n_187),
.B1(n_190),
.B2(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_177),
.B(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_177),
.B(n_217),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_176),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_189),
.A2(n_186),
.B1(n_196),
.B2(n_185),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_274),
.C(n_220),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_276),
.B(n_277),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_268),
.A2(n_280),
.B(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_192),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_183),
.B(n_196),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_277),
.B(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_199),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_189),
.A3(n_204),
.B1(n_215),
.B2(n_174),
.C1(n_207),
.C2(n_212),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_229),
.C(n_238),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_282),
.A2(n_286),
.B1(n_291),
.B2(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_239),
.A2(n_202),
.B1(n_181),
.B2(n_197),
.Y(n_286)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_227),
.A2(n_239),
.A3(n_260),
.B1(n_259),
.B2(n_226),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_288),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_253),
.B1(n_221),
.B2(n_256),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_253),
.B1(n_227),
.B2(n_232),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_294),
.A2(n_282),
.B1(n_275),
.B2(n_283),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_244),
.A2(n_233),
.B1(n_243),
.B2(n_235),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_295),
.A2(n_274),
.B1(n_266),
.B2(n_276),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_297),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_304),
.C(n_312),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_309),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_234),
.Y(n_302)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_222),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_303),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_224),
.C(n_238),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_238),
.Y(n_305)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_306),
.A2(n_310),
.B1(n_313),
.B2(n_269),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_252),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_315),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_289),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_285),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_265),
.B(n_262),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_293),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_264),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_318),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_314),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_320),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_268),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_323),
.C(n_280),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_284),
.C(n_275),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_331),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_286),
.B1(n_273),
.B2(n_279),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_328),
.A2(n_340),
.B1(n_343),
.B2(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_337),
.B(n_338),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_299),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_316),
.A2(n_273),
.B1(n_271),
.B2(n_285),
.Y(n_340)
);

OAI22x1_ASAP7_75t_L g341 ( 
.A1(n_307),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_341),
.A2(n_317),
.B1(n_310),
.B2(n_306),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_267),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_344),
.C(n_345),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_296),
.A2(n_272),
.B1(n_285),
.B2(n_301),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_319),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_298),
.B(n_304),
.C(n_323),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_337),
.A2(n_315),
.B1(n_307),
.B2(n_305),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_351),
.B1(n_356),
.B2(n_359),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_332),
.A2(n_311),
.B(n_318),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_361),
.B(n_351),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_341),
.A2(n_299),
.B1(n_317),
.B2(n_297),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_327),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_334),
.B(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_353),
.B(n_362),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_322),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_350),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_355),
.A2(n_329),
.B1(n_335),
.B2(n_362),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_310),
.B1(n_330),
.B2(n_339),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_345),
.C(n_326),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_363),
.C(n_347),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_339),
.B1(n_328),
.B2(n_331),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_343),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_360),
.A2(n_361),
.B1(n_359),
.B2(n_349),
.Y(n_367)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_342),
.C(n_324),
.Y(n_363)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_366),
.B(n_374),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_370),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_356),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_372),
.Y(n_378)
);

INVx11_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_363),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_348),
.Y(n_372)
);

AOI21xp33_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_354),
.B(n_350),
.Y(n_376)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_374),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_370),
.C(n_357),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_382),
.B(n_347),
.C(n_381),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_383),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_SL g385 ( 
.A(n_379),
.B(n_367),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_385),
.A2(n_368),
.B1(n_380),
.B2(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_386),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_387),
.A2(n_384),
.B(n_365),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_389),
.B(n_382),
.Y(n_391)
);

AOI321xp33_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_388),
.A3(n_390),
.B1(n_373),
.B2(n_368),
.C(n_375),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_375),
.B1(n_366),
.B2(n_372),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_369),
.Y(n_394)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_378),
.B(n_364),
.Y(n_395)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_395),
.A2(n_378),
.B(n_364),
.Y(n_396)
);


endmodule