module fake_jpeg_7874_n_17 (n_3, n_2, n_1, n_0, n_4, n_17);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_17;

wire n_13;
wire n_11;
wire n_14;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

INVx1_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

NOR2x1_ASAP7_75t_R g6 ( 
.A(n_1),
.B(n_3),
.Y(n_6)
);

AND2x2_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_2),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_10),
.C(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

AOI22xp5_ASAP7_75t_L g11 ( 
.A1(n_6),
.A2(n_5),
.B1(n_7),
.B2(n_2),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_6),
.B1(n_7),
.B2(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_15),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_1),
.Y(n_15)
);

AOI322xp5_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_4),
.A3(n_11),
.B1(n_14),
.B2(n_15),
.C1(n_10),
.C2(n_9),
.Y(n_17)
);


endmodule