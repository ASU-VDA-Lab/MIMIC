module fake_ariane_1441_n_788 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_788);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_788;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_424;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_557;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_62),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_0),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_11),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_51),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_34),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_25),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_82),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_39),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_22),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_91),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_101),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_74),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_21),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_45),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_90),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_125),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_24),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_93),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_37),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_133),
.Y(n_187)
);

BUFx2_ASAP7_75t_SL g188 ( 
.A(n_56),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_68),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_92),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_20),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_42),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_142),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_0),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_22),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_14),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_140),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_46),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_143),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_1),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_1),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_2),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_2),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_3),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_195),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_157),
.Y(n_222)
);

CKINVDCx6p67_ASAP7_75t_R g223 ( 
.A(n_160),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_5),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_6),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_150),
.B(n_6),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_8),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_9),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_152),
.Y(n_236)
);

BUFx8_ASAP7_75t_SL g237 ( 
.A(n_163),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_152),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_204),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

BUFx8_ASAP7_75t_SL g244 ( 
.A(n_175),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_9),
.Y(n_247)
);

BUFx8_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_199),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_202),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_183),
.B1(n_190),
.B2(n_191),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_210),
.A2(n_149),
.B1(n_201),
.B2(n_200),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_205),
.B1(n_201),
.B2(n_200),
.Y(n_253)
);

AO22x2_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_188),
.B1(n_11),
.B2(n_12),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_10),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_205),
.B1(n_198),
.B2(n_153),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_153),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_209),
.A2(n_198),
.B1(n_194),
.B2(n_187),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_169),
.Y(n_262)
);

AO22x2_ASAP7_75t_L g263 ( 
.A1(n_216),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_184),
.B1(n_182),
.B2(n_180),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_215),
.A2(n_179),
.B1(n_177),
.B2(n_176),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_239),
.Y(n_267)
);

OR2x6_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_13),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_174),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_215),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_240),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_223),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_216),
.A2(n_233),
.B1(n_230),
.B2(n_232),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_233),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

AO22x2_ASAP7_75t_L g277 ( 
.A1(n_227),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_230),
.A2(n_234),
.B1(n_232),
.B2(n_235),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_227),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_29),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_206),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_237),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_30),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_R g289 ( 
.A1(n_247),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_230),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_44),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_148),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_47),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_223),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_R g309 ( 
.A(n_267),
.B(n_241),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_240),
.B(n_241),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_246),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_269),
.Y(n_315)
);

XNOR2x2_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_221),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_248),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_279),
.B(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_257),
.B(n_246),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_255),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_274),
.B(n_246),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_254),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_261),
.B(n_229),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_280),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_R g342 ( 
.A(n_268),
.B(n_234),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_246),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_252),
.B(n_246),
.Y(n_346)
);

BUFx2_ASAP7_75t_R g347 ( 
.A(n_285),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_271),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_244),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_253),
.B(n_246),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_265),
.B(n_248),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_258),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_258),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_302),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_227),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_305),
.B(n_234),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_227),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_235),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_235),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_211),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_315),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_324),
.B(n_225),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_310),
.B(n_211),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_307),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_212),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_225),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_336),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_212),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_347),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_224),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_224),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_344),
.B(n_217),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_217),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_338),
.B(n_224),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_R g403 ( 
.A(n_356),
.B(n_218),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_R g404 ( 
.A(n_357),
.B(n_218),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_335),
.B(n_224),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_320),
.B(n_248),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_248),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_207),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_207),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_231),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g412 ( 
.A(n_346),
.B(n_228),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_346),
.B(n_213),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_353),
.B(n_231),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_353),
.B(n_231),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_298),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_311),
.B(n_327),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_231),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_311),
.B(n_219),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_341),
.B(n_231),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_327),
.B(n_219),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_354),
.B(n_245),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_362),
.B(n_219),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_343),
.A2(n_219),
.B(n_231),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_363),
.B(n_219),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_355),
.B(n_219),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_322),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_369),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_366),
.B(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

BUFx12f_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_358),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_366),
.B(n_354),
.Y(n_442)
);

NAND2x1p5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_333),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_390),
.B(n_323),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_390),
.B(n_395),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_412),
.B(n_316),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_325),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_384),
.B(n_412),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

CKINVDCx8_ASAP7_75t_R g454 ( 
.A(n_406),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_245),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_391),
.B(n_245),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_365),
.B(n_387),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_426),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_319),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_378),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_326),
.Y(n_469)
);

NAND2x1p5_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_334),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_328),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_387),
.B(n_352),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_375),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_373),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_378),
.B(n_206),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_407),
.B(n_213),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_395),
.B(n_213),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_397),
.B(n_219),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_418),
.B(n_213),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_380),
.B(n_213),
.Y(n_486)
);

NAND2x1p5_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_214),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_380),
.B(n_214),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g489 ( 
.A(n_421),
.B(n_214),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_454),
.Y(n_494)
);

INVx3_ASAP7_75t_SL g495 ( 
.A(n_455),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_438),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_395),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

NAND2x1p5_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_430),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_430),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx6_ASAP7_75t_SL g505 ( 
.A(n_455),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_423),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_478),
.Y(n_508)
);

BUFx4f_ASAP7_75t_SL g509 ( 
.A(n_438),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_461),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_485),
.Y(n_512)
);

BUFx2_ASAP7_75t_SL g513 ( 
.A(n_478),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_458),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_452),
.B(n_373),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_457),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_444),
.B(n_397),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_462),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_435),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_457),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_376),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_443),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_465),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_484),
.A2(n_469),
.B(n_486),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_479),
.B(n_415),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_479),
.B(n_377),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_447),
.B(n_398),
.Y(n_535)
);

BUFx2_ASAP7_75t_SL g536 ( 
.A(n_477),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_506),
.Y(n_537)
);

OAI22x1_ASAP7_75t_SL g538 ( 
.A1(n_494),
.A2(n_449),
.B1(n_474),
.B2(n_456),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_521),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_510),
.Y(n_541)
);

CKINVDCx11_ASAP7_75t_R g542 ( 
.A(n_492),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_490),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_530),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_492),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_534),
.A2(n_473),
.B1(n_475),
.B2(n_464),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_449),
.B1(n_440),
.B2(n_441),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_499),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_535),
.A2(n_367),
.B(n_483),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

BUFx12f_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_494),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_507),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_519),
.A2(n_436),
.B1(n_400),
.B2(n_388),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_414),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_514),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_511),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_532),
.A2(n_414),
.B1(n_375),
.B2(n_460),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_509),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_512),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_529),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_528),
.A2(n_428),
.B(n_430),
.Y(n_567)
);

INVx8_ASAP7_75t_L g568 ( 
.A(n_498),
.Y(n_568)
);

OAI21xp33_ASAP7_75t_L g569 ( 
.A1(n_533),
.A2(n_381),
.B(n_383),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_511),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_533),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

CKINVDCx8_ASAP7_75t_R g573 ( 
.A(n_536),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

BUFx8_ASAP7_75t_L g575 ( 
.A(n_520),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_496),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_505),
.A2(n_375),
.B1(n_460),
.B2(n_382),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_520),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_505),
.A2(n_375),
.B1(n_460),
.B2(n_382),
.Y(n_579)
);

INVx8_ASAP7_75t_L g580 ( 
.A(n_498),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_547),
.A2(n_504),
.B1(n_442),
.B2(n_392),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_572),
.A2(n_375),
.B1(n_505),
.B2(n_460),
.Y(n_583)
);

AND2x4_ASAP7_75t_SL g584 ( 
.A(n_541),
.B(n_559),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_539),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_540),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_563),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_549),
.A2(n_375),
.B1(n_460),
.B2(n_410),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_544),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_551),
.A2(n_483),
.B(n_481),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_569),
.A2(n_375),
.B1(n_460),
.B2(n_410),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_568),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_551),
.A2(n_547),
.B1(n_558),
.B2(n_571),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_576),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_548),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_569),
.A2(n_495),
.B1(n_471),
.B2(n_364),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_558),
.A2(n_495),
.B1(n_471),
.B2(n_364),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_504),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_552),
.B(n_524),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_L g601 ( 
.A1(n_557),
.A2(n_564),
.B(n_566),
.Y(n_601)
);

BUFx12f_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_557),
.A2(n_393),
.B1(n_368),
.B2(n_401),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_537),
.B(n_524),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_538),
.A2(n_525),
.B1(n_498),
.B2(n_536),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_562),
.A2(n_525),
.B1(n_450),
.B2(n_446),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_565),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_574),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_554),
.A2(n_405),
.B(n_376),
.Y(n_611)
);

AOI21xp33_ASAP7_75t_L g612 ( 
.A1(n_577),
.A2(n_488),
.B(n_528),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_578),
.Y(n_613)
);

INVx5_ASAP7_75t_SL g614 ( 
.A(n_541),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_560),
.A2(n_393),
.B1(n_401),
.B2(n_368),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_546),
.A2(n_416),
.B1(n_415),
.B2(n_526),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_537),
.B(n_480),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_541),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_559),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_553),
.A2(n_400),
.B1(n_392),
.B2(n_416),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_546),
.A2(n_513),
.B1(n_419),
.B2(n_389),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_579),
.A2(n_419),
.B1(n_467),
.B2(n_463),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_568),
.A2(n_472),
.B1(n_467),
.B2(n_463),
.Y(n_624)
);

OAI222xp33_ASAP7_75t_L g625 ( 
.A1(n_573),
.A2(n_408),
.B1(n_459),
.B2(n_472),
.C1(n_453),
.C2(n_389),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_561),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_575),
.A2(n_513),
.B1(n_404),
.B2(n_403),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_568),
.A2(n_459),
.B1(n_379),
.B2(n_446),
.Y(n_630)
);

OAI221xp5_ASAP7_75t_SL g631 ( 
.A1(n_593),
.A2(n_405),
.B1(n_399),
.B2(n_394),
.C(n_433),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_588),
.A2(n_379),
.B1(n_453),
.B2(n_482),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_588),
.A2(n_379),
.B1(n_482),
.B2(n_545),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_596),
.A2(n_379),
.B1(n_545),
.B2(n_450),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_596),
.A2(n_411),
.B1(n_575),
.B2(n_409),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_597),
.A2(n_409),
.B1(n_413),
.B2(n_570),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_600),
.B(n_543),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_582),
.A2(n_580),
.B1(n_404),
.B2(n_403),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_597),
.A2(n_413),
.B1(n_214),
.B2(n_580),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_593),
.A2(n_413),
.B1(n_214),
.B2(n_580),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_616),
.A2(n_214),
.B1(n_508),
.B2(n_372),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_590),
.A2(n_581),
.B1(n_543),
.B2(n_508),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_610),
.A2(n_617),
.B1(n_621),
.B2(n_583),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_621),
.A2(n_372),
.B1(n_399),
.B2(n_394),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_611),
.A2(n_376),
.B1(n_470),
.B2(n_443),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_608),
.A2(n_430),
.B1(n_517),
.B2(n_522),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_583),
.A2(n_374),
.B1(n_567),
.B2(n_517),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_615),
.A2(n_601),
.B1(n_623),
.B2(n_612),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_615),
.A2(n_623),
.B1(n_606),
.B2(n_604),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_543),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_591),
.A2(n_374),
.B1(n_567),
.B2(n_517),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_585),
.A2(n_581),
.B1(n_543),
.B2(n_517),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_607),
.A2(n_376),
.B1(n_470),
.B2(n_522),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_591),
.A2(n_374),
.B1(n_489),
.B2(n_487),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_586),
.A2(n_581),
.B1(n_518),
.B2(n_527),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_589),
.A2(n_581),
.B1(n_518),
.B2(n_527),
.Y(n_656)
);

OAI222xp33_ASAP7_75t_L g657 ( 
.A1(n_622),
.A2(n_489),
.B1(n_487),
.B2(n_531),
.C1(n_518),
.C2(n_527),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_630),
.A2(n_522),
.B1(n_500),
.B2(n_501),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_603),
.A2(n_476),
.B1(n_422),
.B2(n_531),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_603),
.A2(n_476),
.B1(n_531),
.B2(n_503),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_605),
.B(n_490),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_599),
.A2(n_476),
.B1(n_503),
.B2(n_493),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_630),
.A2(n_500),
.B1(n_501),
.B2(n_516),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_624),
.A2(n_476),
.B1(n_503),
.B2(n_493),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_613),
.B(n_490),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_624),
.A2(n_594),
.B1(n_598),
.B2(n_628),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_602),
.A2(n_490),
.B1(n_503),
.B2(n_491),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_595),
.A2(n_491),
.B1(n_503),
.B2(n_493),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_595),
.A2(n_493),
.B1(n_491),
.B2(n_424),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_592),
.A2(n_501),
.B1(n_500),
.B2(n_516),
.Y(n_670)
);

OAI21xp33_ASAP7_75t_L g671 ( 
.A1(n_631),
.A2(n_629),
.B(n_627),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_665),
.B(n_618),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_637),
.B(n_620),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_648),
.A2(n_614),
.B1(n_626),
.B2(n_592),
.Y(n_674)
);

NAND4xp25_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_587),
.C(n_619),
.D(n_431),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_SL g676 ( 
.A(n_666),
.B(n_587),
.C(n_614),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_640),
.A2(n_625),
.B(n_425),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_665),
.B(n_584),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g679 ( 
.A1(n_638),
.A2(n_584),
.B(n_592),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_650),
.B(n_614),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_661),
.B(n_592),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_661),
.B(n_427),
.C(n_420),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_643),
.B(n_491),
.Y(n_683)
);

AND2x2_ASAP7_75t_SL g684 ( 
.A(n_634),
.B(n_491),
.Y(n_684)
);

NAND4xp25_ASAP7_75t_SL g685 ( 
.A(n_645),
.B(n_48),
.C(n_49),
.D(n_50),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_656),
.B(n_493),
.C(n_516),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_667),
.B(n_516),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_642),
.B(n_516),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_655),
.B(n_425),
.C(n_53),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_646),
.B(n_52),
.C(n_54),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_649),
.B(n_55),
.Y(n_691)
);

NAND4xp25_ASAP7_75t_L g692 ( 
.A(n_635),
.B(n_645),
.C(n_644),
.D(n_636),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_647),
.B(n_669),
.C(n_651),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_668),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_664),
.B(n_652),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_659),
.B(n_633),
.C(n_662),
.Y(n_696)
);

AOI221xp5_ASAP7_75t_L g697 ( 
.A1(n_641),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_639),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_698)
);

NAND4xp25_ASAP7_75t_L g699 ( 
.A(n_653),
.B(n_146),
.C(n_69),
.D(n_70),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_660),
.B(n_67),
.C(n_71),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_675),
.A2(n_632),
.B1(n_654),
.B2(n_658),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_663),
.C(n_670),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_673),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_672),
.B(n_72),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_678),
.B(n_75),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_680),
.B(n_76),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_694),
.B(n_77),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_683),
.B(n_78),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_681),
.B(n_79),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_676),
.A2(n_685),
.B(n_699),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_692),
.A2(n_657),
.B1(n_84),
.B2(n_85),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_695),
.B(n_81),
.Y(n_712)
);

AND4x1_ASAP7_75t_L g713 ( 
.A(n_686),
.B(n_86),
.C(n_87),
.D(n_88),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_693),
.B(n_89),
.Y(n_714)
);

AOI221xp5_ASAP7_75t_L g715 ( 
.A1(n_691),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.C(n_99),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_684),
.B(n_100),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_691),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_696),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_703),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_714),
.Y(n_720)
);

XOR2x2_ASAP7_75t_L g721 ( 
.A(n_710),
.B(n_700),
.Y(n_721)
);

NAND4xp75_ASAP7_75t_L g722 ( 
.A(n_716),
.B(n_688),
.C(n_687),
.D(n_697),
.Y(n_722)
);

NAND4xp75_ASAP7_75t_SL g723 ( 
.A(n_716),
.B(n_679),
.C(n_674),
.D(n_690),
.Y(n_723)
);

XNOR2xp5_ASAP7_75t_L g724 ( 
.A(n_704),
.B(n_698),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_703),
.B(n_671),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_717),
.Y(n_726)
);

NAND4xp75_ASAP7_75t_SL g727 ( 
.A(n_704),
.B(n_708),
.C(n_709),
.D(n_706),
.Y(n_727)
);

NAND4xp75_ASAP7_75t_SL g728 ( 
.A(n_708),
.B(n_709),
.C(n_706),
.D(n_713),
.Y(n_728)
);

NAND4xp25_ASAP7_75t_L g729 ( 
.A(n_714),
.B(n_682),
.C(n_677),
.D(n_698),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_707),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_725),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_720),
.B(n_712),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_725),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_726),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_730),
.B(n_702),
.Y(n_735)
);

XNOR2xp5_ASAP7_75t_L g736 ( 
.A(n_721),
.B(n_711),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_736),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_731),
.Y(n_738)
);

OA22x2_ASAP7_75t_L g739 ( 
.A1(n_736),
.A2(n_724),
.B1(n_721),
.B2(n_730),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_735),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_740),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_738),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_739),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_743),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_742),
.Y(n_746)
);

AOI22x1_ASAP7_75t_L g747 ( 
.A1(n_741),
.A2(n_734),
.B1(n_735),
.B2(n_739),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_746),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_737),
.B1(n_743),
.B2(n_744),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_745),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_745),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_749),
.A2(n_743),
.B1(n_729),
.B2(n_750),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_749),
.B(n_743),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_749),
.A2(n_733),
.B1(n_732),
.B2(n_722),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_754),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_756),
.A2(n_715),
.B1(n_705),
.B2(n_707),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_752),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_754),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_761),
.A2(n_718),
.B(n_723),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_757),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_719),
.B1(n_701),
.B2(n_728),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_758),
.A2(n_759),
.B1(n_762),
.B2(n_719),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_761),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_765),
.A2(n_719),
.B1(n_727),
.B2(n_689),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_767),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_764),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_763),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_766),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_767),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_769),
.A2(n_677),
.B1(n_107),
.B2(n_108),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_771),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_775)
);

AO22x2_ASAP7_75t_L g776 ( 
.A1(n_772),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_770),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_776),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_777),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_774),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_779),
.B1(n_778),
.B2(n_773),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_780),
.A2(n_768),
.B1(n_775),
.B2(n_122),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_780),
.A2(n_144),
.B1(n_121),
.B2(n_124),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_781),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_784),
.A2(n_782),
.B1(n_783),
.B2(n_128),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_785),
.Y(n_786)
);

AOI221xp5_ASAP7_75t_L g787 ( 
.A1(n_786),
.A2(n_120),
.B1(n_126),
.B2(n_129),
.C(n_130),
.Y(n_787)
);

AOI211xp5_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_132),
.B(n_134),
.C(n_136),
.Y(n_788)
);


endmodule