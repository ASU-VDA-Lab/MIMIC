module fake_jpeg_8122_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

OR2x2_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_10),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_12)
);

NOR2xp67_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_16),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_3),
.B(n_5),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_1),
.Y(n_15)
);

XOR2x1_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_2),
.Y(n_16)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_1),
.B(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_13),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_22),
.B(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_16),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_15),
.B(n_17),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_32)
);

MAJx2_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.C(n_7),
.Y(n_34)
);

NAND5xp2_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_17),
.C(n_7),
.D(n_8),
.E(n_9),
.Y(n_33)
);

OAI321xp33_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.A3(n_33),
.B1(n_32),
.B2(n_31),
.C(n_5),
.Y(n_36)
);

OAI321xp33_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_14),
.C(n_31),
.Y(n_35)
);


endmodule