module real_aes_15478_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_845, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_845;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_0), .Y(n_173) );
AND2x4_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g224 ( .A(n_2), .Y(n_224) );
INVx1_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_4), .A2(n_144), .B1(n_839), .B2(n_840), .Y(n_838) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_4), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_5), .B(n_232), .Y(n_231) );
BUFx2_ASAP7_75t_L g115 ( .A(n_6), .Y(n_115) );
OR2x2_ASAP7_75t_L g126 ( .A(n_6), .B(n_23), .Y(n_126) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_7), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_8), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_9), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_9), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_10), .B(n_194), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_11), .B(n_194), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_12), .B(n_154), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_13), .A2(n_80), .B1(n_191), .B2(n_194), .Y(n_193) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_14), .A2(n_36), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_15), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_16), .B(n_163), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_17), .Y(n_566) );
AO32x1_ASAP7_75t_L g185 ( .A1(n_18), .A2(n_186), .A3(n_187), .B1(n_196), .B2(n_198), .Y(n_185) );
AO32x2_ASAP7_75t_L g302 ( .A1(n_18), .A2(n_186), .A3(n_187), .B1(n_196), .B2(n_198), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_19), .B(n_526), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_20), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_21), .B(n_198), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_22), .Y(n_641) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_23), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_24), .A2(n_42), .B1(n_163), .B2(n_165), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_25), .A2(n_88), .B1(n_191), .B2(n_192), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_26), .B(n_234), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_27), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_28), .B(n_259), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_29), .A2(n_62), .B1(n_192), .B2(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_30), .B(n_194), .Y(n_512) );
INVx2_ASAP7_75t_L g132 ( .A(n_31), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_32), .B(n_195), .Y(n_522) );
INVx1_ASAP7_75t_L g105 ( .A(n_33), .Y(n_105) );
BUFx3_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_34), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_35), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g571 ( .A(n_37), .B(n_531), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_38), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_39), .B(n_174), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_40), .B(n_526), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_41), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_43), .B(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_44), .A2(n_75), .B1(n_174), .B2(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_45), .B(n_203), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_46), .A2(n_171), .B(n_188), .C(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_47), .A2(n_77), .B1(n_191), .B2(n_194), .Y(n_220) );
INVx1_ASAP7_75t_L g158 ( .A(n_48), .Y(n_158) );
AND2x4_ASAP7_75t_L g178 ( .A(n_49), .B(n_179), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_50), .A2(n_51), .B1(n_165), .B2(n_192), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_52), .B(n_198), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_53), .B(n_531), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_54), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_55), .A2(n_100), .B1(n_116), .B2(n_842), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_56), .B(n_192), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_57), .B(n_191), .Y(n_230) );
INVx1_ASAP7_75t_L g179 ( .A(n_58), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_59), .B(n_198), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_60), .A2(n_171), .B(n_172), .C(n_175), .Y(n_170) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_61), .B(n_191), .C(n_236), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_63), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_64), .B(n_198), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_65), .B(n_515), .Y(n_553) );
AND2x2_ASAP7_75t_L g180 ( .A(n_66), .B(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_67), .Y(n_208) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_68), .B(n_163), .C(n_195), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_69), .A2(n_91), .B1(n_174), .B2(n_194), .Y(n_261) );
INVx2_ASAP7_75t_L g169 ( .A(n_70), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_71), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_72), .B(n_515), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_73), .B(n_168), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_74), .B(n_194), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_76), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_78), .B(n_251), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_79), .A2(n_87), .B1(n_526), .B2(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_81), .B(n_194), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_82), .B(n_236), .Y(n_235) );
NAND2xp33_ASAP7_75t_SL g594 ( .A(n_83), .B(n_232), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_84), .B(n_247), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_85), .A2(n_98), .B1(n_165), .B2(n_192), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_86), .B(n_259), .Y(n_277) );
INVx1_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_89), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_90), .B(n_154), .Y(n_283) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_92), .B(n_232), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_93), .B(n_531), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_94), .B(n_168), .C(n_232), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_95), .B(n_515), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_96), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_97), .B(n_526), .Y(n_556) );
CKINVDCx11_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx11_ASAP7_75t_R g843 ( .A(n_101), .Y(n_843) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_111), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NOR2x1p5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND3x2_ASAP7_75t_L g836 ( .A(n_104), .B(n_107), .C(n_125), .Y(n_836) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g124 ( .A(n_105), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g143 ( .A(n_108), .Y(n_143) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1p5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_127), .Y(n_116) );
INVxp67_ASAP7_75t_L g841 ( .A(n_117), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_SL g122 ( .A(n_123), .B(n_125), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_125), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2x1_ASAP7_75t_L g828 ( .A(n_126), .B(n_135), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_829), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_821), .Y(n_128) );
BUFx12f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x6_ASAP7_75t_SL g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_132), .B(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g832 ( .A(n_132), .Y(n_832) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B1(n_499), .B2(n_501), .Y(n_141) );
BUFx12f_ASAP7_75t_L g500 ( .A(n_142), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g827 ( .A(n_143), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g840 ( .A(n_144), .Y(n_840) );
NAND4xp75_ASAP7_75t_L g144 ( .A(n_145), .B(n_373), .C(n_427), .D(n_471), .Y(n_144) );
NOR2x1_ASAP7_75t_L g145 ( .A(n_146), .B(n_326), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_292), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_209), .B(n_213), .C(n_265), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_183), .Y(n_148) );
AND2x2_ASAP7_75t_L g343 ( .A(n_149), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g332 ( .A(n_150), .B(n_268), .Y(n_332) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_151), .Y(n_298) );
AND2x2_ASAP7_75t_L g347 ( .A(n_151), .B(n_199), .Y(n_347) );
INVx1_ASAP7_75t_L g359 ( .A(n_151), .Y(n_359) );
INVx1_ASAP7_75t_L g457 ( .A(n_151), .Y(n_457) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g211 ( .A(n_152), .Y(n_211) );
AOI21x1_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_159), .B(n_180), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp67_ASAP7_75t_SL g561 ( .A(n_154), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_155), .A2(n_533), .A3(n_538), .B(n_539), .Y(n_532) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
INVx2_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_170), .B(n_177), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_161), .B(n_167), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B1(n_165), .B2(n_166), .Y(n_161) );
INVx2_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_164), .Y(n_165) );
INVx1_ASAP7_75t_L g171 ( .A(n_164), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_164), .Y(n_174) );
INVx2_ASAP7_75t_L g191 ( .A(n_164), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_164), .Y(n_232) );
INVx1_ASAP7_75t_L g247 ( .A(n_164), .Y(n_247) );
INVx3_ASAP7_75t_L g515 ( .A(n_164), .Y(n_515) );
INVx1_ASAP7_75t_L g527 ( .A(n_164), .Y(n_527) );
INVx1_ASAP7_75t_L g253 ( .A(n_165), .Y(n_253) );
AOI21x1_ASAP7_75t_L g524 ( .A1(n_167), .A2(n_525), .B(n_528), .Y(n_524) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_SL g260 ( .A(n_168), .Y(n_260) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
INVx1_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
BUFx8_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
INVx1_ASAP7_75t_L g582 ( .A(n_171), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
INVx2_ASAP7_75t_L g537 ( .A(n_175), .Y(n_537) );
BUFx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g252 ( .A(n_176), .Y(n_252) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g197 ( .A(n_178), .Y(n_197) );
AO31x2_ASAP7_75t_L g199 ( .A1(n_178), .A2(n_200), .A3(n_201), .B(n_207), .Y(n_199) );
BUFx10_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
BUFx10_ASAP7_75t_L g538 ( .A(n_178), .Y(n_538) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_182), .B(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_182), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g285 ( .A(n_184), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_199), .Y(n_184) );
AND2x2_ASAP7_75t_L g212 ( .A(n_185), .B(n_199), .Y(n_212) );
INVx1_ASAP7_75t_L g325 ( .A(n_185), .Y(n_325) );
INVx1_ASAP7_75t_L g436 ( .A(n_185), .Y(n_436) );
INVx4_ASAP7_75t_L g198 ( .A(n_186), .Y(n_198) );
BUFx3_ASAP7_75t_L g200 ( .A(n_186), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_186), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_186), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g242 ( .A(n_186), .Y(n_242) );
INVx2_ASAP7_75t_SL g274 ( .A(n_186), .Y(n_274) );
AND2x4_ASAP7_75t_SL g584 ( .A(n_186), .B(n_218), .Y(n_584) );
INVx1_ASAP7_75t_SL g587 ( .A(n_186), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B1(n_193), .B2(n_195), .Y(n_187) );
O2A1O1Ixp5_ASAP7_75t_L g244 ( .A1(n_188), .A2(n_245), .B(n_246), .C(n_248), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_188), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_188), .A2(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_188), .A2(n_578), .B(n_579), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_188), .A2(n_593), .B(n_594), .Y(n_592) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g236 ( .A(n_189), .Y(n_236) );
INVx2_ASAP7_75t_SL g259 ( .A(n_191), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_191), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g234 ( .A(n_192), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_192), .A2(n_522), .B(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g535 ( .A(n_192), .Y(n_535) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_192), .A2(n_515), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx3_ASAP7_75t_L g282 ( .A(n_194), .Y(n_282) );
INVx1_ASAP7_75t_L g529 ( .A(n_194), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_194), .A2(n_590), .B(n_591), .Y(n_589) );
INVx6_ASAP7_75t_L g204 ( .A(n_195), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_195), .A2(n_204), .B1(n_220), .B2(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_195), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_195), .A2(n_514), .B(n_516), .Y(n_513) );
O2A1O1Ixp5_ASAP7_75t_L g640 ( .A1(n_195), .A2(n_246), .B(n_641), .C(n_642), .Y(n_640) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_196), .A2(n_276), .B(n_279), .Y(n_275) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_SL g262 ( .A(n_197), .Y(n_262) );
INVx2_ASAP7_75t_L g217 ( .A(n_198), .Y(n_217) );
INVx3_ASAP7_75t_L g268 ( .A(n_199), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_199), .B(n_272), .Y(n_323) );
AND2x2_ASAP7_75t_L g358 ( .A(n_199), .B(n_359), .Y(n_358) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_200), .A2(n_257), .A3(n_262), .B(n_263), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B1(n_205), .B2(n_206), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_204), .A2(n_258), .B1(n_260), .B2(n_261), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_204), .A2(n_280), .B(n_281), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_204), .A2(n_534), .B1(n_536), .B2(n_537), .Y(n_533) );
AOI21x1_ASAP7_75t_L g276 ( .A1(n_206), .A2(n_277), .B(n_278), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_206), .A2(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
INVx1_ASAP7_75t_L g398 ( .A(n_210), .Y(n_398) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g267 ( .A(n_211), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_211), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
OR2x2_ASAP7_75t_L g364 ( .A(n_211), .B(n_272), .Y(n_364) );
OR2x2_ASAP7_75t_L g435 ( .A(n_211), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g372 ( .A(n_212), .Y(n_372) );
AND2x2_ASAP7_75t_L g424 ( .A(n_212), .B(n_287), .Y(n_424) );
AND2x2_ASAP7_75t_L g481 ( .A(n_212), .B(n_398), .Y(n_481) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_239), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_214), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g490 ( .A(n_214), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
INVx2_ASAP7_75t_L g291 ( .A(n_215), .Y(n_291) );
AND2x2_ASAP7_75t_L g316 ( .A(n_215), .B(n_295), .Y(n_316) );
AND2x2_ASAP7_75t_L g386 ( .A(n_215), .B(n_256), .Y(n_386) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g340 ( .A(n_216), .Y(n_340) );
AOI31xp67_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .A3(n_219), .B(n_222), .Y(n_216) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_218), .A2(n_229), .B(n_233), .Y(n_228) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_218), .A2(n_244), .B(n_249), .Y(n_243) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_218), .A2(n_510), .B(n_513), .Y(n_509) );
OAI21x1_ASAP7_75t_L g520 ( .A1(n_218), .A2(n_521), .B(n_524), .Y(n_520) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_218), .A2(n_552), .B(n_555), .Y(n_551) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_218), .A2(n_589), .B(n_592), .Y(n_588) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_218), .A2(n_640), .B(n_643), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g294 ( .A(n_225), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g355 ( .A(n_225), .B(n_241), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_228), .B(n_238), .Y(n_225) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_226), .A2(n_228), .B(n_238), .Y(n_311) );
OAI21xp33_ASAP7_75t_SL g550 ( .A1(n_226), .A2(n_551), .B(n_558), .Y(n_550) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_226), .A2(n_551), .B(n_558), .Y(n_620) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_226), .A2(n_639), .B(n_647), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_226), .A2(n_639), .B(n_647), .Y(n_670) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g531 ( .A(n_227), .Y(n_531) );
INVx2_ASAP7_75t_L g646 ( .A(n_232), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .Y(n_233) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g362 ( .A(n_240), .B(n_339), .Y(n_362) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_256), .Y(n_240) );
INVx2_ASAP7_75t_SL g284 ( .A(n_241), .Y(n_284) );
BUFx2_ASAP7_75t_L g337 ( .A(n_241), .Y(n_337) );
INVx1_ASAP7_75t_L g409 ( .A(n_241), .Y(n_409) );
AND2x2_ASAP7_75t_L g442 ( .A(n_241), .B(n_290), .Y(n_442) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_255), .Y(n_241) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_242), .A2(n_243), .B(n_255), .Y(n_295) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_242), .A2(n_509), .B(n_517), .Y(n_508) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_242), .A2(n_520), .B(n_530), .Y(n_519) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_242), .A2(n_509), .B(n_517), .Y(n_600) );
OA21x2_ASAP7_75t_L g635 ( .A1(n_242), .A2(n_520), .B(n_530), .Y(n_635) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_252), .B1(n_253), .B2(n_254), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_251), .A2(n_644), .B(n_645), .Y(n_643) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_252), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_580) );
INVx2_ASAP7_75t_L g270 ( .A(n_256), .Y(n_270) );
INVx1_ASAP7_75t_L g290 ( .A(n_256), .Y(n_290) );
INVx1_ASAP7_75t_L g318 ( .A(n_256), .Y(n_318) );
AND2x2_ASAP7_75t_L g408 ( .A(n_256), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g449 ( .A(n_256), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g465 ( .A(n_256), .B(n_450), .Y(n_465) );
AND2x2_ASAP7_75t_L g491 ( .A(n_256), .B(n_295), .Y(n_491) );
OAI32xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .A3(n_284), .B1(n_285), .B2(n_288), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_267), .B(n_432), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_267), .B(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g301 ( .A(n_268), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g403 ( .A(n_268), .Y(n_403) );
INVx1_ASAP7_75t_L g463 ( .A(n_268), .Y(n_463) );
INVx1_ASAP7_75t_L g401 ( .A(n_269), .Y(n_401) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_SL g305 ( .A(n_270), .Y(n_305) );
AND2x2_ASAP7_75t_L g394 ( .A(n_270), .B(n_309), .Y(n_394) );
AND2x2_ASAP7_75t_L g462 ( .A(n_271), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g287 ( .A(n_272), .Y(n_287) );
AND2x2_ASAP7_75t_L g297 ( .A(n_272), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
AND2x2_ASAP7_75t_L g344 ( .A(n_272), .B(n_302), .Y(n_344) );
AND2x2_ASAP7_75t_L g368 ( .A(n_272), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g378 ( .A(n_272), .B(n_369), .Y(n_378) );
INVxp67_ASAP7_75t_L g432 ( .A(n_272), .Y(n_432) );
BUFx2_ASAP7_75t_L g444 ( .A(n_272), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_272), .Y(n_448) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B(n_283), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_284), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g440 ( .A(n_284), .Y(n_440) );
AND2x2_ASAP7_75t_L g348 ( .A(n_287), .B(n_325), .Y(n_348) );
AND2x2_ASAP7_75t_L g477 ( .A(n_287), .B(n_301), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g365 ( .A1(n_288), .A2(n_366), .B1(n_370), .B2(n_371), .Y(n_365) );
O2A1O1Ixp5_ASAP7_75t_R g439 ( .A1(n_288), .A2(n_440), .B(n_441), .C(n_443), .Y(n_439) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g293 ( .A(n_289), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g307 ( .A(n_291), .Y(n_307) );
INVx1_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_291), .B(n_320), .Y(n_426) );
AND2x2_ASAP7_75t_L g438 ( .A(n_291), .B(n_309), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B1(n_299), .B2(n_303), .C1(n_313), .C2(n_321), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_293), .A2(n_335), .B1(n_413), .B2(n_474), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_293), .A2(n_357), .B1(n_493), .B2(n_495), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_294), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_294), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g468 ( .A(n_294), .Y(n_468) );
INVx1_ASAP7_75t_L g498 ( .A(n_294), .Y(n_498) );
INVx1_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
AOI321xp33_ASAP7_75t_L g445 ( .A1(n_299), .A2(n_343), .A3(n_446), .B1(n_451), .B2(n_452), .C(n_453), .Y(n_445) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
OR2x2_ASAP7_75t_L g377 ( .A(n_300), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g397 ( .A(n_301), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g369 ( .A(n_302), .Y(n_369) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
OR2x2_ASAP7_75t_L g370 ( .A(n_305), .B(n_339), .Y(n_370) );
AND2x2_ASAP7_75t_L g390 ( .A(n_305), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g480 ( .A(n_306), .Y(n_480) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g411 ( .A(n_308), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g320 ( .A(n_310), .Y(n_320) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g339 ( .A(n_311), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_314), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_316), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g451 ( .A(n_320), .Y(n_451) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_322), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g384 ( .A(n_323), .Y(n_384) );
INVx1_ASAP7_75t_L g334 ( .A(n_324), .Y(n_334) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_325), .Y(n_382) );
INVx2_ASAP7_75t_L g416 ( .A(n_325), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_351), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_335), .B(n_341), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_330), .B(n_334), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_331), .A2(n_418), .B1(n_468), .B2(n_469), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g433 ( .A(n_332), .Y(n_433) );
AND2x2_ASAP7_75t_L g357 ( .A(n_333), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g371 ( .A(n_333), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g422 ( .A(n_333), .Y(n_422) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g402 ( .A(n_337), .B(n_338), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_337), .B(n_386), .Y(n_418) );
AND2x2_ASAP7_75t_L g464 ( .A(n_337), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_338), .B(n_442), .Y(n_479) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g391 ( .A(n_339), .Y(n_391) );
INVx1_ASAP7_75t_L g450 ( .A(n_340), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B(n_349), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g412 ( .A(n_344), .B(n_367), .Y(n_412) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_347), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g421 ( .A(n_347), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_350), .B(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_365), .Y(n_351) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_360), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_353), .A2(n_420), .B1(n_423), .B2(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI311xp33_ASAP7_75t_L g453 ( .A1(n_355), .A2(n_454), .A3(n_455), .B(n_458), .C(n_459), .Y(n_453) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g381 ( .A(n_358), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_358), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g452 ( .A(n_362), .Y(n_452) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g458 ( .A(n_368), .Y(n_458) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_372), .Y(n_475) );
NOR2x1_ASAP7_75t_L g373 ( .A(n_374), .B(n_399), .Y(n_373) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_379), .C(n_387), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AO21x1_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B(n_385), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AO221x1_ASAP7_75t_L g460 ( .A1(n_381), .A2(n_461), .B1(n_464), .B2(n_466), .C(n_467), .Y(n_460) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g459 ( .A(n_386), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B(n_395), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B(n_404), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g454 ( .A(n_403), .Y(n_454) );
AOI221x1_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_412), .B1(n_413), .B2(n_417), .C(n_419), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_410), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g437 ( .A(n_408), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AO22x1_ASAP7_75t_L g484 ( .A1(n_412), .A2(n_485), .B1(n_487), .B2(n_490), .Y(n_484) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g461 ( .A(n_415), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_416), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp33_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_460), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_445), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_437), .B(n_439), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .C(n_435), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
AND2x2_ASAP7_75t_L g456 ( .A(n_436), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g466 ( .A(n_442), .B(n_451), .Y(n_466) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_448), .B(n_456), .Y(n_494) );
INVx2_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g489 ( .A(n_457), .Y(n_489) );
AND2x2_ASAP7_75t_L g485 ( .A(n_465), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g497 ( .A(n_465), .Y(n_497) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_478), .B1(n_480), .B2(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx4_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2x1p5_ASAP7_75t_SL g501 ( .A(n_502), .B(n_755), .Y(n_501) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_691), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_504), .B(n_612), .C(n_652), .D(n_681), .Y(n_503) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_541), .B(n_548), .C(n_596), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_518), .Y(n_505) );
INVx2_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
AND2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_506), .B(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_506), .B(n_598), .Y(n_774) );
OR2x2_ASAP7_75t_L g810 ( .A(n_506), .B(n_726), .Y(n_810) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g707 ( .A(n_507), .B(n_519), .Y(n_707) );
NOR2xp67_ASAP7_75t_L g733 ( .A(n_507), .B(n_546), .Y(n_733) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g668 ( .A(n_508), .Y(n_668) );
AND2x2_ASAP7_75t_L g606 ( .A(n_518), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_518), .B(n_636), .Y(n_651) );
AND2x2_ASAP7_75t_L g659 ( .A(n_518), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_518), .Y(n_682) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_532), .Y(n_518) );
INVx1_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
INVx1_ASAP7_75t_L g598 ( .A(n_519), .Y(n_598) );
AND2x2_ASAP7_75t_L g669 ( .A(n_519), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g730 ( .A(n_519), .B(n_637), .Y(n_730) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g547 ( .A(n_532), .Y(n_547) );
AND2x2_ASAP7_75t_L g599 ( .A(n_532), .B(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_532), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_532), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g713 ( .A(n_532), .B(n_668), .Y(n_713) );
OR2x2_ASAP7_75t_L g726 ( .A(n_532), .B(n_635), .Y(n_726) );
OR2x2_ASAP7_75t_L g736 ( .A(n_532), .B(n_600), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_537), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_544), .B(n_752), .Y(n_798) );
INVx1_ASAP7_75t_L g654 ( .A(n_545), .Y(n_654) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x2_ASAP7_75t_L g738 ( .A(n_547), .B(n_600), .Y(n_738) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_572), .Y(n_548) );
AND2x2_ASAP7_75t_L g610 ( .A(n_549), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g673 ( .A(n_549), .Y(n_673) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_559), .Y(n_549) );
BUFx2_ASAP7_75t_L g780 ( .A(n_550), .Y(n_780) );
AND2x2_ASAP7_75t_L g618 ( .A(n_559), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g604 ( .A(n_560), .B(n_586), .Y(n_604) );
INVx2_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
AOI21x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B(n_571), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
AND2x2_ASAP7_75t_L g777 ( .A(n_572), .B(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_585), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx4_ASAP7_75t_L g603 ( .A(n_574), .Y(n_603) );
BUFx2_ASAP7_75t_L g611 ( .A(n_574), .Y(n_611) );
OR2x2_ASAP7_75t_L g615 ( .A(n_574), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g676 ( .A(n_574), .B(n_619), .Y(n_676) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B(n_584), .Y(n_576) );
INVx1_ASAP7_75t_L g663 ( .A(n_585), .Y(n_663) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_585), .Y(n_677) );
INVx2_ASAP7_75t_L g702 ( .A(n_585), .Y(n_702) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g616 ( .A(n_586), .Y(n_616) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_595), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B1(n_605), .B2(n_609), .Y(n_596) );
INVx1_ASAP7_75t_L g687 ( .A(n_597), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g698 ( .A(n_598), .Y(n_698) );
AND2x2_ASAP7_75t_L g715 ( .A(n_599), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_599), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g608 ( .A(n_600), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_601), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_602), .B(n_618), .Y(n_710) );
AND2x2_ASAP7_75t_L g718 ( .A(n_602), .B(n_684), .Y(n_718) );
AND2x2_ASAP7_75t_L g794 ( .A(n_602), .B(n_741), .Y(n_794) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g628 ( .A(n_603), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g650 ( .A(n_603), .B(n_619), .Y(n_650) );
OR2x2_ASAP7_75t_L g662 ( .A(n_603), .B(n_663), .Y(n_662) );
NAND2x1_ASAP7_75t_L g696 ( .A(n_603), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g701 ( .A(n_603), .Y(n_701) );
INVx2_ASAP7_75t_L g695 ( .A(n_604), .Y(n_695) );
AND2x2_ASAP7_75t_L g721 ( .A(n_604), .B(n_685), .Y(n_721) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_607), .Y(n_657) );
INVx1_ASAP7_75t_L g724 ( .A(n_607), .Y(n_724) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g708 ( .A(n_608), .B(n_637), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_609), .A2(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g781 ( .A(n_611), .B(n_721), .Y(n_781) );
INVx1_ASAP7_75t_L g817 ( .A(n_611), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_621), .B(n_625), .Y(n_612) );
AOI322xp5_ASAP7_75t_L g765 ( .A1(n_613), .A2(n_661), .A3(n_766), .B1(n_767), .B2(n_768), .C1(n_769), .C2(n_772), .Y(n_765) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_615), .B(n_617), .C(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g631 ( .A(n_616), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g761 ( .A(n_616), .B(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_616), .Y(n_813) );
OR2x2_ASAP7_75t_L g709 ( .A(n_617), .B(n_662), .Y(n_709) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g697 ( .A(n_619), .Y(n_697) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g632 ( .A(n_620), .Y(n_632) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_622), .Y(n_758) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g729 ( .A(n_623), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g792 ( .A(n_624), .B(n_752), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_633), .B(n_648), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_627), .B(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
AND2x2_ASAP7_75t_L g684 ( .A(n_629), .B(n_685), .Y(n_684) );
AND3x2_ASAP7_75t_L g728 ( .A(n_629), .B(n_631), .C(n_701), .Y(n_728) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g690 ( .A(n_630), .Y(n_690) );
AND2x2_ASAP7_75t_L g741 ( .A(n_630), .B(n_702), .Y(n_741) );
INVx2_ASAP7_75t_L g764 ( .A(n_630), .Y(n_764) );
AND2x2_ASAP7_75t_L g768 ( .A(n_631), .B(n_764), .Y(n_768) );
INVx2_ASAP7_75t_L g685 ( .A(n_632), .Y(n_685) );
OR2x2_ASAP7_75t_L g819 ( .A(n_632), .B(n_702), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_633), .B(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g771 ( .A(n_634), .Y(n_771) );
AND2x2_ASAP7_75t_L g680 ( .A(n_635), .B(n_670), .Y(n_680) );
AND2x2_ASAP7_75t_L g716 ( .A(n_635), .B(n_637), .Y(n_716) );
AND2x2_ASAP7_75t_L g712 ( .A(n_636), .B(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_636), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g784 ( .A(n_636), .Y(n_784) );
BUFx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g655 ( .A(n_637), .Y(n_655) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_637), .Y(n_660) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_637), .Y(n_706) );
INVx1_ASAP7_75t_L g752 ( .A(n_637), .Y(n_752) );
INVx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_661), .B(n_664), .Y(n_652) );
OAI31xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .A3(n_656), .B(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g735 ( .A(n_655), .Y(n_735) );
OAI32xp33_ASAP7_75t_L g693 ( .A1(n_656), .A2(n_665), .A3(n_694), .B1(n_698), .B2(n_699), .Y(n_693) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g686 ( .A(n_662), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_671), .B1(n_674), .B2(n_678), .Y(n_664) );
OAI22xp33_ASAP7_75t_SL g749 ( .A1(n_665), .A2(n_710), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g807 ( .A(n_667), .Y(n_807) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g762 ( .A(n_670), .Y(n_762) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AND2x2_ASAP7_75t_L g688 ( .A(n_676), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g763 ( .A(n_676), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g814 ( .A(n_676), .Y(n_814) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g754 ( .A(n_680), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_687), .B2(n_688), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_683), .B(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
AND2x2_ASAP7_75t_L g740 ( .A(n_685), .B(n_701), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g745 ( .A1(n_688), .A2(n_746), .B(n_749), .C(n_753), .Y(n_745) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_690), .Y(n_803) );
INVx1_ASAP7_75t_L g820 ( .A(n_690), .Y(n_820) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_714), .C(n_727), .D(n_745), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_703), .Y(n_692) );
OR2x6_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_697), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g802 ( .A(n_700), .B(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_703) );
NOR2xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_708), .Y(n_704) );
BUFx2_ASAP7_75t_L g717 ( .A(n_705), .Y(n_717) );
AND2x4_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_711), .B(n_797), .Y(n_796) );
INVx3_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g766 ( .A(n_713), .B(n_752), .Y(n_766) );
O2A1O1Ixp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B(n_718), .C(n_719), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_716), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g776 ( .A(n_723), .B(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_739), .C(n_742), .Y(n_727) );
AND2x2_ASAP7_75t_L g806 ( .A(n_730), .B(n_807), .Y(n_806) );
NAND3xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_734), .C(n_737), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_735), .B(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_735), .B(n_771), .Y(n_801) );
INVx1_ASAP7_75t_L g744 ( .A(n_736), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_736), .Y(n_748) );
AND2x2_ASAP7_75t_L g789 ( .A(n_738), .B(n_778), .Y(n_789) );
NAND2xp33_ASAP7_75t_SL g790 ( .A(n_738), .B(n_760), .Y(n_790) );
AND2x4_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g750 ( .A(n_741), .Y(n_750) );
NOR3x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_785), .C(n_804), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_765), .C(n_775), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_763), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g778 ( .A(n_762), .Y(n_778) );
INVx2_ASAP7_75t_L g767 ( .A(n_764), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_766), .A2(n_809), .B1(n_816), .B2(n_845), .Y(n_815) );
O2A1O1Ixp5_ASAP7_75t_L g787 ( .A1(n_767), .A2(n_779), .B(n_788), .C(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AO21x1_ASAP7_75t_L g791 ( .A1(n_770), .A2(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g783 ( .A(n_774), .B(n_784), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_779), .B1(n_781), .B2(n_782), .Y(n_775) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g785 ( .A(n_786), .B(n_791), .C(n_795), .D(n_799), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .C(n_815), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVxp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x4_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
NOR2x1p5_ASAP7_75t_SL g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx6_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx10_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
CKINVDCx11_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_837), .B(n_841), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx4_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVxp33_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
CKINVDCx11_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
endmodule