module fake_netlist_1_5484_n_25 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_25);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
INVx3_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
BUFx2_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
INVxp67_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_2), .B(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_9), .B(n_11), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_9), .B(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
OAI22xp33_ASAP7_75t_L g17 ( .A1(n_13), .A2(n_10), .B1(n_8), .B2(n_12), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_14), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_18), .B(n_16), .Y(n_19) );
AOI32xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_15), .A3(n_9), .B1(n_14), .B2(n_2), .Y(n_20) );
NAND3xp33_ASAP7_75t_L g21 ( .A(n_20), .B(n_0), .C(n_1), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_3), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx2_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
endmodule