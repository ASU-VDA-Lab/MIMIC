module fake_netlist_1_4364_n_581 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_581);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_581;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_20), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_51), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_69), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_72), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_22), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_60), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_47), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_25), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_42), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_53), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_78), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_27), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_36), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_13), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_55), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_45), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_63), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_44), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_52), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_19), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_57), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_50), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_7), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_0), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_46), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_30), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_11), .B(n_58), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_43), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_1), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_5), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_16), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_68), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_2), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_0), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_86), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_121), .Y(n_124) );
NOR2xp33_ASAP7_75t_SL g125 ( .A(n_87), .B(n_34), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_121), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_99), .B(n_1), .Y(n_127) );
AND3x2_ASAP7_75t_L g128 ( .A(n_117), .B(n_2), .C(n_3), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_82), .B(n_3), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_108), .B(n_110), .Y(n_130) );
CKINVDCx6p67_ASAP7_75t_R g131 ( .A(n_88), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_110), .B(n_4), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_116), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_83), .B(n_39), .Y(n_135) );
INVx6_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_116), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_90), .B(n_8), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_111), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_130), .B(n_97), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_130), .B(n_84), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_131), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_143), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_135), .B(n_87), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
NAND2xp33_ASAP7_75t_L g164 ( .A(n_134), .B(n_109), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_134), .B(n_84), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_137), .B(n_105), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_137), .B(n_107), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_127), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_135), .B(n_107), .Y(n_173) );
OR2x6_ASAP7_75t_L g174 ( .A(n_155), .B(n_133), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_171), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_166), .B(n_141), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g177 ( .A1(n_155), .A2(n_111), .B1(n_135), .B2(n_112), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_149), .B(n_141), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_171), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
OR2x6_ASAP7_75t_L g181 ( .A(n_155), .B(n_138), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_148), .B(n_145), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
BUFx12f_ASAP7_75t_L g186 ( .A(n_163), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_162), .B(n_142), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_168), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_168), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_173), .A2(n_132), .B1(n_112), .B2(n_119), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_168), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_169), .B(n_142), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_163), .B(n_125), .Y(n_193) );
NAND2xp33_ASAP7_75t_L g194 ( .A(n_170), .B(n_95), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_172), .B(n_129), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_168), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_164), .A2(n_119), .B1(n_139), .B2(n_122), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_167), .B(n_126), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_156), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_157), .A2(n_106), .B(n_115), .Y(n_207) );
BUFx4f_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
OR2x6_ASAP7_75t_L g210 ( .A(n_186), .B(n_114), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_195), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_182), .B(n_128), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_182), .A2(n_100), .B(n_126), .C(n_124), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_195), .B(n_124), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_197), .B(n_124), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_177), .A2(n_124), .B1(n_93), .B2(n_120), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_186), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_198), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_180), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_175), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_180), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_184), .B(n_109), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_192), .B(n_98), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g228 ( .A1(n_174), .A2(n_98), .B1(n_95), .B2(n_118), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_174), .A2(n_102), .B1(n_104), .B2(n_96), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_203), .A2(n_103), .B(n_113), .C(n_101), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_178), .A2(n_88), .B1(n_106), .B2(n_115), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_178), .B(n_9), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_174), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_201), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_181), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_189), .B(n_86), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_184), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_204), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_187), .A2(n_150), .B(n_151), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_176), .B(n_123), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_189), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_184), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_225), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_237), .Y(n_247) );
OAI21x1_ASAP7_75t_SL g248 ( .A1(n_245), .A2(n_207), .B(n_191), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_217), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_221), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_234), .B(n_188), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_233), .A2(n_187), .B(n_179), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_230), .A2(n_193), .B(n_223), .C(n_235), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_216), .A2(n_181), .B1(n_190), .B2(n_194), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_242), .A2(n_193), .B(n_179), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_242), .A2(n_183), .B(n_185), .Y(n_256) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_243), .A2(n_123), .B(n_203), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_213), .A2(n_188), .B(n_151), .Y(n_258) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_202), .B(n_196), .Y(n_259) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_240), .A2(n_150), .B(n_153), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_216), .A2(n_181), .B1(n_194), .B2(n_206), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_227), .B(n_206), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_219), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_241), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_221), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_212), .B(n_209), .Y(n_267) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_229), .A2(n_153), .B(n_150), .Y(n_268) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_219), .Y(n_269) );
OAI22x1_ASAP7_75t_L g270 ( .A1(n_236), .A2(n_209), .B1(n_206), .B2(n_205), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_244), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_238), .A2(n_153), .B(n_151), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
AO32x2_ASAP7_75t_L g274 ( .A1(n_228), .A2(n_209), .A3(n_208), .B1(n_136), .B2(n_146), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_220), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_255), .A2(n_238), .B(n_226), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_254), .A2(n_232), .B1(n_214), .B2(n_212), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_246), .Y(n_279) );
OAI21xp33_ASAP7_75t_L g280 ( .A1(n_262), .A2(n_227), .B(n_231), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_249), .Y(n_281) );
INVx4_ASAP7_75t_L g282 ( .A(n_275), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_249), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_211), .B1(n_214), .B2(n_215), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_211), .B1(n_220), .B2(n_224), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_250), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_239), .B(n_222), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_249), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_266), .B(n_245), .Y(n_290) );
OAI211xp5_ASAP7_75t_L g291 ( .A1(n_266), .A2(n_218), .B(n_210), .C(n_159), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_259), .B(n_224), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_259), .B(n_224), .Y(n_293) );
AO21x1_ASAP7_75t_L g294 ( .A1(n_258), .A2(n_146), .B(n_237), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
AOI222xp33_ASAP7_75t_L g297 ( .A1(n_267), .A2(n_237), .B1(n_208), .B2(n_210), .C1(n_12), .C2(n_13), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_259), .A2(n_210), .B1(n_237), .B2(n_146), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_253), .A2(n_160), .B(n_152), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_265), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_283), .B(n_273), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_282), .Y(n_303) );
AO31x2_ASAP7_75t_L g304 ( .A1(n_294), .A2(n_270), .A3(n_271), .B(n_263), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_283), .B(n_271), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_281), .B(n_257), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_281), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_289), .B(n_257), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_286), .B(n_259), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_289), .Y(n_314) );
AO31x2_ASAP7_75t_L g315 ( .A1(n_294), .A2(n_270), .A3(n_263), .B(n_264), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_279), .B(n_257), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_282), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_288), .B(n_257), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_279), .B(n_252), .Y(n_321) );
AOI31xp33_ASAP7_75t_L g322 ( .A1(n_297), .A2(n_269), .A3(n_274), .B(n_252), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_278), .A2(n_251), .B1(n_248), .B2(n_270), .C(n_268), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_295), .B(n_274), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_306), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_318), .B(n_292), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_318), .B(n_293), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g328 ( .A(n_312), .B(n_297), .C(n_298), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_303), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_310), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_324), .B(n_293), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_324), .B(n_295), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_310), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_324), .B(n_300), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_320), .B(n_290), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_317), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_307), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_321), .B(n_300), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
OAI33xp33_ASAP7_75t_L g345 ( .A1(n_320), .A2(n_284), .A3(n_290), .B1(n_285), .B2(n_280), .B3(n_14), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_303), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_311), .B(n_287), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_316), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_303), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_323), .A2(n_280), .B1(n_251), .B2(n_268), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_302), .B(n_287), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_302), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_302), .B(n_287), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_303), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_333), .B(n_304), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_353), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_355), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_338), .B(n_313), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_338), .B(n_313), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_341), .B(n_313), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_325), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_333), .B(n_304), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_347), .B(n_304), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_347), .B(n_304), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_334), .B(n_305), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_341), .B(n_304), .Y(n_368) );
OR2x6_ASAP7_75t_L g369 ( .A(n_336), .B(n_308), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_343), .B(n_304), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_343), .B(n_304), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_330), .B(n_322), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_353), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_344), .B(n_326), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_344), .B(n_314), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_326), .B(n_314), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_327), .B(n_315), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_334), .B(n_305), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_329), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_329), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_331), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_331), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_327), .B(n_314), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_337), .B(n_339), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_337), .B(n_315), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_339), .B(n_315), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_342), .B(n_321), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_342), .B(n_322), .Y(n_392) );
AND3x2_ASAP7_75t_L g393 ( .A(n_336), .B(n_247), .C(n_323), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_340), .B(n_315), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_346), .B(n_291), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g396 ( .A1(n_328), .A2(n_319), .B(n_308), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_335), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_340), .B(n_315), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
BUFx12f_ASAP7_75t_L g400 ( .A(n_355), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_360), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_388), .B(n_352), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_352), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_396), .B(n_349), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_377), .B(n_349), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_356), .B(n_354), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_364), .B(n_354), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_377), .B(n_332), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_364), .B(n_351), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_388), .B(n_328), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_357), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_387), .B(n_332), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_400), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_372), .A2(n_345), .B1(n_350), .B2(n_301), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_365), .B(n_351), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_395), .B(n_345), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_365), .B(n_351), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_375), .B(n_351), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_375), .B(n_308), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_400), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_387), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_389), .B(n_308), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_392), .B(n_319), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_366), .B(n_389), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_367), .B(n_319), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_380), .B(n_319), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_391), .B(n_316), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_359), .B(n_316), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_366), .B(n_315), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_386), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_378), .B(n_315), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_359), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_383), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_378), .B(n_301), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_361), .B(n_301), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_361), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_386), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_369), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_368), .B(n_301), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_383), .B(n_9), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_362), .B(n_287), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_373), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_368), .B(n_268), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_370), .B(n_268), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_394), .B(n_10), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_369), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_362), .B(n_285), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g453 ( .A(n_396), .B(n_251), .C(n_299), .D(n_12), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_369), .Y(n_454) );
AOI321xp33_ASAP7_75t_L g455 ( .A1(n_418), .A2(n_371), .A3(n_370), .B1(n_394), .B2(n_398), .C(n_385), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_412), .B(n_398), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_401), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_453), .A2(n_369), .B(n_370), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_415), .A2(n_369), .B1(n_374), .B2(n_358), .Y(n_459) );
AOI211xp5_ASAP7_75t_L g460 ( .A1(n_418), .A2(n_370), .B(n_371), .C(n_390), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_407), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_404), .A2(n_374), .B(n_358), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_426), .B(n_371), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_422), .B(n_384), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_450), .A2(n_390), .B(n_385), .C(n_384), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_416), .A2(n_445), .B(n_422), .Y(n_467) );
NAND3xp33_ASAP7_75t_SL g468 ( .A(n_416), .B(n_247), .C(n_376), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_425), .A2(n_371), .B1(n_393), .B2(n_358), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_409), .B(n_414), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_443), .A2(n_358), .B1(n_374), .B2(n_376), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_432), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_445), .A2(n_374), .B(n_399), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_426), .B(n_399), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_454), .B(n_397), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_437), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_413), .A2(n_146), .B1(n_381), .B2(n_379), .C(n_382), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_403), .B(n_382), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_436), .Y(n_482) );
NOR2xp67_ASAP7_75t_SL g483 ( .A(n_404), .B(n_282), .Y(n_483) );
AOI211xp5_ASAP7_75t_SL g484 ( .A1(n_427), .A2(n_381), .B(n_379), .C(n_269), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g486 ( .A1(n_451), .A2(n_10), .B(n_11), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_435), .A2(n_258), .B(n_251), .C(n_276), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_421), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_435), .A2(n_146), .B(n_276), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_428), .A2(n_296), .B1(n_273), .B2(n_264), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_423), .B(n_146), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_440), .A2(n_255), .B(n_251), .Y(n_492) );
AOI21xp33_ASAP7_75t_L g493 ( .A1(n_446), .A2(n_14), .B(n_15), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_403), .B(n_296), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_433), .B(n_255), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_424), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_433), .B(n_256), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_402), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_406), .B(n_260), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_410), .A2(n_248), .B1(n_152), .B2(n_160), .C(n_147), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_439), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_482), .B(n_408), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_485), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_482), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_471), .A2(n_410), .B1(n_417), .B2(n_419), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_455), .B(n_419), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_467), .A2(n_452), .B1(n_405), .B2(n_448), .C(n_444), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_455), .A2(n_417), .B(n_438), .C(n_408), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_488), .Y(n_510) );
AND2x2_ASAP7_75t_SL g511 ( .A(n_469), .B(n_406), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_460), .A2(n_429), .B1(n_431), .B2(n_449), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_468), .A2(n_449), .B(n_442), .C(n_441), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_476), .B(n_441), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_457), .Y(n_515) );
AOI211xp5_ASAP7_75t_L g516 ( .A1(n_459), .A2(n_442), .B(n_434), .C(n_274), .Y(n_516) );
OAI22xp33_ASAP7_75t_SL g517 ( .A1(n_470), .A2(n_274), .B1(n_273), .B2(n_264), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_464), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_480), .B(n_496), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_502), .Y(n_520) );
AO22x1_ASAP7_75t_L g521 ( .A1(n_458), .A2(n_274), .B1(n_263), .B2(n_275), .Y(n_521) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_484), .B(n_17), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_486), .A2(n_274), .B(n_260), .C(n_23), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_494), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_461), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_465), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_474), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_478), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_463), .B(n_274), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_498), .B(n_260), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_484), .A2(n_256), .B(n_272), .C(n_275), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_456), .B(n_260), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_472), .B(n_18), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_475), .A2(n_275), .B1(n_260), .B2(n_256), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_515), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_508), .A2(n_466), .B1(n_493), .B2(n_481), .C(n_473), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_508), .A2(n_462), .B1(n_477), .B2(n_497), .C(n_479), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_507), .A2(n_491), .B(n_489), .Y(n_538) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_511), .B(n_500), .Y(n_539) );
NOR4xp25_ASAP7_75t_L g540 ( .A(n_505), .B(n_501), .C(n_487), .D(n_499), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_525), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_512), .A2(n_477), .B1(n_492), .B2(n_495), .C(n_483), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_513), .A2(n_490), .B(n_272), .C(n_275), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_509), .A2(n_275), .B1(n_160), .B2(n_152), .C(n_147), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_510), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g546 ( .A1(n_516), .A2(n_272), .B(n_160), .C(n_152), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_503), .Y(n_547) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_506), .A2(n_160), .B1(n_152), .B2(n_147), .C(n_29), .Y(n_548) );
AOI21xp33_ASAP7_75t_L g549 ( .A1(n_533), .A2(n_21), .B(n_26), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_524), .B(n_28), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_531), .A2(n_32), .B(n_33), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_522), .A2(n_147), .B(n_38), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_535), .Y(n_554) );
OAI211xp5_ASAP7_75t_SL g555 ( .A1(n_536), .A2(n_518), .B(n_520), .C(n_523), .Y(n_555) );
AOI211xp5_ASAP7_75t_L g556 ( .A1(n_540), .A2(n_521), .B(n_517), .C(n_523), .Y(n_556) );
AOI211xp5_ASAP7_75t_L g557 ( .A1(n_540), .A2(n_529), .B(n_504), .C(n_532), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g558 ( .A1(n_542), .A2(n_527), .B1(n_528), .B2(n_519), .C1(n_532), .C2(n_530), .Y(n_558) );
OAI321xp33_ASAP7_75t_L g559 ( .A1(n_544), .A2(n_530), .A3(n_514), .B1(n_534), .B2(n_147), .C(n_54), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_541), .Y(n_560) );
AOI211xp5_ASAP7_75t_L g561 ( .A1(n_538), .A2(n_37), .B(n_40), .C(n_41), .Y(n_561) );
AOI211xp5_ASAP7_75t_L g562 ( .A1(n_552), .A2(n_49), .B(n_56), .C(n_59), .Y(n_562) );
OA22x2_ASAP7_75t_SL g563 ( .A1(n_539), .A2(n_61), .B1(n_62), .B2(n_64), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_550), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_560), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_555), .B(n_543), .C(n_546), .Y(n_566) );
NOR2x1p5_ASAP7_75t_L g567 ( .A(n_564), .B(n_547), .Y(n_567) );
NAND4xp75_ASAP7_75t_L g568 ( .A(n_563), .B(n_537), .C(n_551), .D(n_549), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_556), .A2(n_545), .B(n_548), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_558), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_565), .Y(n_571) );
NAND5xp2_ASAP7_75t_L g572 ( .A(n_569), .B(n_557), .C(n_562), .D(n_561), .E(n_559), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_570), .A2(n_554), .B1(n_553), .B2(n_67), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_571), .Y(n_574) );
OA22x2_ASAP7_75t_L g575 ( .A1(n_572), .A2(n_567), .B1(n_568), .B2(n_566), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g576 ( .A1(n_575), .A2(n_573), .B1(n_66), .B2(n_73), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_574), .A2(n_65), .B(n_74), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_576), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_578), .A2(n_577), .B1(n_76), .B2(n_77), .Y(n_579) );
XOR2xp5_ASAP7_75t_L g580 ( .A(n_579), .B(n_75), .Y(n_580) );
AOI22xp5_ASAP7_75t_SL g581 ( .A1(n_580), .A2(n_81), .B1(n_79), .B2(n_80), .Y(n_581) );
endmodule