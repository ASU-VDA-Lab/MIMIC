module fake_jpeg_2569_n_648 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_576;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_59),
.B(n_60),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_24),
.B(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_79),
.Y(n_132)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_72),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_73),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_76),
.B(n_91),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_8),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_80),
.Y(n_201)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_90),
.Y(n_149)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_29),
.Y(n_89)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_23),
.B(n_8),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_37),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_103),
.Y(n_150)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_7),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_105),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_41),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_113),
.B(n_126),
.Y(n_187)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_45),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_116),
.B(n_18),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_45),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_45),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_122),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_123),
.Y(n_211)
);

BUFx4f_ASAP7_75t_SL g124 ( 
.A(n_48),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g127 ( 
.A(n_48),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_28),
.B(n_7),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_28),
.Y(n_130)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_131),
.A2(n_41),
.B(n_50),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_29),
.B1(n_51),
.B2(n_55),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_135),
.A2(n_140),
.B1(n_146),
.B2(n_147),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_51),
.C(n_58),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_137),
.B(n_181),
.C(n_66),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_34),
.B1(n_57),
.B2(n_56),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_138),
.A2(n_173),
.B1(n_191),
.B2(n_110),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_62),
.A2(n_34),
.B1(n_57),
.B2(n_56),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_74),
.A2(n_29),
.B1(n_51),
.B2(n_55),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_36),
.B1(n_29),
.B2(n_58),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_74),
.A2(n_32),
.B1(n_49),
.B2(n_39),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_148),
.A2(n_159),
.B1(n_170),
.B2(n_197),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_72),
.A2(n_36),
.B1(n_40),
.B2(n_49),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_40),
.B1(n_55),
.B2(n_33),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_217),
.C(n_15),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_83),
.A2(n_39),
.B1(n_49),
.B2(n_33),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_39),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_178),
.B(n_184),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_114),
.A2(n_38),
.B1(n_33),
.B2(n_35),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_179),
.A2(n_148),
.B(n_212),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_64),
.A2(n_38),
.B(n_35),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_124),
.B(n_38),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_86),
.B(n_35),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_185),
.B(n_199),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_92),
.A2(n_32),
.B1(n_50),
.B2(n_45),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_0),
.B(n_3),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_73),
.A2(n_118),
.B1(n_125),
.B2(n_96),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_94),
.A2(n_97),
.B1(n_106),
.B2(n_104),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_214),
.B1(n_222),
.B2(n_110),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_108),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_73),
.A2(n_32),
.B1(n_50),
.B2(n_45),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_225),
.B1(n_139),
.B2(n_201),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_99),
.A2(n_44),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_86),
.B(n_44),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_67),
.B(n_44),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_127),
.B(n_10),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_218),
.B(n_221),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_71),
.B(n_10),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_75),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_105),
.A2(n_80),
.B1(n_66),
.B2(n_131),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_80),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_227),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_68),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_228),
.B(n_243),
.Y(n_328)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_229),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_151),
.B(n_0),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_230),
.B(n_267),
.Y(n_341)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_231),
.Y(n_348)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_232),
.Y(n_347)
);

BUFx4f_ASAP7_75t_SL g233 ( 
.A(n_174),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_233),
.Y(n_344)
);

OA22x2_ASAP7_75t_L g312 ( 
.A1(n_235),
.A2(n_240),
.B1(n_280),
.B2(n_197),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_237),
.Y(n_334)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_238),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_239),
.B(n_258),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_145),
.A2(n_131),
.B1(n_3),
.B2(n_5),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_241),
.A2(n_252),
.B1(n_261),
.B2(n_272),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_242),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_132),
.B(n_5),
.Y(n_244)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_244),
.Y(n_321)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_245),
.Y(n_359)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_139),
.Y(n_248)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_150),
.A2(n_5),
.B1(n_11),
.B2(n_13),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_168),
.A2(n_171),
.B1(n_217),
.B2(n_158),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_253),
.B(n_275),
.Y(n_339)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_254),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_201),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_156),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_262),
.Y(n_315)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_134),
.Y(n_257)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_162),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_259),
.Y(n_369)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_141),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_260),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_137),
.A2(n_16),
.B1(n_18),
.B2(n_176),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_263),
.A2(n_264),
.B1(n_307),
.B2(n_309),
.Y(n_317)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_149),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_277),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_160),
.B(n_16),
.Y(n_267)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_269),
.Y(n_353)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_270),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_190),
.B(n_216),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_282),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_142),
.A2(n_181),
.B1(n_165),
.B2(n_195),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_192),
.B(n_203),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_273),
.B(n_276),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_146),
.A2(n_135),
.B(n_225),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_274),
.A2(n_243),
.B(n_246),
.C(n_262),
.Y(n_330)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_166),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_155),
.B(n_224),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_167),
.B(n_195),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_177),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_281),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_165),
.A2(n_186),
.B1(n_223),
.B2(n_219),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_213),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_287),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_193),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_286),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_169),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_285),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_163),
.B(n_143),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_188),
.B(n_206),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_289),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_163),
.B(n_206),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_294),
.Y(n_357)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_292),
.B(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_169),
.B(n_177),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_186),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_295),
.B(n_300),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_226),
.B(n_179),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_301),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_133),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_204),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_299),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_152),
.B(n_175),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_166),
.B(n_194),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_161),
.B(n_220),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_304),
.Y(n_367)
);

OR2x2_ASAP7_75t_SL g303 ( 
.A(n_161),
.B(n_220),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_189),
.C(n_144),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_152),
.B(n_175),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_133),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_305),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_180),
.B(n_200),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_305),
.Y(n_361)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_164),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_180),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_308),
.Y(n_365)
);

INVx4_ASAP7_75t_SL g309 ( 
.A(n_211),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_194),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_310),
.A2(n_248),
.B1(n_309),
.B2(n_290),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_269),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_223),
.B1(n_164),
.B2(n_219),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_313),
.A2(n_310),
.B1(n_308),
.B2(n_297),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_296),
.A2(n_200),
.B1(n_189),
.B2(n_204),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_316),
.A2(n_322),
.B1(n_332),
.B2(n_242),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_L g384 ( 
.A1(n_320),
.A2(n_351),
.B(n_275),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_235),
.A2(n_144),
.B1(n_202),
.B2(n_283),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_258),
.A2(n_202),
.B(n_254),
.C(n_281),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_324),
.A2(n_350),
.B(n_320),
.C(n_334),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_230),
.B(n_228),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_325),
.B(n_345),
.C(n_284),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_330),
.A2(n_278),
.B(n_291),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_240),
.A2(n_246),
.B1(n_234),
.B2(n_274),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_271),
.B(n_246),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_340),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_265),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_279),
.A2(n_303),
.B1(n_249),
.B2(n_247),
.Y(n_351)
);

AOI22x1_ASAP7_75t_L g360 ( 
.A1(n_301),
.A2(n_306),
.B1(n_267),
.B2(n_251),
.Y(n_360)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_366),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_268),
.B(n_298),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_371),
.A2(n_374),
.B1(n_381),
.B2(n_384),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_337),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_372),
.B(n_383),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_356),
.A2(n_261),
.B1(n_252),
.B2(n_259),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_325),
.B(n_236),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_402),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_324),
.A2(n_292),
.B(n_287),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_376),
.A2(n_389),
.B(n_413),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_260),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_380),
.Y(n_423)
);

OAI22x1_ASAP7_75t_L g451 ( 
.A1(n_378),
.A2(n_347),
.B1(n_368),
.B2(n_359),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_366),
.B(n_250),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_379),
.B(n_387),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_257),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_229),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_386),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_321),
.C(n_315),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_355),
.A2(n_232),
.B(n_248),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_293),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_318),
.A2(n_231),
.B1(n_245),
.B2(n_307),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_395),
.A2(n_314),
.B1(n_329),
.B2(n_336),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_233),
.B(n_270),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_396),
.A2(n_417),
.B(n_317),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_284),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_403),
.C(n_328),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_346),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_407),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_333),
.B(n_233),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_400),
.B(n_401),
.Y(n_424)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_328),
.B(n_238),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_264),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_404),
.B(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_333),
.B(n_341),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_406),
.B(n_411),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_318),
.B(n_360),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_369),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_412),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_322),
.A2(n_332),
.B1(n_330),
.B2(n_343),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_340),
.B1(n_343),
.B2(n_312),
.Y(n_431)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_410),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_341),
.B(n_363),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_361),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_355),
.A2(n_350),
.B(n_339),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_345),
.B(n_367),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_414),
.B(n_416),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_323),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_319),
.Y(n_443)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_339),
.B(n_357),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_418),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_378),
.A2(n_334),
.B1(n_339),
.B2(n_354),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_425),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_403),
.Y(n_463)
);

OAI32xp33_ASAP7_75t_L g430 ( 
.A1(n_407),
.A2(n_340),
.A3(n_316),
.B1(n_354),
.B2(n_313),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_431),
.A2(n_437),
.B1(n_444),
.B2(n_450),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_412),
.A2(n_342),
.B(n_340),
.C(n_312),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_432),
.B(n_439),
.Y(n_477)
);

OAI21xp33_ASAP7_75t_SL g469 ( 
.A1(n_434),
.A2(n_435),
.B(n_438),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_385),
.A2(n_311),
.B1(n_327),
.B2(n_364),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_409),
.A2(n_312),
.B1(n_327),
.B2(n_364),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_385),
.A2(n_311),
.B1(n_358),
.B2(n_319),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_375),
.B(n_402),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_445),
.C(n_427),
.Y(n_468)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_392),
.A2(n_358),
.B1(n_365),
.B2(n_352),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_352),
.C(n_370),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_392),
.A2(n_365),
.B1(n_314),
.B2(n_329),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_452),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_451),
.A2(n_386),
.B1(n_395),
.B2(n_371),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_373),
.B(n_399),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_344),
.B(n_370),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_454),
.A2(n_455),
.B(n_396),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_389),
.A2(n_344),
.B(n_347),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_378),
.A2(n_336),
.B1(n_348),
.B2(n_359),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_415),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_455),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_461),
.B(n_471),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_420),
.C(n_414),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_462),
.B(n_472),
.C(n_476),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_463),
.B(n_464),
.C(n_468),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_426),
.B(n_373),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_426),
.B(n_398),
.C(n_401),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_470),
.B(n_482),
.C(n_488),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_443),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_408),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_436),
.Y(n_474)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_475),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_424),
.B(n_377),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_477),
.B(n_430),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_419),
.A2(n_376),
.B(n_417),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_487),
.B(n_419),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_440),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_481),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_445),
.C(n_457),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_439),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_483),
.B(n_486),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_457),
.B(n_380),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_484),
.B(n_441),
.Y(n_502)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_382),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_381),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_429),
.B(n_458),
.Y(n_489)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_440),
.B(n_416),
.Y(n_490)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_491),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_424),
.Y(n_492)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_444),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_423),
.Y(n_524)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_421),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_495),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_432),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_499),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_441),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_502),
.B(n_530),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_460),
.A2(n_422),
.B1(n_434),
.B2(n_428),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_507),
.A2(n_469),
.B1(n_478),
.B2(n_473),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_431),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_528),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_513),
.A2(n_487),
.B(n_473),
.Y(n_550)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_467),
.Y(n_514)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_514),
.Y(n_535)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_516),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_459),
.A2(n_437),
.B1(n_422),
.B2(n_428),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_517),
.A2(n_526),
.B1(n_494),
.B2(n_471),
.Y(n_541)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_475),
.Y(n_518)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_518),
.Y(n_548)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_523),
.Y(n_532)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_465),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_524),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_460),
.A2(n_447),
.B1(n_451),
.B2(n_374),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_468),
.B(n_425),
.C(n_391),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_488),
.C(n_484),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_386),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_483),
.B(n_453),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_466),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_533),
.B(n_542),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_506),
.B(n_480),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_534),
.B(n_543),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_536),
.A2(n_544),
.B1(n_551),
.B2(n_519),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_498),
.B(n_465),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_538),
.B(n_503),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_539),
.B(n_509),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_541),
.A2(n_556),
.B1(n_526),
.B2(n_511),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_481),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_501),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_515),
.A2(n_461),
.B1(n_466),
.B2(n_491),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_476),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_545),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_505),
.B(n_525),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_546),
.Y(n_576)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_547),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_550),
.A2(n_509),
.B(n_513),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_515),
.A2(n_486),
.B1(n_479),
.B2(n_451),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_508),
.B(n_493),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_552),
.B(n_555),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_410),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_553),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_520),
.B(n_527),
.C(n_528),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_520),
.C(n_502),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_517),
.A2(n_456),
.B1(n_453),
.B2(n_495),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_501),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_558),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_499),
.B(n_449),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_529),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_522),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_510),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_561),
.B(n_572),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_562),
.B(n_564),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_563),
.B(n_581),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_524),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_565),
.B(n_566),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_567),
.Y(n_584)
);

A2O1A1O1Ixp25_ASAP7_75t_L g568 ( 
.A1(n_554),
.A2(n_522),
.B(n_507),
.C(n_519),
.D(n_504),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_568),
.A2(n_574),
.B(n_548),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_569),
.A2(n_541),
.B1(n_554),
.B2(n_556),
.Y(n_585)
);

XNOR2x1_ASAP7_75t_L g596 ( 
.A(n_570),
.B(n_535),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_500),
.Y(n_574)
);

CKINVDCx11_ASAP7_75t_R g578 ( 
.A(n_532),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_578),
.B(n_393),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_540),
.B(n_496),
.C(n_449),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_580),
.B(n_538),
.C(n_533),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_550),
.A2(n_415),
.B(n_405),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_582),
.B(n_598),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_585),
.B(n_594),
.Y(n_601)
);

AOI211xp5_ASAP7_75t_L g586 ( 
.A1(n_569),
.A2(n_544),
.B(n_536),
.C(n_551),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_586),
.A2(n_583),
.B1(n_564),
.B2(n_598),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_571),
.B(n_552),
.C(n_540),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_592),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_537),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_593),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_566),
.B(n_537),
.C(n_531),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_531),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_561),
.B(n_548),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_570),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_SL g608 ( 
.A(n_595),
.B(n_596),
.Y(n_608)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_597),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_563),
.B(n_549),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_573),
.A2(n_549),
.B(n_535),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_599),
.A2(n_576),
.B(n_560),
.Y(n_604)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_600),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_602),
.A2(n_586),
.B1(n_585),
.B2(n_595),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_604),
.A2(n_605),
.B(n_596),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_590),
.A2(n_575),
.B(n_565),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_584),
.B(n_587),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_607),
.B(n_609),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_591),
.C(n_594),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_588),
.B(n_581),
.C(n_579),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_610),
.B(n_612),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_600),
.B(n_577),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_562),
.C(n_575),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_615),
.C(n_394),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_568),
.C(n_578),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_617),
.A2(n_620),
.B1(n_622),
.B2(n_616),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_SL g634 ( 
.A(n_618),
.B(n_608),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_603),
.B(n_592),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_619),
.B(n_626),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_606),
.A2(n_614),
.B1(n_615),
.B2(n_601),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_609),
.B(n_593),
.Y(n_621)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_621),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_601),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_610),
.B(n_421),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_624),
.B(n_625),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_613),
.B(n_421),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_605),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_628),
.B(n_446),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_623),
.B(n_611),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_632),
.B(n_633),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_634),
.A2(n_388),
.B(n_390),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_SL g639 ( 
.A1(n_635),
.A2(n_624),
.B(n_617),
.C(n_625),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_446),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_636),
.B(n_621),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_630),
.B(n_627),
.C(n_626),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_638),
.B(n_639),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_640),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_641),
.B(n_631),
.C(n_629),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_637),
.C(n_634),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_642),
.B(n_643),
.Y(n_646)
);

AOI221xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_629),
.B1(n_446),
.B2(n_348),
.C(n_362),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_362),
.Y(n_648)
);


endmodule