module fake_jpeg_6494_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_26),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_21),
.B(n_14),
.C(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_24),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_15),
.B1(n_35),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_53),
.B1(n_24),
.B2(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_15),
.B1(n_16),
.B2(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_66),
.B1(n_53),
.B2(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_41),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_43),
.B1(n_26),
.B2(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_0),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_69),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_39),
.B(n_44),
.C(n_47),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_78),
.B(n_83),
.C(n_60),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_57),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_84),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_85),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_41),
.B(n_45),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_17),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_63),
.B(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_102),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_91),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_99),
.B1(n_86),
.B2(n_87),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_65),
.C(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_69),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_64),
.B1(n_69),
.B2(n_51),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_87),
.B1(n_81),
.B2(n_86),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_66),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_57),
.B1(n_60),
.B2(n_51),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_48),
.B1(n_29),
.B2(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_51),
.B1(n_48),
.B2(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_14),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_14),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_13),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_133),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_103),
.C(n_97),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_128),
.C(n_132),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_91),
.C(n_48),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_0),
.C(n_1),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_12),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_116),
.C(n_104),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_104),
.C(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_111),
.C(n_110),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_115),
.B(n_105),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_140),
.B1(n_109),
.B2(n_139),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_107),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_130),
.B(n_121),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_154),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_122),
.B(n_131),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_150),
.B(n_151),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_R g152 ( 
.A1(n_137),
.A2(n_11),
.B(n_10),
.C(n_3),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_138),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_153),
.A2(n_134),
.B1(n_10),
.B2(n_4),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_136),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_158),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_147),
.B(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_2),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_3),
.B(n_4),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_6),
.B1(n_8),
.B2(n_155),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_6),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.C(n_8),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_163),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.C(n_172),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_164),
.C(n_167),
.Y(n_176)
);


endmodule