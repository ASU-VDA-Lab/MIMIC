module real_aes_18180_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g889 ( .A(n_0), .B(n_890), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_1), .A2(n_516), .B1(n_517), .B2(n_519), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_1), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_2), .A2(n_36), .B1(n_143), .B2(n_235), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_3), .A2(n_12), .B1(n_548), .B2(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g890 ( .A(n_4), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_5), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_6), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_7), .A2(n_13), .B1(n_549), .B2(n_585), .Y(n_584) );
XNOR2xp5_ASAP7_75t_L g517 ( .A(n_8), .B(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g122 ( .A(n_9), .B(n_32), .Y(n_122) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_10), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_11), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_14), .B(n_158), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_15), .A2(n_102), .B1(n_188), .B2(n_548), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_16), .A2(n_33), .B1(n_566), .B2(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_17), .B(n_158), .Y(n_563) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_18), .A2(n_49), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_19), .B(n_239), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_20), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_20), .A2(n_95), .B1(n_621), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_21), .A2(n_40), .B1(n_195), .B2(n_210), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_22), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_23), .A2(n_46), .B1(n_210), .B2(n_548), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_24), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_25), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_26), .B(n_218), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_27), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_28), .Y(n_892) );
XNOR2x1_ASAP7_75t_L g518 ( .A(n_29), .B(n_41), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_30), .B(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_31), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_34), .A2(n_86), .B1(n_143), .B2(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_35), .A2(n_39), .B1(n_143), .B2(n_551), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_37), .A2(n_52), .B1(n_548), .B2(n_603), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_38), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_42), .B(n_158), .Y(n_206) );
INVx2_ASAP7_75t_L g117 ( .A(n_43), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_44), .B(n_191), .Y(n_233) );
BUFx3_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
INVx1_ASAP7_75t_L g871 ( .A(n_45), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_47), .B(n_177), .Y(n_241) );
XOR2x2_ASAP7_75t_L g125 ( .A(n_48), .B(n_126), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_48), .A2(n_859), .B1(n_860), .B2(n_863), .Y(n_858) );
INVx1_ASAP7_75t_L g863 ( .A(n_48), .Y(n_863) );
AND2x2_ASAP7_75t_L g269 ( .A(n_50), .B(n_177), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_51), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_53), .B(n_218), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_54), .B(n_195), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_55), .A2(n_73), .B1(n_195), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_56), .A2(n_76), .B1(n_143), .B2(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_57), .B(n_299), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_58), .A2(n_147), .B(n_156), .C(n_262), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_59), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_60), .A2(n_99), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
AND2x4_ASAP7_75t_L g161 ( .A(n_62), .B(n_162), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_63), .A2(n_64), .B1(n_210), .B2(n_222), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_65), .A2(n_83), .B1(n_861), .B2(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_65), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_66), .B(n_136), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_67), .B(n_177), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_68), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_69), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g162 ( .A(n_70), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_71), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_72), .B(n_136), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_74), .B(n_143), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_75), .B(n_191), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_77), .B(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g149 ( .A(n_78), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_79), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_80), .B(n_158), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_81), .B(n_152), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_82), .A2(n_98), .B1(n_156), .B2(n_210), .Y(n_535) );
INVx1_ASAP7_75t_L g862 ( .A(n_83), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_84), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_85), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_87), .A2(n_92), .B1(n_217), .B2(n_218), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_88), .B(n_158), .Y(n_190) );
NAND2xp33_ASAP7_75t_SL g175 ( .A(n_89), .B(n_146), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_90), .B(n_189), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_91), .B(n_136), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_93), .Y(n_588) );
INVx1_ASAP7_75t_L g113 ( .A(n_94), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_94), .B(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g857 ( .A(n_95), .Y(n_857) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_96), .B(n_158), .Y(n_567) );
NAND2xp33_ASAP7_75t_L g145 ( .A(n_97), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_100), .B(n_177), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g171 ( .A(n_101), .B(n_146), .C(n_170), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_103), .B(n_143), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_104), .B(n_218), .Y(n_297) );
AOI21xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_882), .B(n_891), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_872), .Y(n_106) );
OAI211xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_123), .B(n_520), .C(n_849), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2xp67_ASAP7_75t_SL g109 ( .A(n_110), .B(n_114), .Y(n_109) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g842 ( .A(n_112), .B(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g848 ( .A(n_113), .Y(n_848) );
NOR2x1_ASAP7_75t_R g846 ( .A(n_114), .B(n_847), .Y(n_846) );
INVx5_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x6_ASAP7_75t_SL g115 ( .A(n_116), .B(n_118), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_117), .B(n_841), .Y(n_840) );
INVx3_ASAP7_75t_L g852 ( .A(n_117), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_120), .B(n_122), .Y(n_843) );
AND3x2_ASAP7_75t_L g869 ( .A(n_121), .B(n_848), .C(n_870), .Y(n_869) );
AND2x6_ASAP7_75t_SL g874 ( .A(n_121), .B(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g886 ( .A(n_122), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_514), .B2(n_515), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_126), .Y(n_866) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_446), .Y(n_126) );
NAND4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_321), .C(n_361), .D(n_410), .Y(n_127) );
NOR2xp67_ASAP7_75t_L g128 ( .A(n_129), .B(n_270), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_180), .B1(n_242), .B2(n_251), .Y(n_129) );
INVx1_ASAP7_75t_L g442 ( .A(n_130), .Y(n_442) );
INVx1_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_131), .B(n_289), .Y(n_358) );
AND2x2_ASAP7_75t_L g389 ( .A(n_131), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_163), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_132), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g313 ( .A(n_132), .Y(n_313) );
AND2x2_ASAP7_75t_L g488 ( .A(n_132), .B(n_356), .Y(n_488) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx2_ASAP7_75t_L g253 ( .A(n_133), .Y(n_253) );
AND2x2_ASAP7_75t_L g341 ( .A(n_133), .B(n_303), .Y(n_341) );
AND2x2_ASAP7_75t_L g385 ( .A(n_133), .B(n_290), .Y(n_385) );
OR2x2_ASAP7_75t_L g403 ( .A(n_133), .B(n_404), .Y(n_403) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g307 ( .A(n_134), .B(n_290), .Y(n_307) );
BUFx2_ASAP7_75t_L g364 ( .A(n_134), .Y(n_364) );
OR2x2_ASAP7_75t_L g372 ( .A(n_134), .B(n_330), .Y(n_372) );
INVx1_ASAP7_75t_L g427 ( .A(n_134), .Y(n_427) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
INVx2_ASAP7_75t_L g575 ( .A(n_136), .Y(n_575) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_SL g159 ( .A(n_137), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_SL g166 ( .A(n_137), .Y(n_166) );
INVx2_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
BUFx3_ASAP7_75t_L g531 ( .A(n_137), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_137), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g559 ( .A(n_137), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_137), .B(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_137), .B(n_598), .Y(n_597) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_150), .B(n_159), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_147), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_143), .A2(n_210), .B1(n_267), .B2(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g549 ( .A(n_143), .Y(n_549) );
INVx4_ASAP7_75t_L g551 ( .A(n_143), .Y(n_551) );
INVx1_ASAP7_75t_L g603 ( .A(n_143), .Y(n_603) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_144), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_144), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx1_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
INVx1_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
INVx1_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_144), .Y(n_222) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
INVx2_ASAP7_75t_L g264 ( .A(n_144), .Y(n_264) );
INVx2_ASAP7_75t_L g195 ( .A(n_146), .Y(n_195) );
INVx1_ASAP7_75t_L g566 ( .A(n_146), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_147), .A2(n_173), .B(n_175), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_147), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_147), .A2(n_294), .B(n_295), .Y(n_293) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
INVx1_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
BUFx8_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B1(n_155), .B2(n_157), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_152), .A2(n_193), .B(n_194), .Y(n_192) );
INVx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g224 ( .A(n_154), .Y(n_224) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_158), .A2(n_169), .B(n_171), .Y(n_168) );
INVx1_ASAP7_75t_L g239 ( .A(n_158), .Y(n_239) );
INVx3_ASAP7_75t_L g548 ( .A(n_158), .Y(n_548) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_160), .A2(n_168), .B(n_172), .Y(n_167) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_160), .A2(n_186), .B(n_192), .Y(n_185) );
OAI21x1_ASAP7_75t_L g203 ( .A1(n_160), .A2(n_204), .B(n_207), .Y(n_203) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_160), .A2(n_232), .B(n_236), .Y(n_231) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_160), .A2(n_293), .B(n_296), .Y(n_292) );
BUFx10_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx10_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
INVx1_ASAP7_75t_L g538 ( .A(n_161), .Y(n_538) );
AND2x2_ASAP7_75t_L g254 ( .A(n_163), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g366 ( .A(n_163), .B(n_343), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_163), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g404 ( .A(n_164), .Y(n_404) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_164), .Y(n_409) );
AND2x2_ASAP7_75t_L g426 ( .A(n_164), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g316 ( .A(n_165), .B(n_256), .Y(n_316) );
INVx1_ASAP7_75t_L g330 ( .A(n_165), .Y(n_330) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_176), .Y(n_165) );
INVx1_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
INVx1_ASAP7_75t_L g536 ( .A(n_170), .Y(n_536) );
INVx1_ASAP7_75t_SL g552 ( .A(n_170), .Y(n_552) );
INVx1_ASAP7_75t_L g594 ( .A(n_174), .Y(n_594) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g184 ( .A(n_178), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_178), .B(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_178), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g225 ( .A(n_179), .Y(n_225) );
INVx2_ASAP7_75t_L g229 ( .A(n_179), .Y(n_229) );
NAND2x1_ASAP7_75t_L g180 ( .A(n_181), .B(n_197), .Y(n_180) );
AND2x4_ASAP7_75t_L g491 ( .A(n_181), .B(n_419), .Y(n_491) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
INVxp67_ASAP7_75t_SL g250 ( .A(n_182), .Y(n_250) );
BUFx3_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
INVx1_ASAP7_75t_L g351 ( .A(n_182), .Y(n_351) );
AND2x2_ASAP7_75t_L g354 ( .A(n_182), .B(n_200), .Y(n_354) );
AND2x2_ASAP7_75t_L g379 ( .A(n_182), .B(n_230), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_182), .Y(n_382) );
AND2x2_ASAP7_75t_L g414 ( .A(n_182), .B(n_279), .Y(n_414) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OAI21x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_196), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_184), .A2(n_185), .B(n_196), .Y(n_280) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_184), .A2(n_292), .B(n_301), .Y(n_291) );
OAI21xp33_ASAP7_75t_SL g319 ( .A1(n_184), .A2(n_292), .B(n_301), .Y(n_319) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_190), .C(n_191), .Y(n_186) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_191), .A2(n_208), .B(n_209), .Y(n_207) );
INVx6_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
O2A1O1Ixp5_ASAP7_75t_L g561 ( .A1(n_191), .A2(n_551), .B(n_562), .C(n_563), .Y(n_561) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_212), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g323 ( .A(n_199), .B(n_309), .Y(n_323) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g349 ( .A(n_201), .B(n_336), .Y(n_349) );
AND2x2_ASAP7_75t_L g378 ( .A(n_201), .B(n_214), .Y(n_378) );
OR2x2_ASAP7_75t_L g474 ( .A(n_201), .B(n_214), .Y(n_474) );
OAI21x1_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_202), .A2(n_231), .B(n_241), .Y(n_230) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_248) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_202), .A2(n_231), .B(n_241), .Y(n_279) );
INVx2_ASAP7_75t_L g217 ( .A(n_210), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_210), .A2(n_233), .B(n_234), .Y(n_232) );
AND2x2_ASAP7_75t_L g353 ( .A(n_212), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g502 ( .A(n_212), .Y(n_502) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_213), .Y(n_244) );
OR2x2_ASAP7_75t_L g436 ( .A(n_213), .B(n_246), .Y(n_436) );
INVx1_ASAP7_75t_L g458 ( .A(n_213), .Y(n_458) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_230), .Y(n_213) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g309 ( .A(n_214), .B(n_279), .Y(n_309) );
INVx1_ASAP7_75t_L g336 ( .A(n_214), .Y(n_336) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_214), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_214), .B(n_230), .Y(n_423) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_225), .A3(n_226), .B(n_227), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B1(n_221), .B2(n_223), .Y(n_215) );
INVx1_ASAP7_75t_L g585 ( .A(n_218), .Y(n_585) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_220), .A2(n_533), .B1(n_535), .B2(n_536), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_220), .A2(n_547), .B1(n_550), .B2(n_552), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_220), .A2(n_565), .B(n_567), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_220), .A2(n_223), .B1(n_573), .B2(n_574), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_220), .A2(n_552), .B1(n_584), .B2(n_586), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_220), .A2(n_223), .B1(n_593), .B2(n_595), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_220), .A2(n_223), .B1(n_602), .B2(n_604), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_220), .A2(n_223), .B1(n_618), .B2(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g596 ( .A(n_222), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_223), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g300 ( .A(n_224), .Y(n_300) );
INVx2_ASAP7_75t_L g258 ( .A(n_225), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_225), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_SL g587 ( .A(n_225), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
AO31x2_ASAP7_75t_L g571 ( .A1(n_226), .A2(n_572), .A3(n_575), .B(n_576), .Y(n_571) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_226), .A2(n_545), .A3(n_583), .B(n_587), .Y(n_582) );
AO31x2_ASAP7_75t_L g591 ( .A1(n_226), .A2(n_531), .A3(n_592), .B(n_597), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
BUFx2_ASAP7_75t_L g545 ( .A(n_229), .Y(n_545) );
AND2x2_ASAP7_75t_L g360 ( .A(n_230), .B(n_280), .Y(n_360) );
INVx2_ASAP7_75t_L g299 ( .A(n_235), .Y(n_299) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .Y(n_236) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR3x1_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .C(n_249), .Y(n_243) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_246), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g308 ( .A(n_246), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g359 ( .A(n_246), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g399 ( .A(n_246), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_246), .B(n_422), .Y(n_454) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_247), .B(n_335), .Y(n_395) );
AND2x2_ASAP7_75t_L g419 ( .A(n_247), .B(n_279), .Y(n_419) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g275 ( .A(n_248), .Y(n_275) );
BUFx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g430 ( .A(n_250), .B(n_309), .Y(n_430) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_253), .B(n_316), .Y(n_495) );
AND2x4_ASAP7_75t_L g487 ( .A(n_254), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_254), .B(n_307), .Y(n_501) );
INVx2_ASAP7_75t_L g303 ( .A(n_255), .Y(n_303) );
INVx1_ASAP7_75t_L g306 ( .A(n_255), .Y(n_306) );
INVx2_ASAP7_75t_L g391 ( .A(n_255), .Y(n_391) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g375 ( .A(n_256), .Y(n_375) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B(n_269), .Y(n_256) );
NOR2xp67_ASAP7_75t_SL g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g600 ( .A(n_258), .Y(n_600) );
INVx1_ASAP7_75t_L g553 ( .A(n_259), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_SL g534 ( .A(n_264), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_310), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_286), .B1(n_304), .B2(n_308), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_281), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g338 ( .A(n_274), .B(n_285), .Y(n_338) );
AND2x2_ASAP7_75t_L g498 ( .A(n_274), .B(n_379), .Y(n_498) );
BUFx2_ASAP7_75t_L g369 ( .A(n_275), .Y(n_369) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g368 ( .A(n_278), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g283 ( .A(n_279), .Y(n_283) );
INVx1_ASAP7_75t_L g335 ( .A(n_279), .Y(n_335) );
INVx1_ASAP7_75t_L g460 ( .A(n_280), .Y(n_460) );
AOI31xp33_ASAP7_75t_L g478 ( .A1(n_281), .A2(n_479), .A3(n_480), .B(n_481), .Y(n_478) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_282), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_283), .B(n_378), .Y(n_477) );
INVx2_ASAP7_75t_L g505 ( .A(n_283), .Y(n_505) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_284), .Y(n_320) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g333 ( .A(n_285), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_285), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g463 ( .A(n_285), .B(n_423), .Y(n_463) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_302), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g374 ( .A(n_290), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_300), .Y(n_296) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_306), .Y(n_327) );
INVx1_ASAP7_75t_L g367 ( .A(n_306), .Y(n_367) );
INVx1_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
AND2x2_ASAP7_75t_L g408 ( .A(n_307), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g464 ( .A(n_307), .B(n_391), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_308), .A2(n_381), .B(n_383), .Y(n_380) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_320), .Y(n_310) );
NAND3x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .C(n_317), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g482 ( .A(n_313), .B(n_402), .Y(n_482) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2x1_ASAP7_75t_SL g435 ( .A(n_315), .B(n_347), .Y(n_435) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g355 ( .A(n_316), .B(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_317), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_317), .B(n_426), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_317), .B(n_426), .Y(n_499) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g402 ( .A(n_319), .B(n_375), .Y(n_402) );
AND2x2_ASAP7_75t_L g322 ( .A(n_320), .B(n_323), .Y(n_322) );
AOI221x1_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B1(n_331), .B2(n_340), .C(n_344), .Y(n_321) );
AOI32xp33_ASAP7_75t_L g503 ( .A1(n_323), .A2(n_504), .A3(n_509), .B1(n_510), .B2(n_512), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_328), .B(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g342 ( .A(n_330), .B(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
OR2x2_ASAP7_75t_L g459 ( .A(n_330), .B(n_460), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_337), .C(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g381 ( .A(n_334), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g398 ( .A(n_334), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_337), .A2(n_434), .B1(n_436), .B2(n_437), .Y(n_433) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g511 ( .A(n_341), .Y(n_511) );
INVx2_ASAP7_75t_L g356 ( .A(n_343), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B(n_352), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g480 ( .A(n_349), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_350), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B1(n_357), .B2(n_359), .Y(n_352) );
AND2x4_ASAP7_75t_L g449 ( .A(n_355), .B(n_364), .Y(n_449) );
INVx1_ASAP7_75t_L g508 ( .A(n_356), .Y(n_508) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g387 ( .A(n_360), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_360), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_360), .B(n_388), .Y(n_479) );
AOI211x1_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_368), .B(n_370), .C(n_396), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR3x2_ASAP7_75t_L g471 ( .A(n_364), .B(n_366), .C(n_367), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_365), .A2(n_387), .B1(n_389), .B2(n_392), .Y(n_386) );
NOR2x1p5_ASAP7_75t_SL g365 ( .A(n_366), .B(n_367), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_366), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
INVx2_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_376), .B(n_380), .C(n_386), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_378), .B(n_382), .Y(n_393) );
INVx1_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_378), .B(n_485), .Y(n_493) );
OAI32xp33_ASAP7_75t_L g468 ( .A1(n_379), .A2(n_424), .A3(n_469), .B1(n_471), .B2(n_472), .Y(n_468) );
INVx1_ASAP7_75t_L g485 ( .A(n_379), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_379), .B(n_399), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_382), .B(n_416), .Y(n_451) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g429 ( .A(n_388), .B(n_414), .Y(n_429) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g438 ( .A(n_391), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g406 ( .A(n_394), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B1(n_405), .B2(n_407), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g444 ( .A(n_401), .Y(n_444) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g425 ( .A(n_402), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_402), .B(n_409), .Y(n_513) );
INVx1_ASAP7_75t_SL g439 ( .A(n_403), .Y(n_439) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_433), .C(n_440), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_424), .B(n_428), .Y(n_411) );
NOR2xp33_ASAP7_75t_SL g412 ( .A(n_413), .B(n_417), .Y(n_412) );
INVxp67_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g432 ( .A(n_426), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g441 ( .A(n_429), .Y(n_441) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_434), .A2(n_485), .B1(n_486), .B2(n_489), .C(n_490), .Y(n_484) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI32xp33_ASAP7_75t_L g440 ( .A1(n_437), .A2(n_441), .A3(n_442), .B1(n_443), .B2(n_445), .Y(n_440) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_443), .A2(n_453), .B1(n_454), .B2(n_455), .C(n_461), .Y(n_452) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_465), .C(n_483), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B(n_452), .Y(n_447) );
AOI211x1_ASAP7_75t_L g465 ( .A1(n_448), .A2(n_466), .B(n_468), .C(n_475), .Y(n_465) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2x1_ASAP7_75t_SL g456 ( .A(n_457), .B(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g467 ( .A(n_458), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AO21x1_ASAP7_75t_L g475 ( .A1(n_464), .A2(n_476), .B(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g509 ( .A(n_480), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI21xp33_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_492), .B(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g506 ( .A(n_505), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_514), .A2(n_521), .B(n_833), .C(n_844), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_514), .A2(n_834), .B(n_835), .Y(n_833) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g834 ( .A(n_523), .Y(n_834) );
NAND4xp75_ASAP7_75t_L g523 ( .A(n_524), .B(n_673), .C(n_749), .D(n_801), .Y(n_523) );
AND3x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_646), .C(n_659), .Y(n_524) );
AOI221x1_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_578), .B1(n_607), .B2(n_611), .C(n_623), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_526), .A2(n_647), .B(n_649), .C(n_650), .Y(n_646) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_541), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g610 ( .A(n_530), .Y(n_610) );
BUFx2_ASAP7_75t_L g628 ( .A(n_530), .Y(n_628) );
OR2x2_ASAP7_75t_L g670 ( .A(n_530), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g677 ( .A(n_530), .B(n_544), .Y(n_677) );
AND2x4_ASAP7_75t_L g712 ( .A(n_530), .B(n_543), .Y(n_712) );
OR2x2_ASAP7_75t_L g755 ( .A(n_530), .B(n_571), .Y(n_755) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .A3(n_537), .B(n_539), .Y(n_530) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_537), .A2(n_600), .A3(n_601), .B(n_605), .Y(n_599) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g568 ( .A(n_538), .Y(n_568) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_556), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_543), .B(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_543), .Y(n_642) );
INVx2_ASAP7_75t_L g669 ( .A(n_543), .Y(n_669) );
INVx3_ASAP7_75t_L g682 ( .A(n_543), .Y(n_682) );
AND2x2_ASAP7_75t_L g800 ( .A(n_543), .B(n_629), .Y(n_800) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g609 ( .A(n_544), .B(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g665 ( .A(n_544), .Y(n_665) );
AO31x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .A3(n_553), .B(n_554), .Y(n_544) );
AO31x2_ASAP7_75t_L g616 ( .A1(n_553), .A2(n_600), .A3(n_617), .B(n_620), .Y(n_616) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g685 ( .A(n_557), .Y(n_685) );
INVx1_ASAP7_75t_L g812 ( .A(n_557), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_570), .Y(n_557) );
AND2x2_ASAP7_75t_L g608 ( .A(n_558), .B(n_571), .Y(n_608) );
INVx1_ASAP7_75t_L g671 ( .A(n_558), .Y(n_671) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_569), .Y(n_558) );
OAI21x1_ASAP7_75t_L g630 ( .A1(n_559), .A2(n_560), .B(n_569), .Y(n_630) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B(n_568), .Y(n_560) );
INVx2_ASAP7_75t_L g626 ( .A(n_570), .Y(n_626) );
AND2x2_ASAP7_75t_L g678 ( .A(n_570), .B(n_629), .Y(n_678) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g640 ( .A(n_571), .Y(n_640) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_571), .Y(n_700) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_580), .A2(n_672), .B1(n_676), .B2(n_679), .Y(n_675) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_589), .Y(n_580) );
INVx1_ASAP7_75t_L g693 ( .A(n_581), .Y(n_693) );
BUFx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g613 ( .A(n_582), .B(n_591), .Y(n_613) );
AND2x2_ASAP7_75t_L g644 ( .A(n_582), .B(n_599), .Y(n_644) );
INVx4_ASAP7_75t_SL g655 ( .A(n_582), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_582), .B(n_689), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_582), .B(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g726 ( .A(n_590), .B(n_704), .Y(n_726) );
OR2x2_ASAP7_75t_L g759 ( .A(n_590), .B(n_741), .Y(n_759) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_599), .Y(n_590) );
INVx2_ASAP7_75t_L g633 ( .A(n_591), .Y(n_633) );
INVx1_ASAP7_75t_L g638 ( .A(n_591), .Y(n_638) );
AND2x2_ASAP7_75t_L g645 ( .A(n_591), .B(n_615), .Y(n_645) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_591), .Y(n_661) );
INVx1_ASAP7_75t_L g689 ( .A(n_591), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_591), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g622 ( .A(n_599), .Y(n_622) );
AND2x4_ASAP7_75t_L g632 ( .A(n_599), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g658 ( .A(n_599), .Y(n_658) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_599), .Y(n_735) );
INVx1_ASAP7_75t_L g828 ( .A(n_599), .Y(n_828) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_608), .B(n_681), .Y(n_748) );
AND2x2_ASAP7_75t_L g761 ( .A(n_608), .B(n_677), .Y(n_761) );
AND2x2_ASAP7_75t_L g831 ( .A(n_608), .B(n_682), .Y(n_831) );
AND2x4_ASAP7_75t_L g666 ( .A(n_610), .B(n_629), .Y(n_666) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g733 ( .A(n_613), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g747 ( .A(n_613), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_613), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g649 ( .A(n_614), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_614), .B(n_687), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g743 ( .A1(n_614), .A2(n_744), .B(n_747), .C(n_748), .Y(n_743) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_622), .Y(n_614) );
AND2x2_ASAP7_75t_L g714 ( .A(n_615), .B(n_655), .Y(n_714) );
INVx3_ASAP7_75t_L g741 ( .A(n_615), .Y(n_741) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g636 ( .A(n_616), .Y(n_636) );
AND2x4_ASAP7_75t_L g662 ( .A(n_616), .B(n_622), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_622), .B(n_655), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_631), .B1(n_639), .B2(n_643), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g780 ( .A(n_625), .Y(n_780) );
AND2x4_ASAP7_75t_L g691 ( .A(n_626), .B(n_671), .Y(n_691) );
INVx1_ASAP7_75t_L g711 ( .A(n_626), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_628), .A2(n_684), .B1(n_694), .B2(n_696), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_628), .B(n_685), .Y(n_742) );
NAND2x1_ASAP7_75t_L g799 ( .A(n_628), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g814 ( .A(n_628), .Y(n_814) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx2_ASAP7_75t_L g753 ( .A(n_630), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
AND2x2_ASAP7_75t_L g672 ( .A(n_632), .B(n_654), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_632), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_632), .B(n_714), .Y(n_713) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_632), .Y(n_787) );
NAND2x1p5_ASAP7_75t_L g794 ( .A(n_632), .B(n_695), .Y(n_794) );
AND2x4_ASAP7_75t_L g817 ( .A(n_632), .B(n_745), .Y(n_817) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx3_ASAP7_75t_L g695 ( .A(n_635), .Y(n_695) );
AND2x2_ASAP7_75t_L g707 ( .A(n_635), .B(n_700), .Y(n_707) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g657 ( .A(n_636), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g705 ( .A(n_636), .Y(n_705) );
INVx1_ASAP7_75t_L g648 ( .A(n_637), .Y(n_648) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g805 ( .A(n_638), .B(n_655), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g731 ( .A(n_640), .B(n_712), .Y(n_731) );
INVx2_ASAP7_75t_L g772 ( .A(n_640), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_640), .B(n_666), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_641), .B(n_691), .Y(n_821) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_644), .B(n_704), .Y(n_703) );
AND2x4_ASAP7_75t_L g716 ( .A(n_644), .B(n_661), .Y(n_716) );
INVx1_ASAP7_75t_L g808 ( .A(n_644), .Y(n_808) );
AND2x2_ASAP7_75t_L g807 ( .A(n_645), .B(n_734), .Y(n_807) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_649), .A2(n_779), .B1(n_781), .B2(n_783), .Y(n_778) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g687 ( .A(n_655), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g723 ( .A(n_655), .Y(n_723) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_655), .Y(n_729) );
INVx2_ASAP7_75t_L g746 ( .A(n_655), .Y(n_746) );
OR2x2_ASAP7_75t_L g767 ( .A(n_655), .B(n_730), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_655), .B(n_725), .Y(n_777) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g744 ( .A(n_657), .B(n_745), .Y(n_744) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_657), .Y(n_798) );
INVx1_ASAP7_75t_L g725 ( .A(n_658), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_667), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_662), .B(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g730 ( .A(n_662), .Y(n_730) );
AND2x2_ASAP7_75t_L g804 ( .A(n_662), .B(n_805), .Y(n_804) );
AOI211x1_ASAP7_75t_SL g732 ( .A1(n_663), .A2(n_733), .B(n_736), .C(n_743), .Y(n_732) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g789 ( .A(n_665), .B(n_666), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_666), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_666), .Y(n_782) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_672), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g697 ( .A(n_669), .Y(n_697) );
NOR2x1p5_ASAP7_75t_L g754 ( .A(n_669), .B(n_755), .Y(n_754) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_670), .B(n_699), .Y(n_698) );
NOR2xp67_ASAP7_75t_SL g771 ( .A(n_670), .B(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g832 ( .A(n_672), .B(n_740), .Y(n_832) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_717), .Y(n_673) );
NAND3xp33_ASAP7_75t_SL g674 ( .A(n_675), .B(n_683), .C(n_701), .Y(n_674) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_677), .Y(n_708) );
AND2x2_ASAP7_75t_L g715 ( .A(n_677), .B(n_711), .Y(n_715) );
AND2x4_ASAP7_75t_SL g829 ( .A(n_677), .B(n_691), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_678), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_680), .A2(n_722), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g811 ( .A(n_682), .B(n_812), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_690), .B2(n_692), .Y(n_684) );
NAND2x1_ASAP7_75t_L g760 ( .A(n_687), .B(n_740), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_687), .B(n_734), .Y(n_770) );
INVx1_ASAP7_75t_L g797 ( .A(n_687), .Y(n_797) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_690), .A2(n_816), .B(n_819), .Y(n_815) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_691), .A2(n_703), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g776 ( .A(n_695), .Y(n_776) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g720 ( .A(n_698), .Y(n_720) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_708), .B1(n_709), .B2(n_713), .C1(n_715), .C2(n_716), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g736 ( .A1(n_703), .A2(n_737), .B(n_742), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_704), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g818 ( .A(n_704), .Y(n_818) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_705), .Y(n_824) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
AND2x2_ASAP7_75t_L g788 ( .A(n_710), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g781 ( .A(n_711), .B(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_732), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_727), .B2(n_731), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_726), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g738 ( .A(n_724), .Y(n_738) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx4_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g766 ( .A(n_741), .B(n_758), .Y(n_766) );
OR2x2_ASAP7_75t_L g826 ( .A(n_741), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND5xp2_ASAP7_75t_L g802 ( .A(n_747), .B(n_794), .C(n_803), .D(n_806), .E(n_808), .Y(n_802) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_785), .Y(n_749) );
NAND2xp67_ASAP7_75t_SL g750 ( .A(n_751), .B(n_768), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_756), .B1(n_761), .B2(n_762), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND3xp33_ASAP7_75t_SL g756 ( .A(n_757), .B(n_759), .C(n_760), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g791 ( .A(n_760), .Y(n_791) );
NAND3xp33_ASAP7_75t_SL g762 ( .A(n_763), .B(n_766), .C(n_767), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g784 ( .A(n_765), .Y(n_784) );
O2A1O1Ixp33_ASAP7_75t_SL g796 ( .A1(n_766), .A2(n_797), .B(n_798), .C(n_799), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_773), .B2(n_774), .C(n_778), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_775), .B(n_823), .Y(n_822) );
OR2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
INVx1_ASAP7_75t_L g792 ( .A(n_779), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_790), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g795 ( .A(n_789), .Y(n_795) );
AOI211xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B(n_793), .C(n_796), .Y(n_790) );
AOI211x1_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_809), .B(n_815), .C(n_830), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2x1p5_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NAND2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_822), .B1(n_825), .B2(n_829), .Y(n_819) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g844 ( .A(n_835), .B(n_845), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx5_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx10_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_848), .B(n_889), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_853), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx8_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_878), .Y(n_853) );
AOI31xp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_866), .A3(n_867), .B(n_872), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_855), .B(n_880), .Y(n_879) );
AO22x1_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_858), .B1(n_864), .B2(n_865), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_856), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_858), .Y(n_865) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g881 ( .A(n_866), .Y(n_881) );
INVx1_ASAP7_75t_L g880 ( .A(n_867), .Y(n_880) );
BUFx2_ASAP7_75t_SL g867 ( .A(n_868), .Y(n_867) );
INVx4_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NOR2x1p5_ASAP7_75t_L g887 ( .A(n_870), .B(n_888), .Y(n_887) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g876 ( .A(n_871), .Y(n_876) );
NOR2xp33_ASAP7_75t_SL g872 ( .A(n_873), .B(n_877), .Y(n_872) );
INVx5_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_881), .Y(n_878) );
BUFx10_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
BUFx6f_ASAP7_75t_L g893 ( .A(n_883), .Y(n_893) );
INVx6_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NAND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
endmodule