module fake_jpeg_25373_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_34),
.B1(n_42),
.B2(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_66),
.B1(n_72),
.B2(n_79),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_37),
.B1(n_42),
.B2(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

HAxp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_21),
.CON(n_69),
.SN(n_69)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_83),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_77),
.Y(n_91)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_43),
.B1(n_40),
.B2(n_32),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_39),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_22),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_31),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_20),
.B1(n_22),
.B2(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_25),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_0),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_62),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_39),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_104),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_22),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_36),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_81),
.B1(n_61),
.B2(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_123),
.B1(n_132),
.B2(n_103),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_72),
.B1(n_79),
.B2(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_92),
.B1(n_93),
.B2(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_118),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_16),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_129),
.Y(n_149)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_16),
.B(n_65),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_131),
.B(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_76),
.B1(n_65),
.B2(n_80),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_67),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_59),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_2),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_155),
.B1(n_120),
.B2(n_130),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_114),
.B1(n_121),
.B2(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_146),
.B(n_116),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_91),
.C(n_96),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_145),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_89),
.B1(n_91),
.B2(n_108),
.C(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_153),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_96),
.A3(n_104),
.B1(n_89),
.B2(n_111),
.C1(n_105),
.C2(n_100),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_101),
.C(n_111),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_111),
.B1(n_103),
.B2(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_90),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_162),
.B1(n_167),
.B2(n_168),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_173),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_118),
.B1(n_119),
.B2(n_127),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_169),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_3),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_11),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_172),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_10),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_10),
.B(n_11),
.Y(n_174)
);

NAND2xp67_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_168),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_139),
.C(n_141),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_154),
.C(n_153),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_188),
.B1(n_170),
.B2(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_156),
.C(n_137),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_137),
.C(n_151),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_160),
.B(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_176),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_173),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_169),
.B(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_164),
.B1(n_159),
.B2(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_198),
.A2(n_176),
.B1(n_183),
.B2(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_203),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_195),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_177),
.B1(n_181),
.B2(n_140),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_186),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_181),
.B(n_12),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_189),
.B(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_189),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_204),
.B(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_208),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_12),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_214),
.A2(n_210),
.B(n_200),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_218),
.B(n_219),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_215),
.C(n_12),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_221),
.B(n_13),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_13),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_220),
.Y(n_224)
);


endmodule