module fake_aes_8359_n_741 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_741, n_389);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_741;
output n_389;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_79), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_26), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_32), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_57), .Y(n_84) );
INVxp33_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_10), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_13), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_62), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_36), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_76), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_61), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_38), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_43), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_39), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_45), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_9), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_51), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_67), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_68), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_46), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_27), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_4), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_3), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_29), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_35), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_54), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_52), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_5), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_3), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_37), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_22), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_16), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_50), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_34), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_66), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_16), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_33), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_44), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_101), .B(n_0), .Y(n_132) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_89), .A2(n_40), .B(n_78), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
CKINVDCx6p67_ASAP7_75t_R g135 ( .A(n_105), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_107), .B(n_0), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_101), .B(n_1), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
BUFx12f_ASAP7_75t_L g140 ( .A(n_113), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_128), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_128), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_109), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_88), .B(n_94), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_87), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_120), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_107), .B(n_2), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_85), .B(n_5), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_120), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_92), .B(n_47), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_88), .B(n_6), .Y(n_160) );
AND2x6_ASAP7_75t_L g161 ( .A(n_93), .B(n_49), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_102), .B(n_53), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_109), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_95), .Y(n_165) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_95), .B(n_80), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_96), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_94), .B(n_7), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_96), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_106), .B(n_7), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_97), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_97), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_111), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_137), .B(n_98), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
BUFx2_ASAP7_75t_SL g179 ( .A(n_170), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_144), .B(n_108), .Y(n_182) );
INVx4_ASAP7_75t_SL g183 ( .A(n_159), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_160), .B(n_86), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_144), .B(n_113), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_164), .B(n_121), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_164), .B(n_110), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_160), .B(n_116), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_135), .B(n_121), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_137), .B(n_130), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_141), .B(n_129), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_173), .B(n_112), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_140), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_170), .B(n_118), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_154), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_141), .B(n_127), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_140), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_135), .A2(n_87), .B1(n_99), .B2(n_123), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_140), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_166), .B(n_98), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_154), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_147), .B(n_126), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
AO22x2_ASAP7_75t_L g214 ( .A1(n_152), .A2(n_125), .B1(n_124), .B2(n_81), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_134), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_135), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_160), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
AO22x2_ASAP7_75t_L g220 ( .A1(n_152), .A2(n_100), .B1(n_117), .B2(n_115), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_156), .B(n_99), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_147), .B(n_104), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_160), .B(n_103), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_148), .B(n_84), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_159), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_148), .B(n_83), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_149), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_149), .B(n_82), .Y(n_229) );
INVxp67_ASAP7_75t_L g230 ( .A(n_156), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_151), .Y(n_231) );
INVxp33_ASAP7_75t_L g232 ( .A(n_132), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_151), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_132), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_165), .B(n_122), .Y(n_237) );
INVx5_ASAP7_75t_L g238 ( .A(n_159), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_167), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_167), .B(n_42), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_210), .A2(n_166), .B1(n_138), .B2(n_168), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_190), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_224), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_189), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
INVx3_ASAP7_75t_SL g249 ( .A(n_216), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_210), .A2(n_166), .B1(n_161), .B2(n_159), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
BUFx12f_ASAP7_75t_L g252 ( .A(n_200), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_226), .B(n_171), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_232), .B(n_171), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_226), .B(n_169), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_179), .B(n_138), .Y(n_257) );
BUFx4f_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_178), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_232), .B(n_169), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_182), .B(n_145), .Y(n_261) );
AND2x6_ASAP7_75t_SL g262 ( .A(n_197), .B(n_145), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_207), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_230), .B(n_168), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_198), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_236), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_208), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_225), .A2(n_161), .B1(n_159), .B2(n_163), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_225), .A2(n_161), .B1(n_159), .B2(n_172), .Y(n_271) );
BUFx12f_ASAP7_75t_L g272 ( .A(n_191), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_221), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_197), .Y(n_275) );
OR2x2_ASAP7_75t_SL g276 ( .A(n_214), .B(n_133), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_191), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_205), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_203), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_201), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_190), .Y(n_282) );
NOR2xp67_ASAP7_75t_L g283 ( .A(n_186), .B(n_158), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_188), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_182), .B(n_157), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_211), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_230), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_228), .B(n_161), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_213), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_214), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_184), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_231), .B(n_161), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_184), .B(n_157), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_184), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_233), .B(n_161), .Y(n_295) );
BUFx8_ASAP7_75t_L g296 ( .A(n_223), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_214), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_237), .B(n_155), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_192), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_220), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_183), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_192), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_205), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_192), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_209), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_238), .B(n_172), .Y(n_306) );
NOR2xp33_ASAP7_75t_R g307 ( .A(n_234), .B(n_161), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_223), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_183), .Y(n_309) );
INVx5_ASAP7_75t_L g310 ( .A(n_224), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_183), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_227), .B(n_158), .Y(n_312) );
AOI21xp5_ASAP7_75t_SL g313 ( .A1(n_242), .A2(n_234), .B(n_133), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
NOR3xp33_ASAP7_75t_L g315 ( .A(n_275), .B(n_212), .C(n_222), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_243), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_263), .A2(n_220), .B1(n_218), .B2(n_161), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_296), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_264), .B(n_235), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_243), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_284), .B(n_239), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_266), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_268), .B(n_238), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_275), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_296), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_264), .B(n_261), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_244), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_264), .B(n_196), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_248), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_277), .A2(n_220), .B1(n_212), .B2(n_238), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_261), .A2(n_195), .B1(n_229), .B2(n_222), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_257), .B(n_177), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_251), .Y(n_335) );
BUFx12f_ASAP7_75t_L g336 ( .A(n_272), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_282), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_256), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_241), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_290), .A2(n_229), .B1(n_204), .B2(n_196), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_297), .A2(n_204), .B1(n_195), .B2(n_177), .Y(n_342) );
OAI22x1_ASAP7_75t_L g343 ( .A1(n_300), .A2(n_133), .B1(n_158), .B2(n_153), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_257), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_250), .A2(n_240), .B1(n_153), .B2(n_150), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_282), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_272), .B(n_238), .Y(n_347) );
OAI22xp5_ASAP7_75t_SL g348 ( .A1(n_263), .A2(n_133), .B1(n_157), .B2(n_155), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_241), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_257), .B(n_157), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_291), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_282), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_291), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_304), .A2(n_240), .B1(n_150), .B2(n_153), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_254), .B(n_155), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_287), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_274), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_282), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_277), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_294), .A2(n_172), .B1(n_150), .B2(n_155), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_247), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_252), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_299), .A2(n_172), .B1(n_142), .B2(n_143), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_301), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_302), .A2(n_172), .B1(n_142), .B2(n_143), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_273), .A2(n_172), .B1(n_142), .B2(n_143), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_281), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_336), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_319), .A2(n_246), .B1(n_269), .B2(n_252), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_355), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_359), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_328), .B(n_260), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_321), .B(n_308), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_313), .A2(n_295), .B(n_292), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_364), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_313), .A2(n_288), .B(n_255), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_364), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_319), .A2(n_269), .B1(n_249), .B2(n_258), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_318), .A2(n_285), .B1(n_293), .B2(n_258), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_336), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_362), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_323), .A2(n_276), .B1(n_270), .B2(n_271), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_330), .B(n_285), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_333), .B(n_298), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_339), .A2(n_255), .B(n_253), .Y(n_387) );
AOI211x1_ASAP7_75t_L g388 ( .A1(n_332), .A2(n_259), .B(n_289), .C(n_286), .Y(n_388) );
UNKNOWN g389 ( );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_321), .A2(n_249), .B1(n_283), .B2(n_262), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_351), .A2(n_293), .B1(n_279), .B2(n_280), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_356), .A2(n_253), .B1(n_306), .B2(n_307), .C(n_131), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
INVx4_ASAP7_75t_L g394 ( .A(n_364), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_349), .Y(n_395) );
INVx5_ASAP7_75t_L g396 ( .A(n_364), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_355), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_359), .B(n_312), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_317), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_396), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_386), .A2(n_351), .B1(n_315), .B2(n_353), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_381), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_386), .B(n_320), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_371), .A2(n_327), .B1(n_326), .B2(n_334), .Y(n_405) );
OR2x2_ASAP7_75t_SL g406 ( .A(n_399), .B(n_340), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_372), .B(n_333), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_389), .B(n_357), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_396), .B(n_344), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_396), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
OAI211xp5_ASAP7_75t_L g412 ( .A1(n_369), .A2(n_342), .B(n_326), .C(n_353), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_393), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_350), .B1(n_327), .B2(n_334), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_385), .B(n_329), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_393), .B(n_350), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_384), .A2(n_334), .B1(n_348), .B2(n_345), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_395), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_366), .B(n_345), .C(n_367), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_370), .A2(n_350), .B1(n_334), .B2(n_357), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_396), .B(n_350), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_397), .A2(n_334), .B1(n_348), .B2(n_338), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_373), .A2(n_362), .B1(n_314), .B2(n_324), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_373), .A2(n_335), .B1(n_338), .B2(n_329), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_390), .A2(n_354), .B1(n_331), .B2(n_360), .C(n_335), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_399), .B(n_373), .Y(n_429) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_403), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_404), .B(n_375), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_404), .B(n_375), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_416), .B(n_400), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_417), .A2(n_407), .B(n_377), .Y(n_435) );
OAI21x1_ASAP7_75t_L g436 ( .A1(n_417), .A2(n_374), .B(n_376), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_416), .B(n_400), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_413), .A2(n_374), .B(n_387), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_423), .A2(n_373), .B1(n_331), .B2(n_379), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_415), .B(n_388), .Y(n_440) );
OA21x2_ASAP7_75t_L g441 ( .A1(n_403), .A2(n_187), .B(n_180), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_413), .B(n_394), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_418), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_418), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_421), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_415), .A2(n_366), .B(n_314), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_425), .A2(n_396), .B1(n_394), .B2(n_378), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_412), .A2(n_383), .B1(n_368), .B2(n_382), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_421), .B(n_376), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_414), .A2(n_394), .B1(n_376), .B2(n_324), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
OAI222xp33_ASAP7_75t_L g454 ( .A1(n_405), .A2(n_383), .B1(n_368), .B2(n_382), .C1(n_361), .C2(n_14), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_402), .A2(n_343), .B1(n_392), .B2(n_347), .C1(n_325), .C2(n_378), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_427), .B(n_419), .C(n_420), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_408), .B(n_365), .C(n_363), .D(n_142), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_401), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_401), .B(n_378), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_411), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_426), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_429), .A2(n_378), .B1(n_352), .B2(n_316), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_411), .A2(n_343), .B(n_378), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_401), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_406), .A2(n_322), .B1(n_316), .B2(n_352), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_424), .A2(n_322), .B1(n_316), .B2(n_346), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_454), .B(n_408), .C(n_410), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_432), .B(n_428), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_457), .A2(n_406), .B1(n_422), .B2(n_409), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_439), .A2(n_422), .B1(n_409), .B2(n_316), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_445), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_431), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_466), .B(n_422), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_445), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_450), .B(n_143), .C(n_131), .D(n_422), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_466), .B(n_409), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_432), .B(n_409), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_456), .B(n_139), .C(n_134), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_433), .B(n_8), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_466), .B(n_10), .Y(n_484) );
NAND3xp33_ASAP7_75t_SL g485 ( .A(n_455), .B(n_307), .C(n_12), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_458), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_433), .B(n_11), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_446), .B(n_11), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_456), .A2(n_322), .B1(n_316), .B2(n_346), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_447), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_457), .A2(n_322), .B1(n_358), .B2(n_346), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_458), .Y(n_493) );
NAND3xp33_ASAP7_75t_SL g494 ( .A(n_455), .B(n_14), .C(n_15), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_444), .B(n_17), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_453), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_463), .A2(n_449), .B(n_444), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_444), .B(n_17), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_458), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_436), .B(n_19), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_460), .B(n_139), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_434), .B(n_364), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_435), .B(n_139), .Y(n_507) );
OR2x6_ASAP7_75t_L g508 ( .A(n_465), .B(n_322), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_435), .B(n_453), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_434), .B(n_437), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_464), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_452), .A2(n_440), .B1(n_465), .B2(n_467), .C(n_448), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_461), .B(n_139), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_440), .B(n_131), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_451), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_442), .B(n_139), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_467), .B(n_358), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_464), .B(n_131), .C(n_180), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_442), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_486), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_468), .B(n_134), .C(n_139), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_472), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_509), .B(n_436), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_516), .B(n_459), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_485), .A2(n_448), .B1(n_449), .B2(n_438), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_511), .B(n_459), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_509), .B(n_438), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_503), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_494), .A2(n_462), .B(n_459), .Y(n_534) );
OAI21xp5_ASAP7_75t_SL g535 ( .A1(n_478), .A2(n_459), .B(n_134), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_507), .B(n_438), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_507), .B(n_438), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_469), .B(n_441), .Y(n_538) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_475), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_503), .B(n_441), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_491), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_489), .A2(n_441), .B(n_187), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_480), .B(n_441), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_474), .B(n_134), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_522), .B(n_358), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
AND2x4_ASAP7_75t_SL g549 ( .A(n_479), .B(n_337), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_510), .Y(n_550) );
OAI33xp33_ASAP7_75t_L g551 ( .A1(n_483), .A2(n_219), .A3(n_209), .B1(n_306), .B2(n_25), .B3(n_30), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_473), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_517), .B(n_337), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_484), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_475), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_521), .B(n_337), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_481), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_489), .A2(n_219), .B(n_278), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_474), .B(n_185), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_487), .B(n_20), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_479), .B(n_174), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_500), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_481), .B(n_502), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_484), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_21), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_488), .B(n_174), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_500), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_493), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_493), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_512), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_495), .B(n_174), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_495), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_499), .B(n_506), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_499), .B(n_174), .Y(n_574) );
BUFx3_ASAP7_75t_L g575 ( .A(n_500), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_508), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_470), .A2(n_175), .B1(n_185), .B2(n_176), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_512), .B(n_175), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_488), .B(n_23), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_514), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_501), .B(n_175), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_501), .B(n_175), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_515), .B(n_247), .C(n_265), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_502), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_518), .B(n_185), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_533), .B(n_515), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_525), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_543), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_530), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_541), .B(n_518), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_544), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_532), .B(n_498), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_555), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_535), .B(n_482), .C(n_513), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_532), .B(n_504), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_539), .B(n_500), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_570), .B(n_471), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_531), .B(n_508), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_528), .A2(n_492), .B(n_504), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_560), .A2(n_504), .B(n_490), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_526), .B(n_505), .Y(n_603) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_545), .B(n_520), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_568), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_548), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_550), .B(n_505), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_526), .B(n_508), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_528), .B(n_519), .C(n_508), .D(n_303), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_554), .B(n_519), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_564), .B(n_185), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_572), .B(n_527), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_540), .B(n_176), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_546), .B(n_176), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_546), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_536), .B(n_176), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_585), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_580), .B(n_31), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_582), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_563), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_536), .B(n_537), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_536), .B(n_55), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_563), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_523), .B(n_56), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_569), .B(n_58), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_537), .B(n_59), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_560), .A2(n_217), .B1(n_215), .B2(n_305), .C(n_303), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_573), .B(n_63), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_538), .B(n_64), .Y(n_629) );
NOR2x1p5_ASAP7_75t_L g630 ( .A(n_524), .B(n_217), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_543), .B(n_69), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_552), .B(n_70), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_537), .B(n_71), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_552), .B(n_72), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_557), .Y(n_635) );
OAI32xp33_ASAP7_75t_L g636 ( .A1(n_565), .A2(n_73), .A3(n_74), .B1(n_75), .B2(n_77), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_567), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_557), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_576), .B(n_215), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_566), .Y(n_640) );
OAI31xp33_ASAP7_75t_L g641 ( .A1(n_577), .A2(n_278), .A3(n_305), .B(n_267), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_566), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_601), .A2(n_534), .B1(n_577), .B2(n_584), .C(n_558), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_588), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_590), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_603), .B(n_576), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_591), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_594), .B(n_576), .Y(n_648) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_596), .B(n_562), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_594), .B(n_567), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_619), .B(n_575), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_604), .B(n_549), .Y(n_652) );
XNOR2xp5_ASAP7_75t_L g653 ( .A(n_605), .B(n_549), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_593), .B(n_575), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_620), .B(n_553), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_606), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_623), .B(n_542), .Y(n_658) );
XOR2x2_ASAP7_75t_L g659 ( .A(n_597), .B(n_547), .Y(n_659) );
NAND2x1_ASAP7_75t_L g660 ( .A(n_595), .B(n_562), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_SL g661 ( .A1(n_602), .A2(n_579), .B(n_578), .C(n_556), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_603), .B(n_562), .Y(n_662) );
AOI31xp33_ASAP7_75t_L g663 ( .A1(n_599), .A2(n_551), .A3(n_561), .B(n_559), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_595), .B(n_562), .Y(n_664) );
XOR2x2_ASAP7_75t_L g665 ( .A(n_597), .B(n_561), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_612), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_615), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_607), .Y(n_668) );
XNOR2x1_ASAP7_75t_L g669 ( .A(n_608), .B(n_559), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_599), .A2(n_574), .B(n_571), .C(n_586), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_592), .Y(n_671) );
XNOR2x2_ASAP7_75t_L g672 ( .A(n_609), .B(n_586), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_621), .B(n_583), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_635), .Y(n_674) );
XNOR2x2_ASAP7_75t_L g675 ( .A(n_622), .B(n_583), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_638), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_641), .A2(n_636), .B(n_627), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_587), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_589), .B(n_581), .Y(n_679) );
AND3x1_ASAP7_75t_L g680 ( .A(n_608), .B(n_267), .C(n_265), .Y(n_680) );
OA22x2_ASAP7_75t_L g681 ( .A1(n_622), .A2(n_301), .B1(n_309), .B2(n_311), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_610), .B(n_215), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_600), .B(n_215), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_611), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_637), .B(n_217), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_640), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_630), .B(n_301), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_626), .B(n_309), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_616), .A2(n_217), .B(n_245), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_626), .A2(n_309), .B1(n_311), .B2(n_310), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_640), .Y(n_691) );
OR2x6_ASAP7_75t_L g692 ( .A(n_633), .B(n_311), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_642), .B(n_245), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_598), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_642), .B(n_245), .Y(n_695) );
XNOR2x2_ASAP7_75t_SL g696 ( .A(n_633), .B(n_245), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_598), .A2(n_628), .B(n_625), .C(n_624), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_613), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_616), .A2(n_310), .B1(n_639), .B2(n_618), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_629), .A2(n_310), .B1(n_614), .B2(n_639), .C1(n_631), .C2(n_632), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_613), .B(n_310), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_634), .B(n_620), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_588), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_666), .B(n_678), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_694), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_652), .B(n_653), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_662), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_671), .B(n_668), .Y(n_708) );
AOI21xp33_ASAP7_75t_SL g709 ( .A1(n_649), .A2(n_663), .B(n_681), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_663), .A2(n_643), .B(n_677), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_680), .A2(n_643), .B1(n_692), .B2(n_670), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_692), .A2(n_669), .B1(n_688), .B2(n_648), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_696), .A2(n_660), .B(n_661), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_648), .A2(n_650), .B1(n_675), .B2(n_699), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_672), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_646), .B(n_673), .Y(n_716) );
XOR2x2_ASAP7_75t_L g717 ( .A(n_659), .B(n_665), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_650), .A2(n_658), .B1(n_664), .B2(n_651), .Y(n_718) );
AO22x2_ASAP7_75t_L g719 ( .A1(n_714), .A2(n_644), .B1(n_645), .B2(n_647), .Y(n_719) );
AO22x2_ASAP7_75t_L g720 ( .A1(n_710), .A2(n_656), .B1(n_703), .B2(n_657), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_713), .A2(n_677), .B(n_651), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_711), .B(n_700), .C(n_697), .D(n_690), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_715), .B(n_687), .Y(n_723) );
XNOR2x2_ASAP7_75t_L g724 ( .A(n_717), .B(n_683), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_718), .A2(n_703), .B1(n_667), .B2(n_691), .C(n_686), .Y(n_725) );
AO22x2_ASAP7_75t_L g726 ( .A1(n_712), .A2(n_676), .B1(n_674), .B2(n_702), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_721), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_722), .A2(n_711), .B1(n_706), .B2(n_704), .Y(n_728) );
O2A1O1Ixp33_ASAP7_75t_L g729 ( .A1(n_724), .A2(n_709), .B(n_708), .C(n_705), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_725), .B(n_716), .Y(n_730) );
OAI322xp33_ASAP7_75t_L g731 ( .A1(n_719), .A2(n_707), .A3(n_654), .B1(n_655), .B2(n_684), .C1(n_698), .C2(n_693), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_730), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_727), .A2(n_723), .B1(n_726), .B2(n_720), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_729), .A2(n_689), .B1(n_655), .B2(n_695), .C(n_685), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_732), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_733), .A2(n_728), .B1(n_731), .B2(n_679), .Y(n_736) );
INVx2_ASAP7_75t_SL g737 ( .A(n_735), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_736), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_734), .B1(n_701), .B2(n_682), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_739), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_740), .A2(n_737), .B(n_679), .Y(n_741) );
endmodule