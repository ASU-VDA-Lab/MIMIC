module fake_jpeg_12210_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_61),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_0),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_77),
.B1(n_84),
.B2(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_76),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_19),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_54),
.B1(n_60),
.B2(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_94),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_55),
.B(n_59),
.C(n_70),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_100),
.B(n_25),
.Y(n_120)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_69),
.C(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_56),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_5),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_50),
.B1(n_48),
.B2(n_4),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_1),
.B(n_2),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_112),
.B1(n_27),
.B2(n_28),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_118),
.B1(n_32),
.B2(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_114),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_15),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_30),
.C(n_31),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_129),
.C(n_107),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_35),
.C(n_42),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_114),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_127),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_123),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_139),
.B1(n_123),
.B2(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_131),
.C(n_129),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_138),
.B(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_103),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_136),
.B1(n_104),
.B2(n_117),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_146),
.Y(n_147)
);


endmodule