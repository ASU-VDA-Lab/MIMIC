module real_jpeg_31059_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_0),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_7),
.B1(n_15),
.B2(n_18),
.Y(n_14)
);

CKINVDCx11_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_73),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_2),
.A2(n_73),
.B1(n_259),
.B2(n_263),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_5),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_6),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_6),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_77),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22x1_ASAP7_75t_SL g199 ( 
.A1(n_8),
.A2(n_77),
.B1(n_200),
.B2(n_204),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_8),
.B(n_227),
.Y(n_226)
);

AOI22x1_ASAP7_75t_SL g270 ( 
.A1(n_8),
.A2(n_77),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

OAI32xp33_ASAP7_75t_L g285 ( 
.A1(n_8),
.A2(n_286),
.A3(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_8),
.B(n_210),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_55),
.B1(n_120),
.B2(n_166),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_55),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g311 ( 
.A1(n_10),
.A2(n_55),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_12),
.Y(n_178)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_251),
.Y(n_18)
);

NAND2xp33_ASAP7_75t_R g19 ( 
.A(n_20),
.B(n_247),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_212),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_21),
.B(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_149),
.Y(n_21)
);

XOR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_110),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_76),
.C(n_86),
.Y(n_23)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_24),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_64),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_54),
.Y(n_25)
);

NAND2x1_ASAP7_75t_L g208 ( 
.A(n_26),
.B(n_68),
.Y(n_208)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_27),
.B(n_270),
.Y(n_269)
);

AO21x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_35),
.B(n_44),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_47),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_51),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_54),
.B(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_61),
.Y(n_273)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_67),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_72),
.Y(n_272)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_76),
.A2(n_86),
.B1(n_87),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_76),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_76),
.A2(n_86),
.B1(n_87),
.B2(n_216),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_77),
.A2(n_133),
.B(n_153),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g220 ( 
.A1(n_77),
.A2(n_221),
.A3(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_77),
.B(n_287),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_R g332 ( 
.A(n_77),
.B(n_188),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_77),
.B(n_90),
.Y(n_341)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2x1p5_ASAP7_75t_L g155 ( 
.A(n_79),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_79),
.B(n_165),
.Y(n_164)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_99),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_88),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_89),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_89),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_93),
.Y(n_314)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_94),
.Y(n_313)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_94),
.Y(n_340)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_95),
.B(n_307),
.Y(n_306)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_100),
.B(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_136),
.Y(n_110)
);

OAI31xp33_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.A3(n_119),
.B(n_124),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_129),
.B(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_142),
.B(n_148),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_141),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_148),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_171),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_206),
.B1(n_207),
.B2(n_211),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_172),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_198),
.B(n_199),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_173),
.B(n_199),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_188),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_182),
.B2(n_184),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_181),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_194),
.B2(n_197),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_240),
.Y(n_266)
);

NAND2x1p5_ASAP7_75t_L g318 ( 
.A(n_198),
.B(n_258),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_238),
.Y(n_237)
);

BUFx4f_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2x1p5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_219),
.C(n_236),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_213),
.B(n_279),
.Y(n_278)
);

OAI22x1_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_214),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_236),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_231),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_220),
.A2(n_231),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_231),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_234),
.B(n_235),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_239),
.B(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_280),
.B(n_352),
.Y(n_252)
);

NOR2xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_278),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_254),
.B(n_278),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_267),
.C(n_274),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_256),
.B(n_267),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.Y(n_256)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_303),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_350),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_345),
.B(n_351),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_321),
.B(n_344),
.Y(n_281)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_304),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_304),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_301),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_285),
.B1(n_301),
.B2(n_302),
.Y(n_323)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_315),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

AND2x4_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_347),
.C(n_348),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_330),
.B(n_343),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_324),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI21x1_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_334),
.B(n_342),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_333),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_337),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_349),
.Y(n_351)
);


endmodule