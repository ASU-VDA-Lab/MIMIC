module real_aes_913_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g206 ( .A(n_0), .B(n_153), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_1), .B(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_2), .B(n_137), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_3), .B(n_155), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_4), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g144 ( .A(n_5), .Y(n_144) );
NAND2xp33_ASAP7_75t_SL g250 ( .A(n_6), .B(n_143), .Y(n_250) );
INVx1_ASAP7_75t_L g242 ( .A(n_7), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_8), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_9), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g131 ( .A(n_10), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g476 ( .A(n_11), .B(n_248), .Y(n_476) );
AND2x2_ASAP7_75t_L g540 ( .A(n_12), .B(n_182), .Y(n_540) );
INVx2_ASAP7_75t_L g133 ( .A(n_13), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_14), .B(n_155), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_15), .Y(n_114) );
NOR3xp33_ASAP7_75t_L g785 ( .A(n_15), .B(n_786), .C(n_788), .Y(n_785) );
AOI221x1_ASAP7_75t_L g245 ( .A1(n_16), .A2(n_146), .B1(n_246), .B2(n_248), .C(n_249), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_17), .B(n_137), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_18), .B(n_137), .Y(n_495) );
INVx1_ASAP7_75t_L g118 ( .A(n_19), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_20), .A2(n_66), .B1(n_442), .B2(n_443), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_20), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_21), .A2(n_93), .B1(n_137), .B2(n_186), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_22), .A2(n_146), .B(n_151), .Y(n_145) );
AOI221xp5_ASAP7_75t_SL g216 ( .A1(n_23), .A2(n_37), .B1(n_137), .B2(n_146), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_24), .B(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g134 ( .A(n_25), .B(n_91), .Y(n_134) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_25), .A2(n_91), .B(n_133), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_26), .B(n_155), .Y(n_233) );
INVxp67_ASAP7_75t_L g244 ( .A(n_27), .Y(n_244) );
AND2x2_ASAP7_75t_L g177 ( .A(n_28), .B(n_167), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_29), .B(n_779), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_30), .A2(n_146), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_31), .A2(n_248), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_32), .B(n_155), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_33), .A2(n_146), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_34), .B(n_155), .Y(n_511) );
AND2x2_ASAP7_75t_L g143 ( .A(n_35), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g147 ( .A(n_35), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g194 ( .A(n_35), .Y(n_194) );
OR2x6_ASAP7_75t_L g116 ( .A(n_36), .B(n_117), .Y(n_116) );
INVxp67_ASAP7_75t_L g788 ( .A(n_36), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_38), .B(n_137), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_39), .A2(n_83), .B1(n_146), .B2(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_40), .B(n_155), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_41), .B(n_137), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_42), .B(n_153), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_43), .A2(n_146), .B(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_44), .A2(n_52), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_44), .Y(n_769) );
AND2x2_ASAP7_75t_L g209 ( .A(n_45), .B(n_167), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_46), .B(n_153), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_47), .B(n_167), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_48), .B(n_137), .Y(n_519) );
INVx1_ASAP7_75t_L g140 ( .A(n_49), .Y(n_140) );
INVx1_ASAP7_75t_L g150 ( .A(n_49), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_50), .A2(n_53), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_50), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_51), .B(n_155), .Y(n_474) );
INVx1_ASAP7_75t_L g768 ( .A(n_52), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_53), .Y(n_122) );
AND2x2_ASAP7_75t_L g486 ( .A(n_53), .B(n_167), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_54), .B(n_137), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_55), .B(n_153), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_56), .B(n_153), .Y(n_510) );
AND2x2_ASAP7_75t_L g168 ( .A(n_57), .B(n_167), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_58), .B(n_137), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_59), .B(n_155), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_60), .B(n_137), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_61), .A2(n_146), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_62), .B(n_153), .Y(n_164) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_63), .B(n_132), .Y(n_234) );
AND2x2_ASAP7_75t_L g501 ( .A(n_64), .B(n_132), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_65), .A2(n_146), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_66), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_67), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_68), .B(n_182), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_69), .B(n_153), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_70), .B(n_153), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_71), .A2(n_95), .B1(n_146), .B2(n_192), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_72), .B(n_155), .Y(n_498) );
INVx1_ASAP7_75t_L g142 ( .A(n_73), .Y(n_142) );
INVx1_ASAP7_75t_L g148 ( .A(n_73), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_74), .B(n_153), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_75), .A2(n_146), .B(n_490), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_76), .A2(n_146), .B(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_77), .A2(n_146), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g513 ( .A(n_78), .B(n_132), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_79), .B(n_167), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_80), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_80), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_81), .B(n_137), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_82), .A2(n_85), .B1(n_137), .B2(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_86), .A2(n_105), .B1(n_781), .B2(n_790), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_87), .B(n_153), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_88), .B(n_153), .Y(n_219) );
AND2x2_ASAP7_75t_L g467 ( .A(n_89), .B(n_182), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_90), .A2(n_146), .B(n_162), .Y(n_161) );
XNOR2xp5_ASAP7_75t_L g763 ( .A(n_92), .B(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_94), .B(n_155), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_96), .A2(n_146), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_97), .B(n_155), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_98), .B(n_137), .Y(n_208) );
INVxp67_ASAP7_75t_L g247 ( .A(n_99), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_100), .B(n_155), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_101), .A2(n_146), .B(n_231), .Y(n_230) );
BUFx2_ASAP7_75t_L g500 ( .A(n_102), .Y(n_500) );
BUFx2_ASAP7_75t_L g109 ( .A(n_103), .Y(n_109) );
BUFx2_ASAP7_75t_SL g777 ( .A(n_103), .Y(n_777) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B(n_448), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_107), .A2(n_444), .B1(n_776), .B2(n_778), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_109), .B(n_116), .Y(n_770) );
OAI21x1_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_120), .B(n_444), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g447 ( .A(n_113), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_114), .Y(n_451) );
OR2x2_ASAP7_75t_L g780 ( .A(n_114), .B(n_116), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_118), .B(n_119), .Y(n_789) );
XOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
XNOR2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_441), .Y(n_124) );
INVx3_ASAP7_75t_SL g760 ( .A(n_125), .Y(n_760) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_371), .Y(n_125) );
NOR4xp25_ASAP7_75t_SL g126 ( .A(n_127), .B(n_264), .C(n_308), .D(n_335), .Y(n_126) );
OAI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_225), .B1(n_235), .B2(n_252), .C(n_254), .Y(n_127) );
AOI32xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_178), .A3(n_198), .B1(n_210), .B2(n_221), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_129), .B(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_129), .A2(n_377), .B1(n_435), .B2(n_438), .Y(n_434) );
AND2x4_ASAP7_75t_SL g129 ( .A(n_130), .B(n_158), .Y(n_129) );
INVx5_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
OR2x2_ASAP7_75t_L g253 ( .A(n_130), .B(n_223), .Y(n_253) );
AND2x4_ASAP7_75t_L g255 ( .A(n_130), .B(n_170), .Y(n_255) );
INVx2_ASAP7_75t_L g270 ( .A(n_130), .Y(n_270) );
OR2x2_ASAP7_75t_L g282 ( .A(n_130), .B(n_179), .Y(n_282) );
AND2x2_ASAP7_75t_L g289 ( .A(n_130), .B(n_169), .Y(n_289) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_130), .B(n_212), .Y(n_331) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_130), .Y(n_388) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x4_ASAP7_75t_L g157 ( .A(n_133), .B(n_134), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_145), .B(n_157), .Y(n_135) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
INVx1_ASAP7_75t_L g251 ( .A(n_138), .Y(n_251) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
AND2x6_ASAP7_75t_L g153 ( .A(n_139), .B(n_148), .Y(n_153) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g155 ( .A(n_141), .B(n_150), .Y(n_155) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx5_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
AND2x2_ASAP7_75t_L g149 ( .A(n_144), .B(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
BUFx3_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
INVx2_ASAP7_75t_L g196 ( .A(n_148), .Y(n_196) );
AND2x4_ASAP7_75t_L g192 ( .A(n_149), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B(n_156), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_153), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_156), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_156), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_156), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_156), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_156), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_156), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_156), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_156), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_156), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_156), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_156), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_156), .A2(n_537), .B(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_157), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_157), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_157), .B(n_247), .Y(n_246) );
NOR3xp33_ASAP7_75t_L g249 ( .A(n_157), .B(n_250), .C(n_251), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_157), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_157), .A2(n_519), .B(n_520), .Y(n_518) );
INVx3_ASAP7_75t_SL g283 ( .A(n_158), .Y(n_283) );
AND2x2_ASAP7_75t_L g302 ( .A(n_158), .B(n_224), .Y(n_302) );
AOI32xp33_ASAP7_75t_L g417 ( .A1(n_158), .A2(n_288), .A3(n_318), .B1(n_348), .B2(n_383), .Y(n_417) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_169), .Y(n_158) );
AND2x2_ASAP7_75t_L g257 ( .A(n_159), .B(n_179), .Y(n_257) );
OR2x2_ASAP7_75t_L g273 ( .A(n_159), .B(n_170), .Y(n_273) );
INVx1_ASAP7_75t_L g296 ( .A(n_159), .Y(n_296) );
INVx2_ASAP7_75t_L g312 ( .A(n_159), .Y(n_312) );
AND2x2_ASAP7_75t_L g349 ( .A(n_159), .B(n_212), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_159), .B(n_170), .Y(n_368) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_159), .Y(n_437) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_166), .B(n_168), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_165), .Y(n_160) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_166), .A2(n_171), .B(n_177), .Y(n_170) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_171), .B(n_177), .Y(n_223) );
AOI21x1_ASAP7_75t_L g533 ( .A1(n_166), .A2(n_534), .B(n_540), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_167), .Y(n_166) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_167), .A2(n_216), .B(n_220), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_167), .A2(n_462), .B(n_463), .Y(n_461) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_167), .A2(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g404 ( .A(n_170), .B(n_179), .Y(n_404) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_170), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_176), .Y(n_171) );
OR2x2_ASAP7_75t_L g252 ( .A(n_178), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g258 ( .A(n_178), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g271 ( .A(n_178), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g433 ( .A(n_178), .B(n_302), .Y(n_433) );
BUFx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g362 ( .A(n_179), .B(n_312), .Y(n_362) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_180), .Y(n_212) );
AOI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B(n_197), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_182), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_182), .A2(n_495), .B(n_496), .Y(n_494) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g202 ( .A(n_183), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_191), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_186), .A2(n_192), .B1(n_241), .B2(n_243), .Y(n_240) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_190), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2x1p5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_198), .B(n_329), .Y(n_431) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_199), .B(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g214 ( .A(n_200), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
AND2x2_ASAP7_75t_L g262 ( .A(n_200), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_200), .B(n_238), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_200), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g320 ( .A(n_200), .Y(n_320) );
OR2x2_ASAP7_75t_L g339 ( .A(n_200), .B(n_266), .Y(n_339) );
INVx1_ASAP7_75t_L g346 ( .A(n_200), .Y(n_346) );
NOR2xp33_ASAP7_75t_R g398 ( .A(n_200), .B(n_227), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_200), .B(n_239), .Y(n_402) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AOI21x1_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_209), .Y(n_201) );
INVx4_ASAP7_75t_L g248 ( .A(n_202), .Y(n_248) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_202), .A2(n_470), .B(n_476), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_208), .Y(n_203) );
AOI32xp33_ASAP7_75t_L g425 ( .A1(n_210), .A2(n_261), .A3(n_426), .B1(n_427), .B2(n_428), .Y(n_425) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g292 ( .A(n_212), .Y(n_292) );
AND2x4_ASAP7_75t_L g311 ( .A(n_212), .B(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_212), .B(n_283), .Y(n_340) );
OR2x2_ASAP7_75t_L g394 ( .A(n_212), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g352 ( .A(n_213), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g410 ( .A(n_213), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_214), .B(n_227), .Y(n_376) );
AND2x2_ASAP7_75t_L g413 ( .A(n_214), .B(n_379), .Y(n_413) );
INVx2_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
INVx2_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_215), .B(n_227), .Y(n_286) );
INVx1_ASAP7_75t_L g317 ( .A(n_215), .Y(n_317) );
OR2x2_ASAP7_75t_L g343 ( .A(n_215), .B(n_227), .Y(n_343) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_215), .Y(n_395) );
BUFx3_ASAP7_75t_L g424 ( .A(n_215), .Y(n_424) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_222), .B(n_311), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_222), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_223), .B(n_296), .Y(n_295) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_223), .A2(n_292), .B(n_310), .Y(n_325) );
OAI32xp33_ASAP7_75t_L g347 ( .A1(n_224), .A2(n_348), .A3(n_350), .B1(n_352), .B2(n_354), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_224), .B(n_311), .Y(n_420) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g353 ( .A(n_226), .Y(n_353) );
NOR2x1p5_ASAP7_75t_L g423 ( .A(n_226), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x4_ASAP7_75t_L g237 ( .A(n_227), .B(n_238), .Y(n_237) );
AND2x4_ASAP7_75t_SL g261 ( .A(n_227), .B(n_239), .Y(n_261) );
OR2x2_ASAP7_75t_L g265 ( .A(n_227), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_227), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g329 ( .A(n_227), .B(n_239), .Y(n_329) );
OR2x2_ASAP7_75t_L g391 ( .A(n_227), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g408 ( .A(n_227), .B(n_339), .Y(n_408) );
INVx1_ASAP7_75t_L g440 ( .A(n_227), .Y(n_440) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_236), .B(n_317), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_237), .B(n_351), .Y(n_350) );
AOI222xp33_ASAP7_75t_L g355 ( .A1(n_237), .A2(n_356), .B1(n_361), .B2(n_363), .C1(n_366), .C2(n_369), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_237), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g383 ( .A(n_237), .B(n_262), .Y(n_383) );
AND2x2_ASAP7_75t_L g345 ( .A(n_238), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g360 ( .A(n_238), .B(n_265), .Y(n_360) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_239), .B(n_266), .Y(n_298) );
AND2x4_ASAP7_75t_L g319 ( .A(n_239), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g379 ( .A(n_239), .B(n_300), .Y(n_379) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_245), .Y(n_239) );
INVx3_ASAP7_75t_L g506 ( .A(n_248), .Y(n_506) );
INVx1_ASAP7_75t_SL g259 ( .A(n_253), .Y(n_259) );
NAND2xp33_ASAP7_75t_SL g428 ( .A(n_253), .B(n_283), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_258), .C(n_260), .Y(n_254) );
INVx2_ASAP7_75t_SL g305 ( .A(n_255), .Y(n_305) );
AND2x2_ASAP7_75t_L g309 ( .A(n_256), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_257), .B(n_305), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_257), .A2(n_295), .B(n_331), .C(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g407 ( .A(n_257), .B(n_388), .Y(n_407) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x4_ASAP7_75t_L g306 ( .A(n_261), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g411 ( .A(n_261), .Y(n_411) );
OAI211xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B(n_274), .C(n_301), .Y(n_264) );
INVx2_ASAP7_75t_L g276 ( .A(n_265), .Y(n_276) );
OR2x2_ASAP7_75t_L g323 ( .A(n_265), .B(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_269), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g361 ( .A(n_269), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_269), .B(n_349), .Y(n_415) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_271), .A2(n_374), .B1(n_375), .B2(n_377), .C1(n_380), .C2(n_383), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_272), .A2(n_337), .B1(n_340), .B2(n_341), .C(n_347), .Y(n_336) );
AND2x2_ASAP7_75t_L g374 ( .A(n_272), .B(n_331), .Y(n_374) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp33_ASAP7_75t_SL g287 ( .A(n_273), .B(n_288), .Y(n_287) );
AOI221x1_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B1(n_284), .B2(n_287), .C(n_290), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g427 ( .A(n_277), .B(n_365), .Y(n_427) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g285 ( .A(n_278), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OAI32xp33_ASAP7_75t_L g393 ( .A1(n_283), .A2(n_324), .A3(n_394), .B1(n_396), .B2(n_400), .Y(n_393) );
OAI21xp33_ASAP7_75t_SL g412 ( .A1(n_284), .A2(n_413), .B(n_414), .Y(n_412) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI21xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_294), .B(n_297), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OR2x2_ASAP7_75t_L g294 ( .A(n_292), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g367 ( .A(n_292), .B(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_296), .A2(n_322), .B1(n_325), .B2(n_326), .C(n_330), .Y(n_321) );
INVx1_ASAP7_75t_L g397 ( .A(n_296), .Y(n_397) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_296), .Y(n_403) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_306), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_305), .B(n_370), .Y(n_369) );
OAI21xp5_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_313), .B(n_321), .Y(n_308) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_312), .Y(n_382) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_315), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g334 ( .A(n_317), .Y(n_334) );
INVx1_ASAP7_75t_L g324 ( .A(n_319), .Y(n_324) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_319), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_319), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_319), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g338 ( .A(n_329), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_334), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_336), .B(n_355), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g351 ( .A(n_339), .Y(n_351) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_SL g365 ( .A(n_343), .Y(n_365) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_345), .B(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_346), .Y(n_359) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_357), .B(n_360), .Y(n_356) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g370 ( .A(n_362), .Y(n_370) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g389 ( .A(n_368), .Y(n_389) );
NOR4xp25_ASAP7_75t_L g371 ( .A(n_372), .B(n_405), .C(n_416), .D(n_429), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_384), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_374), .A2(n_385), .B(n_390), .C(n_393), .Y(n_384) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_387), .B(n_389), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_387), .A2(n_397), .B(n_398), .C(n_399), .Y(n_396) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
OAI21xp33_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_404), .B(n_436), .Y(n_435) );
OAI221xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_408), .B1(n_409), .B2(n_410), .C(n_412), .Y(n_405) );
INVx1_ASAP7_75t_SL g409 ( .A(n_407), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_418), .C(n_425), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp33_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_449), .B(n_773), .Y(n_448) );
AOI32xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_758), .A3(n_761), .B1(n_771), .B2(n_772), .Y(n_449) );
INVx1_ASAP7_75t_L g771 ( .A(n_450), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_451), .Y(n_759) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_683), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_455), .B(n_602), .Y(n_454) );
NAND5xp2_ASAP7_75t_L g455 ( .A(n_456), .B(n_546), .C(n_556), .D(n_573), .E(n_589), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_482), .B1(n_524), .B2(n_528), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_468), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g530 ( .A(n_460), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g548 ( .A(n_460), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g569 ( .A(n_460), .B(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g583 ( .A(n_460), .Y(n_583) );
AND2x2_ASAP7_75t_L g592 ( .A(n_460), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_SL g614 ( .A(n_460), .B(n_532), .Y(n_614) );
BUFx2_ASAP7_75t_L g657 ( .A(n_460), .Y(n_657) );
AND2x2_ASAP7_75t_L g672 ( .A(n_460), .B(n_469), .Y(n_672) );
OR2x2_ASAP7_75t_L g704 ( .A(n_460), .B(n_705), .Y(n_704) );
NOR4xp25_ASAP7_75t_L g753 ( .A(n_460), .B(n_754), .C(n_755), .D(n_756), .Y(n_753) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_467), .Y(n_460) );
AOI31xp33_ASAP7_75t_L g621 ( .A1(n_468), .A2(n_622), .A3(n_624), .B(n_626), .Y(n_621) );
INVx2_ASAP7_75t_SL g738 ( .A(n_468), .Y(n_738) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
INVx2_ASAP7_75t_L g545 ( .A(n_469), .Y(n_545) );
AND2x2_ASAP7_75t_L g549 ( .A(n_469), .B(n_533), .Y(n_549) );
INVx2_ASAP7_75t_L g572 ( .A(n_469), .Y(n_572) );
AND2x2_ASAP7_75t_L g591 ( .A(n_469), .B(n_532), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g550 ( .A(n_477), .Y(n_550) );
INVx2_ASAP7_75t_L g568 ( .A(n_477), .Y(n_568) );
AND2x2_ASAP7_75t_L g623 ( .A(n_477), .B(n_583), .Y(n_623) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AND2x4_ASAP7_75t_L g594 ( .A(n_478), .B(n_479), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_514), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_502), .Y(n_483) );
OR2x2_ASAP7_75t_L g524 ( .A(n_484), .B(n_525), .Y(n_524) );
INVx3_ASAP7_75t_L g675 ( .A(n_484), .Y(n_675) );
OR2x2_ASAP7_75t_L g723 ( .A(n_484), .B(n_724), .Y(n_723) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
OR2x2_ASAP7_75t_SL g515 ( .A(n_485), .B(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g553 ( .A(n_485), .Y(n_553) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_485), .Y(n_597) );
INVx2_ASAP7_75t_L g605 ( .A(n_485), .Y(n_605) );
OR2x2_ASAP7_75t_L g640 ( .A(n_485), .B(n_504), .Y(n_640) );
AND2x2_ASAP7_75t_L g752 ( .A(n_485), .B(n_607), .Y(n_752) );
AND2x2_ASAP7_75t_L g757 ( .A(n_485), .B(n_517), .Y(n_757) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OR2x2_ASAP7_75t_L g516 ( .A(n_493), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g581 ( .A(n_493), .B(n_503), .Y(n_581) );
OR2x2_ASAP7_75t_L g588 ( .A(n_493), .B(n_553), .Y(n_588) );
NOR2x1_ASAP7_75t_SL g607 ( .A(n_493), .B(n_527), .Y(n_607) );
BUFx2_ASAP7_75t_L g639 ( .A(n_493), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_493), .B(n_553), .Y(n_648) );
AND2x2_ASAP7_75t_L g681 ( .A(n_493), .B(n_601), .Y(n_681) );
INVx2_ASAP7_75t_SL g690 ( .A(n_493), .Y(n_690) );
AND2x2_ASAP7_75t_L g693 ( .A(n_493), .B(n_504), .Y(n_693) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_501), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_502), .B(n_558), .C(n_643), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_502), .B(n_605), .Y(n_708) );
INVxp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_503), .B(n_690), .Y(n_711) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_504), .Y(n_555) );
AND2x2_ASAP7_75t_L g599 ( .A(n_504), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g664 ( .A(n_504), .B(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_513), .Y(n_505) );
AO21x1_ASAP7_75t_SL g527 ( .A1(n_506), .A2(n_507), .B(n_513), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AND2x4_ASAP7_75t_L g559 ( .A(n_514), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g695 ( .A(n_516), .B(n_640), .Y(n_695) );
AND2x2_ASAP7_75t_L g526 ( .A(n_517), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g563 ( .A(n_517), .Y(n_563) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_517), .Y(n_580) );
INVx2_ASAP7_75t_L g601 ( .A(n_517), .Y(n_601) );
INVx1_ASAP7_75t_L g665 ( .A(n_517), .Y(n_665) );
INVx2_ASAP7_75t_L g747 ( .A(n_524), .Y(n_747) );
OR2x2_ASAP7_75t_L g611 ( .A(n_525), .B(n_588), .Y(n_611) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g751 ( .A(n_526), .B(n_648), .Y(n_751) );
AND2x2_ASAP7_75t_L g644 ( .A(n_527), .B(n_601), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_541), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_530), .A2(n_658), .B1(n_675), .B2(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g571 ( .A(n_532), .Y(n_571) );
AND2x2_ASAP7_75t_L g625 ( .A(n_532), .B(n_545), .Y(n_625) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_532), .Y(n_652) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_533), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
INVxp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_543), .B(n_657), .Y(n_656) );
OAI32xp33_ASAP7_75t_L g673 ( .A1(n_543), .A2(n_674), .A3(n_676), .B1(n_677), .B2(n_679), .Y(n_673) );
BUFx2_ASAP7_75t_L g558 ( .A(n_544), .Y(n_558) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g700 ( .A(n_545), .B(n_594), .Y(n_700) );
OR4x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .C(n_551), .D(n_554), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_547), .A2(n_638), .B1(n_732), .B2(n_733), .Y(n_731) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_548), .Y(n_740) );
AND2x2_ASAP7_75t_L g582 ( .A(n_549), .B(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g662 ( .A(n_549), .Y(n_662) );
INVx1_ASAP7_75t_L g678 ( .A(n_549), .Y(n_678) );
INVx1_ASAP7_75t_L g713 ( .A(n_549), .Y(n_713) );
OR2x2_ASAP7_75t_L g670 ( .A(n_550), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g714 ( .A(n_550), .B(n_715), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_551), .A2(n_588), .B1(n_632), .B2(n_651), .Y(n_653) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g697 ( .A(n_552), .B(n_606), .Y(n_697) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g579 ( .A(n_553), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g560 ( .A(n_554), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g687 ( .A(n_554), .B(n_558), .C(n_639), .D(n_651), .Y(n_687) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g724 ( .A(n_555), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B1(n_561), .B2(n_565), .Y(n_556) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_557), .A2(n_558), .B1(n_708), .B2(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx3_ASAP7_75t_L g586 ( .A(n_563), .Y(n_586) );
AOI32xp33_ASAP7_75t_L g702 ( .A1(n_563), .A2(n_703), .A3(n_707), .B1(n_712), .B2(n_716), .Y(n_702) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_566), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g661 ( .A(n_566), .B(n_662), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_566), .A2(n_574), .B1(n_686), .B2(n_691), .C(n_694), .Y(n_685) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g618 ( .A(n_567), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g733 ( .A(n_567), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_568), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g575 ( .A(n_570), .Y(n_575) );
AND2x2_ASAP7_75t_L g593 ( .A(n_570), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_SL g633 ( .A(n_571), .Y(n_633) );
INVx1_ASAP7_75t_L g617 ( .A(n_572), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B1(n_582), .B2(n_584), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g719 ( .A(n_575), .B(n_649), .Y(n_719) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g659 ( .A(n_578), .Y(n_659) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g590 ( .A(n_583), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_583), .B(n_620), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_583), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_583), .B(n_625), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_584), .A2(n_744), .B1(n_745), .B2(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
OR2x2_ASAP7_75t_L g626 ( .A(n_586), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g636 ( .A(n_586), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_586), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_586), .B(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_SL g691 ( .A(n_586), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g667 ( .A(n_588), .B(n_668), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_595), .Y(n_589) );
INVx1_ASAP7_75t_L g609 ( .A(n_591), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_592), .A2(n_629), .B1(n_636), .B2(n_641), .Y(n_628) );
INVx3_ASAP7_75t_L g631 ( .A(n_594), .Y(n_631) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
OAI32xp33_ASAP7_75t_SL g686 ( .A1(n_597), .A2(n_657), .A3(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g606 ( .A(n_600), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND4xp25_ASAP7_75t_SL g602 ( .A(n_603), .B(n_628), .C(n_645), .D(n_660), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B1(n_610), .B2(n_612), .C(n_621), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx2_ASAP7_75t_L g643 ( .A(n_605), .Y(n_643) );
AND2x2_ASAP7_75t_L g692 ( .A(n_605), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_605), .B(n_644), .Y(n_730) );
AND2x2_ASAP7_75t_L g741 ( .A(n_605), .B(n_664), .Y(n_741) );
INVx2_ASAP7_75t_L g627 ( .A(n_607), .Y(n_627) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_618), .Y(n_612) );
AND2x2_ASAP7_75t_L g744 ( .A(n_613), .B(n_615), .Y(n_744) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_614), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g721 ( .A(n_619), .Y(n_721) );
INVx1_ASAP7_75t_L g706 ( .A(n_620), .Y(n_706) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_623), .B(n_678), .Y(n_677) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_624), .B(n_631), .Y(n_635) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g734 ( .A(n_625), .Y(n_734) );
INVx1_ASAP7_75t_L g716 ( .A(n_627), .Y(n_716) );
OR2x2_ASAP7_75t_L g732 ( .A(n_627), .B(n_643), .Y(n_732) );
NAND2xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_634), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g649 ( .A(n_631), .Y(n_649) );
AND2x2_ASAP7_75t_L g654 ( .A(n_631), .B(n_644), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_631), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g728 ( .A(n_632), .Y(n_728) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_637), .A2(n_718), .B1(n_720), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g682 ( .A(n_640), .Y(n_682) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g668 ( .A(n_644), .Y(n_668) );
AOI322xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .A3(n_650), .B1(n_653), .B2(n_654), .C1(n_655), .C2(n_658), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_646), .A2(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_648), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g720 ( .A(n_649), .B(n_721), .Y(n_720) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_656), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g676 ( .A(n_657), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_657), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B1(n_666), .B2(n_669), .C(n_673), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_662), .A2(n_749), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_664), .B(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g715 ( .A(n_665), .Y(n_715) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_669), .A2(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp33_ASAP7_75t_SL g749 ( .A(n_678), .B(n_750), .Y(n_749) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NOR4xp75_ASAP7_75t_L g683 ( .A(n_684), .B(n_701), .C(n_725), .D(n_742), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_696), .Y(n_684) );
INVx1_ASAP7_75t_L g755 ( .A(n_693), .Y(n_755) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g727 ( .A(n_700), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g754 ( .A(n_700), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_717), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g750 ( .A(n_721), .Y(n_750) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND3x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_735), .C(n_739), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B(n_731), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_748), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g774 ( .A(n_758), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_770), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_763), .B(n_770), .Y(n_772) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_772), .A2(n_774), .B(n_775), .Y(n_773) );
CKINVDCx8_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_783), .Y(n_790) );
INVx3_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_785), .B(n_789), .Y(n_784) );
endmodule