module fake_jpeg_2660_n_570 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_570);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_570;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_17),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_55),
.Y(n_158)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_60),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_0),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_66),
.Y(n_115)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_72),
.Y(n_130)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_75),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_28),
.B(n_10),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_28),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_76),
.B(n_82),
.Y(n_150)
);

INVx2_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_77),
.B(n_29),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_32),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_8),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_23),
.B(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_87),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_51),
.Y(n_148)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_1),
.Y(n_159)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_49),
.B1(n_22),
.B2(n_51),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_112),
.A2(n_126),
.B1(n_47),
.B2(n_30),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_60),
.A2(n_49),
.B1(n_22),
.B2(n_51),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_29),
.B1(n_49),
.B2(n_43),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_138),
.B1(n_165),
.B2(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_42),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_136),
.B(n_155),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_29),
.B1(n_46),
.B2(n_51),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_152),
.B1(n_169),
.B2(n_170),
.Y(n_178)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_163),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_29),
.B1(n_36),
.B2(n_42),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_70),
.B(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_69),
.B(n_52),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_157),
.B(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_121),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_23),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_97),
.Y(n_187)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_68),
.A2(n_36),
.B1(n_24),
.B2(n_27),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_85),
.A2(n_46),
.B1(n_40),
.B2(n_32),
.Y(n_170)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_172),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_179),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_43),
.B1(n_24),
.B2(n_78),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_174),
.A2(n_125),
.B1(n_134),
.B2(n_119),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_176),
.A2(n_181),
.B1(n_184),
.B2(n_198),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_108),
.A2(n_88),
.A3(n_96),
.B1(n_77),
.B2(n_100),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_150),
.B1(n_169),
.B2(n_112),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_126),
.A2(n_80),
.B1(n_98),
.B2(n_104),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_190),
.B(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_110),
.A2(n_73),
.B1(n_71),
.B2(n_65),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_97),
.B1(n_93),
.B2(n_101),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_185),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_115),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_186),
.B(n_189),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_187),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_111),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_128),
.A2(n_55),
.B(n_103),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_130),
.A2(n_56),
.B1(n_94),
.B2(n_59),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_193),
.A2(n_228),
.B1(n_230),
.B2(n_135),
.Y(n_242)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

BUFx24_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_89),
.B1(n_95),
.B2(n_74),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_197),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_131),
.A2(n_83),
.B(n_61),
.C(n_30),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_200),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_124),
.B(n_109),
.C(n_113),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_209),
.C(n_217),
.Y(n_234)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

BUFx2_ASAP7_75t_SL g251 ( 
.A(n_202),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_116),
.A2(n_65),
.B1(n_71),
.B2(n_51),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_203),
.A2(n_205),
.B1(n_208),
.B2(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_116),
.A2(n_40),
.B1(n_32),
.B2(n_46),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_40),
.B1(n_32),
.B2(n_46),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_40),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_117),
.B(n_32),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_213),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_129),
.A2(n_30),
.B1(n_25),
.B2(n_50),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_120),
.B(n_40),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_137),
.Y(n_215)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_111),
.B(n_2),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_142),
.B(n_83),
.C(n_61),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_219),
.C(n_223),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_146),
.B(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_114),
.A2(n_30),
.B1(n_25),
.B2(n_4),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_144),
.B(n_2),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_5),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_30),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_120),
.B(n_2),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_225),
.A2(n_7),
.B(n_11),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_227),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_167),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_232),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_167),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_134),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_139),
.B1(n_156),
.B2(n_119),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_235),
.A2(n_252),
.B1(n_253),
.B2(n_262),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_238),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_156),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_250),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_127),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_243),
.B(n_279),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_195),
.B(n_127),
.CI(n_135),
.CON(n_250),
.SN(n_250)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_183),
.A2(n_160),
.B1(n_107),
.B2(n_140),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_140),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_271),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_178),
.A2(n_160),
.B1(n_107),
.B2(n_11),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_178),
.A2(n_5),
.B1(n_7),
.B2(n_11),
.Y(n_267)
);

AO21x2_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_283),
.B(n_284),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_268),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_178),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_270),
.B1(n_208),
.B2(n_229),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_178),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_7),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_182),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_196),
.B1(n_175),
.B2(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_171),
.B(n_217),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_281),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_228),
.B(n_187),
.C(n_185),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_217),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_188),
.B(n_192),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_191),
.C(n_218),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_15),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_212),
.A2(n_190),
.B1(n_185),
.B2(n_197),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_185),
.A2(n_18),
.B1(n_197),
.B2(n_182),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g285 ( 
.A(n_206),
.B(n_200),
.C(n_197),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_287),
.C(n_209),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_188),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_310),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_239),
.B(n_173),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_290),
.B(n_294),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_184),
.B1(n_187),
.B2(n_210),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_291),
.A2(n_338),
.B(n_298),
.Y(n_367)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_263),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_292),
.B(n_295),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_263),
.B(n_180),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_233),
.A2(n_194),
.B(n_172),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_296),
.A2(n_253),
.B(n_277),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_247),
.A2(n_209),
.B1(n_199),
.B2(n_226),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_302),
.B1(n_309),
.B2(n_314),
.Y(n_339)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_247),
.A2(n_199),
.B1(n_216),
.B2(n_227),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_303),
.B(n_318),
.Y(n_372)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_308),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_175),
.B1(n_214),
.B2(n_207),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_258),
.A2(n_177),
.B1(n_207),
.B2(n_204),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_249),
.Y(n_316)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_239),
.B(n_275),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_317),
.B(n_319),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_255),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_282),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_237),
.B(n_177),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_323),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_265),
.Y(n_321)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_258),
.A2(n_224),
.B1(n_231),
.B2(n_232),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_322),
.A2(n_326),
.B1(n_335),
.B2(n_244),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_238),
.B(n_202),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_327),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_261),
.A2(n_280),
.B1(n_242),
.B2(n_264),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_243),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_267),
.B1(n_270),
.B2(n_269),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_329),
.A2(n_268),
.B1(n_278),
.B2(n_250),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_234),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_330),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_266),
.B(n_234),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_332),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_254),
.B(n_286),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_236),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_333),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_260),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_337),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_264),
.A2(n_287),
.B1(n_285),
.B2(n_262),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_SL g336 ( 
.A(n_233),
.B(n_250),
.C(n_257),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_336),
.Y(n_381)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_279),
.C(n_260),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_340),
.B(n_344),
.C(n_349),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_368),
.B(n_377),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_307),
.B(n_256),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_351),
.B1(n_289),
.B2(n_308),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_342),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_286),
.C(n_236),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_300),
.A2(n_235),
.B1(n_259),
.B2(n_273),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_300),
.A2(n_252),
.B1(n_273),
.B2(n_240),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_352),
.A2(n_358),
.B1(n_371),
.B2(n_374),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_274),
.B(n_241),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_354),
.B(n_375),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_241),
.C(n_276),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_362),
.C(n_364),
.Y(n_399)
);

OA22x2_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_251),
.B1(n_265),
.B2(n_298),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_351),
.B(n_341),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_300),
.A2(n_251),
.B1(n_265),
.B2(n_335),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_265),
.C(n_313),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_315),
.Y(n_364)
);

AO21x2_ASAP7_75t_L g418 ( 
.A1(n_367),
.A2(n_368),
.B(n_357),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_297),
.A2(n_296),
.B(n_293),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_300),
.A2(n_326),
.B1(n_299),
.B2(n_302),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_329),
.A2(n_314),
.B1(n_322),
.B2(n_310),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_293),
.A2(n_289),
.B(n_303),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_289),
.A2(n_315),
.B(n_316),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_309),
.A2(n_289),
.B1(n_306),
.B2(n_320),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_378),
.A2(n_306),
.B1(n_312),
.B2(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_319),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_386),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_383),
.B(n_318),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_387),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_323),
.Y(n_389)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_376),
.B1(n_379),
.B2(n_362),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_305),
.Y(n_391)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_356),
.B(n_328),
.Y(n_392)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_392),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_372),
.A2(n_321),
.B1(n_337),
.B2(n_311),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_393),
.A2(n_394),
.B1(n_401),
.B2(n_402),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_397),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_338),
.C(n_301),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_409),
.C(n_349),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_371),
.A2(n_321),
.B1(n_358),
.B2(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_382),
.B(n_363),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_342),
.A2(n_352),
.B1(n_374),
.B2(n_348),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_404),
.B1(n_405),
.B2(n_414),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_410),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_366),
.C(n_355),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_361),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_347),
.A2(n_369),
.B1(n_365),
.B2(n_381),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_411),
.B(n_413),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_359),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_354),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_360),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_415),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_440)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_375),
.A2(n_377),
.B1(n_369),
.B2(n_365),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_364),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_419),
.A2(n_420),
.B1(n_384),
.B2(n_385),
.Y(n_449)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_356),
.B(n_350),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_421),
.B(n_390),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_394),
.A2(n_381),
.B1(n_339),
.B2(n_367),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_429),
.C(n_432),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_411),
.A2(n_339),
.B1(n_357),
.B2(n_350),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_449),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_427),
.A2(n_444),
.B1(n_446),
.B2(n_439),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_379),
.C(n_357),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_373),
.C(n_380),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_373),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_436),
.C(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_380),
.C(n_409),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_419),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_389),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_388),
.A2(n_401),
.B1(n_403),
.B2(n_404),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_388),
.A2(n_404),
.B1(n_414),
.B2(n_408),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_417),
.C(n_412),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_451),
.C(n_420),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_408),
.C(n_395),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_452),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_395),
.B(n_391),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_454),
.B(n_443),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_456),
.B(n_475),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_410),
.Y(n_458)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_415),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_460),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_424),
.B(n_413),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_450),
.A2(n_418),
.B(n_406),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_462),
.A2(n_479),
.B(n_444),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_428),
.B(n_397),
.C(n_407),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_477),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g466 ( 
.A(n_451),
.B(n_418),
.CI(n_416),
.CON(n_466),
.SN(n_466)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_426),
.B(n_422),
.C(n_437),
.Y(n_504)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_457),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_471),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_418),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_470),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_418),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_418),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_474),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_423),
.C(n_432),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_436),
.C(n_441),
.Y(n_489)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_445),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_476),
.Y(n_484)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_425),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_481),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_438),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_450),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_482),
.B(n_461),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_462),
.A2(n_450),
.B(n_446),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_486),
.A2(n_496),
.B(n_471),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_499),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_475),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_429),
.C(n_448),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_498),
.C(n_468),
.Y(n_508)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_494),
.Y(n_507)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

BUFx12f_ASAP7_75t_SL g496 ( 
.A(n_477),
.Y(n_496)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_497),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_427),
.C(n_454),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_430),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_464),
.B(n_452),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_502),
.B(n_459),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_504),
.A2(n_472),
.B(n_481),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_514),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_516),
.Y(n_526)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_487),
.Y(n_511)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_521),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_513),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_500),
.A2(n_479),
.B1(n_465),
.B2(n_482),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_459),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_523),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_485),
.A2(n_455),
.B1(n_465),
.B2(n_476),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_519),
.A2(n_520),
.B1(n_525),
.B2(n_484),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_455),
.B1(n_458),
.B2(n_460),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_474),
.Y(n_521)
);

AO22x1_ASAP7_75t_L g522 ( 
.A1(n_483),
.A2(n_460),
.B1(n_466),
.B2(n_470),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_504),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_489),
.B(n_456),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_521),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_483),
.B(n_467),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_507),
.A2(n_486),
.B1(n_491),
.B2(n_506),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_531),
.B(n_534),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_532),
.A2(n_522),
.B(n_516),
.Y(n_545)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_533),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_488),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_510),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_535),
.A2(n_539),
.B(n_518),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_499),
.C(n_490),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_498),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_524),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_508),
.B(n_484),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_507),
.A2(n_522),
.B1(n_506),
.B2(n_525),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_540),
.A2(n_491),
.B1(n_501),
.B2(n_466),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_542),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_515),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_545),
.A2(n_549),
.B1(n_531),
.B2(n_538),
.Y(n_552)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_546),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_537),
.A2(n_496),
.B(n_514),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_547),
.A2(n_548),
.B(n_550),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_505),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_532),
.A2(n_501),
.B(n_494),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_551),
.A2(n_528),
.B(n_530),
.Y(n_558)
);

AO21x1_ASAP7_75t_L g560 ( 
.A1(n_552),
.A2(n_556),
.B(n_530),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_544),
.A2(n_526),
.B(n_540),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_553),
.A2(n_545),
.B(n_546),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_529),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_558),
.A2(n_550),
.B(n_512),
.Y(n_562)
);

OAI321xp33_ASAP7_75t_L g565 ( 
.A1(n_559),
.A2(n_555),
.A3(n_511),
.B1(n_497),
.B2(n_493),
.C(n_503),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_560),
.B(n_561),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_557),
.B(n_542),
.C(n_536),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_562),
.A2(n_554),
.B(n_556),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_564),
.A2(n_565),
.B(n_503),
.C(n_497),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_567),
.C(n_480),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_563),
.B(n_478),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_497),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_493),
.Y(n_570)
);


endmodule