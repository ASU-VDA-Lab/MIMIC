module real_aes_3204_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_938;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_954;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_898;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_0), .A2(n_570), .B1(n_571), .B2(n_574), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_0), .Y(n_574) );
INVx1_ASAP7_75t_L g653 ( .A(n_1), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_2), .A2(n_16), .B1(n_174), .B2(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g617 ( .A(n_3), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_4), .A2(n_35), .B1(n_140), .B2(n_226), .Y(n_225) );
INVx1_ASAP7_75t_SL g671 ( .A(n_5), .Y(n_671) );
INVxp67_ASAP7_75t_L g550 ( .A(n_6), .Y(n_550) );
INVx1_ASAP7_75t_L g938 ( .A(n_6), .Y(n_938) );
INVx1_ASAP7_75t_L g942 ( .A(n_6), .Y(n_942) );
NAND3xp33_ASAP7_75t_SL g953 ( .A(n_6), .B(n_954), .C(n_955), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_7), .A2(n_90), .B1(n_214), .B2(n_215), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_8), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_9), .B(n_255), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_10), .A2(n_36), .B1(n_245), .B2(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g181 ( .A(n_11), .Y(n_181) );
OAI22xp33_ASAP7_75t_SL g111 ( .A1(n_12), .A2(n_112), .B1(n_113), .B2(n_114), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_13), .A2(n_63), .B1(n_572), .B2(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_13), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_14), .A2(n_58), .B1(n_251), .B2(n_658), .Y(n_657) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_15), .A2(n_70), .B(n_126), .Y(n_125) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_15), .A2(n_70), .B(n_126), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_17), .B(n_177), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_18), .A2(n_82), .B1(n_227), .B2(n_250), .Y(n_612) );
INVx2_ASAP7_75t_L g607 ( .A(n_19), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_20), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g178 ( .A(n_21), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_22), .B(n_316), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_23), .A2(n_27), .B1(n_214), .B2(n_215), .Y(n_588) );
BUFx3_ASAP7_75t_L g107 ( .A(n_24), .Y(n_107) );
BUFx8_ASAP7_75t_SL g564 ( .A(n_24), .Y(n_564) );
O2A1O1Ixp5_ASAP7_75t_L g603 ( .A1(n_25), .A2(n_140), .B(n_193), .C(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_26), .A2(n_66), .B1(n_141), .B2(n_615), .Y(n_614) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_28), .A2(n_187), .B(n_190), .C(n_192), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_29), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_30), .B(n_231), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_31), .A2(n_83), .B1(n_173), .B2(n_198), .Y(n_663) );
INVx1_ASAP7_75t_L g555 ( .A(n_32), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_32), .B(n_81), .Y(n_952) );
INVx1_ASAP7_75t_L g600 ( .A(n_33), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_34), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_34), .Y(n_567) );
AND2x2_ASAP7_75t_L g955 ( .A(n_37), .B(n_956), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_38), .B(n_310), .Y(n_649) );
INVx2_ASAP7_75t_L g605 ( .A(n_39), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_40), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_41), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_42), .A2(n_105), .B1(n_950), .B2(n_957), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_43), .A2(n_48), .B1(n_217), .B2(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_44), .A2(n_69), .B1(n_133), .B2(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_45), .B(n_227), .Y(n_308) );
INVx2_ASAP7_75t_L g123 ( .A(n_46), .Y(n_123) );
INVx2_ASAP7_75t_L g627 ( .A(n_47), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_49), .B(n_231), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_50), .B(n_203), .Y(n_221) );
INVx1_ASAP7_75t_SL g674 ( .A(n_51), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_52), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_53), .A2(n_146), .B(n_173), .C(n_175), .Y(n_172) );
INVx1_ASAP7_75t_L g275 ( .A(n_54), .Y(n_275) );
INVx1_ASAP7_75t_L g686 ( .A(n_55), .Y(n_686) );
INVx2_ASAP7_75t_L g201 ( .A(n_56), .Y(n_201) );
INVx1_ASAP7_75t_L g126 ( .A(n_57), .Y(n_126) );
AND2x4_ASAP7_75t_L g148 ( .A(n_59), .B(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g205 ( .A(n_59), .B(n_149), .Y(n_205) );
INVx2_ASAP7_75t_L g136 ( .A(n_60), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_61), .A2(n_110), .B1(n_544), .B2(n_545), .Y(n_109) );
INVx1_ASAP7_75t_L g545 ( .A(n_61), .Y(n_545) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_62), .Y(n_138) );
INVx1_ASAP7_75t_L g572 ( .A(n_63), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_64), .A2(n_98), .B1(n_115), .B2(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_64), .Y(n_116) );
INVx1_ASAP7_75t_SL g191 ( .A(n_65), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_67), .B(n_632), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_68), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_71), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_72), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_73), .A2(n_140), .B(n_144), .C(n_146), .Y(n_139) );
OR2x6_ASAP7_75t_L g552 ( .A(n_74), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g954 ( .A(n_74), .Y(n_954) );
INVx1_ASAP7_75t_L g271 ( .A(n_75), .Y(n_271) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_76), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_77), .B(n_169), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_78), .B(n_245), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g167 ( .A(n_79), .B(n_168), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_80), .A2(n_129), .B(n_132), .C(n_137), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_80), .A2(n_129), .B(n_132), .C(n_137), .Y(n_326) );
INVx1_ASAP7_75t_L g554 ( .A(n_81), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_84), .A2(n_95), .B1(n_249), .B2(n_251), .Y(n_248) );
INVx1_ASAP7_75t_L g956 ( .A(n_85), .Y(n_956) );
BUFx5_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_87), .B(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_88), .B(n_632), .Y(n_672) );
INVx2_ASAP7_75t_L g630 ( .A(n_89), .Y(n_630) );
INVx1_ASAP7_75t_L g636 ( .A(n_91), .Y(n_636) );
INVx2_ASAP7_75t_L g693 ( .A(n_92), .Y(n_693) );
INVx2_ASAP7_75t_SL g149 ( .A(n_93), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_94), .B(n_316), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_96), .B(n_125), .Y(n_272) );
INVx1_ASAP7_75t_SL g237 ( .A(n_97), .Y(n_237) );
INVx1_ASAP7_75t_L g115 ( .A(n_98), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_99), .B(n_150), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_100), .Y(n_558) );
AND2x2_ASAP7_75t_L g254 ( .A(n_101), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_SL g199 ( .A(n_102), .Y(n_199) );
AO32x2_ASAP7_75t_L g584 ( .A1(n_103), .A2(n_261), .A3(n_286), .B1(n_585), .B2(n_589), .Y(n_584) );
AO22x2_ASAP7_75t_L g698 ( .A1(n_103), .A2(n_285), .B1(n_585), .B2(n_699), .Y(n_698) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_108), .B(n_561), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI21x1_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_546), .B(n_556), .Y(n_108) );
INVx1_ASAP7_75t_L g544 ( .A(n_110), .Y(n_544) );
XNOR2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_117), .Y(n_110) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AO22x2_ASAP7_75t_L g575 ( .A1(n_117), .A2(n_576), .B1(n_936), .B2(n_939), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_117), .A2(n_576), .B1(n_937), .B2(n_944), .Y(n_943) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_417), .Y(n_117) );
NOR3xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_348), .C(n_387), .Y(n_118) );
OAI211xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_152), .B(n_238), .C(n_331), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_120), .A2(n_423), .B1(n_424), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_121), .B(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g293 ( .A(n_121), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_121), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g410 ( .A(n_121), .Y(n_410) );
AND2x2_ASAP7_75t_L g452 ( .A(n_121), .B(n_241), .Y(n_452) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_122), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g259 ( .A(n_124), .Y(n_259) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
BUFx3_ASAP7_75t_L g255 ( .A(n_125), .Y(n_255) );
INVx1_ASAP7_75t_L g590 ( .A(n_125), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_125), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_125), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_125), .B(n_634), .Y(n_654) );
NOR2xp67_ASAP7_75t_L g660 ( .A(n_125), .B(n_634), .Y(n_660) );
INVx1_ASAP7_75t_L g700 ( .A(n_125), .Y(n_700) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_139), .C(n_147), .D(n_150), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g650 ( .A(n_130), .Y(n_650) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp33_ASAP7_75t_L g165 ( .A(n_131), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g214 ( .A(n_131), .Y(n_214) );
INVx2_ASAP7_75t_L g231 ( .A(n_131), .Y(n_231) );
INVx2_ASAP7_75t_L g245 ( .A(n_131), .Y(n_245) );
INVx2_ASAP7_75t_L g251 ( .A(n_131), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_136), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_133), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g282 ( .A(n_134), .Y(n_282) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
INVx2_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
INVx6_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx1_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx2_ASAP7_75t_SL g219 ( .A(n_137), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_137), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_137), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g613 ( .A(n_137), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_137), .A2(n_217), .B(n_630), .C(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_137), .B(n_660), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g669 ( .A1(n_137), .A2(n_670), .B(n_671), .C(n_672), .Y(n_669) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
INVxp67_ASAP7_75t_L g196 ( .A(n_138), .Y(n_196) );
INVx4_ASAP7_75t_L g283 ( .A(n_138), .Y(n_283) );
INVx1_ASAP7_75t_L g665 ( .A(n_138), .Y(n_665) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_139), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_140), .B(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g632 ( .A(n_142), .Y(n_632) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g218 ( .A(n_143), .Y(n_218) );
INVx3_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_146), .A2(n_626), .B(n_627), .C(n_628), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_146), .A2(n_245), .B(n_674), .C(n_675), .Y(n_673) );
NOR2x1_ASAP7_75t_SL g157 ( .A(n_147), .B(n_158), .Y(n_157) );
AOI221x1_ASAP7_75t_L g594 ( .A1(n_147), .A2(n_595), .B1(n_597), .B2(n_599), .C(n_601), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_147), .B(n_232), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_147), .B(n_232), .C(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_147), .B(n_192), .Y(n_688) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_151), .B(n_237), .Y(n_236) );
NAND2x1_ASAP7_75t_L g152 ( .A(n_153), .B(n_182), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g353 ( .A(n_155), .Y(n_353) );
AND2x2_ASAP7_75t_L g386 ( .A(n_155), .B(n_345), .Y(n_386) );
AND2x2_ASAP7_75t_L g414 ( .A(n_155), .B(n_303), .Y(n_414) );
AND2x2_ASAP7_75t_L g446 ( .A(n_155), .B(n_432), .Y(n_446) );
INVx1_ASAP7_75t_L g534 ( .A(n_155), .Y(n_534) );
OR2x2_ASAP7_75t_L g539 ( .A(n_155), .B(n_532), .Y(n_539) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OR2x2_ASAP7_75t_L g330 ( .A(n_156), .B(n_266), .Y(n_330) );
OR2x2_ASAP7_75t_L g341 ( .A(n_156), .B(n_301), .Y(n_341) );
AND2x4_ASAP7_75t_L g361 ( .A(n_156), .B(n_301), .Y(n_361) );
INVx1_ASAP7_75t_L g369 ( .A(n_156), .Y(n_369) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_156), .Y(n_456) );
AND2x2_ASAP7_75t_L g471 ( .A(n_156), .B(n_266), .Y(n_471) );
AO31x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_163), .A3(n_171), .B(n_179), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g610 ( .A(n_159), .B(n_205), .Y(n_610) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_160), .B(n_634), .Y(n_668) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
BUFx3_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_170), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
INVx2_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
INVx1_ASAP7_75t_L g646 ( .A(n_169), .Y(n_646) );
INVx1_ASAP7_75t_L g658 ( .A(n_169), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_170), .A2(n_312), .B(n_314), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_170), .A2(n_193), .B1(n_586), .B2(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVxp67_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
INVx2_ASAP7_75t_L g246 ( .A(n_174), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_178), .Y(n_175) );
INVx1_ASAP7_75t_L g596 ( .A(n_176), .Y(n_596) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g189 ( .A(n_177), .Y(n_189) );
INVx1_ASAP7_75t_L g277 ( .A(n_177), .Y(n_277) );
INVx1_ASAP7_75t_L g313 ( .A(n_177), .Y(n_313) );
INVx2_ASAP7_75t_SL g587 ( .A(n_177), .Y(n_587) );
INVx1_ASAP7_75t_L g615 ( .A(n_177), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
BUFx3_ASAP7_75t_L g286 ( .A(n_180), .Y(n_286) );
INVx3_ASAP7_75t_L g316 ( .A(n_180), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_180), .B(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_180), .B(n_617), .Y(n_616) );
AOI322xp5_ASAP7_75t_L g401 ( .A1(n_182), .A2(n_389), .A3(n_402), .B1(n_403), .B2(n_405), .C1(n_407), .C2(n_412), .Y(n_401) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_207), .Y(n_182) );
INVx1_ASAP7_75t_L g287 ( .A(n_183), .Y(n_287) );
BUFx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g339 ( .A(n_184), .B(n_304), .Y(n_339) );
INVx2_ASAP7_75t_SL g346 ( .A(n_184), .Y(n_346) );
AND2x2_ASAP7_75t_L g416 ( .A(n_184), .B(n_301), .Y(n_416) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g298 ( .A(n_185), .Y(n_298) );
INVx3_ASAP7_75t_L g433 ( .A(n_185), .Y(n_433) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_194), .B(n_206), .Y(n_185) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_189), .B(n_652), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_189), .A2(n_214), .B1(n_690), .B2(n_691), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_192), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_192), .B(n_248), .Y(n_247) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_193), .A2(n_645), .B(n_647), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_197), .B(n_202), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_195), .A2(n_213), .B1(n_216), .B2(n_219), .Y(n_212) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx3_ASAP7_75t_L g253 ( .A(n_203), .Y(n_253) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g235 ( .A(n_205), .Y(n_235) );
AND2x2_ASAP7_75t_L g252 ( .A(n_205), .B(n_253), .Y(n_252) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_205), .Y(n_261) );
INVx3_ASAP7_75t_L g634 ( .A(n_205), .Y(n_634) );
AND2x2_ASAP7_75t_L g699 ( .A(n_205), .B(n_700), .Y(n_699) );
AND2x6_ASAP7_75t_SL g347 ( .A(n_207), .B(n_240), .Y(n_347) );
AND2x2_ASAP7_75t_L g478 ( .A(n_207), .B(n_441), .Y(n_478) );
AND2x2_ASAP7_75t_L g489 ( .A(n_207), .B(n_459), .Y(n_489) );
AND2x4_ASAP7_75t_L g536 ( .A(n_207), .B(n_293), .Y(n_536) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
OR2x2_ASAP7_75t_L g290 ( .A(n_208), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g320 ( .A(n_208), .Y(n_320) );
AOI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B(n_220), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_209), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_212), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g670 ( .A(n_215), .Y(n_670) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_217), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g250 ( .A(n_218), .Y(n_250) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_221), .A2(n_259), .B(n_260), .Y(n_258) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_222), .B(n_322), .Y(n_321) );
NAND2x1_ASAP7_75t_L g364 ( .A(n_222), .B(n_295), .Y(n_364) );
INVx1_ASAP7_75t_L g485 ( .A(n_222), .Y(n_485) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g292 ( .A(n_223), .Y(n_292) );
AOI21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_228), .B(n_236), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_232), .B(n_233), .Y(n_228) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_232), .B(n_244), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_232), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_611) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_234), .A2(n_307), .B(n_311), .Y(n_306) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_235), .A2(n_272), .B(n_285), .Y(n_284) );
AOI222xp33_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_262), .B1(n_288), .B2(n_296), .C1(n_317), .C2(n_329), .Y(n_238) );
AND2x2_ASAP7_75t_L g484 ( .A(n_239), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_256), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_240), .B(n_321), .Y(n_377) );
INVx1_ASAP7_75t_L g520 ( .A(n_240), .Y(n_520) );
BUFx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_SL g295 ( .A(n_242), .Y(n_295) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_247), .A3(n_252), .B(n_254), .Y(n_242) );
INVx1_ASAP7_75t_L g601 ( .A(n_246), .Y(n_601) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g269 ( .A(n_251), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_253), .B(n_261), .Y(n_323) );
AO21x2_ASAP7_75t_L g709 ( .A1(n_253), .A2(n_679), .B(n_692), .Y(n_709) );
INVx1_ASAP7_75t_L g365 ( .A(n_256), .Y(n_365) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_258), .Y(n_385) );
AND2x2_ASAP7_75t_L g436 ( .A(n_258), .B(n_291), .Y(n_436) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_259), .A2(n_306), .B(n_315), .Y(n_355) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_287), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g438 ( .A(n_265), .B(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_278), .B(n_284), .Y(n_266) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_267), .A2(n_278), .B(n_284), .Y(n_302) );
NAND3x1_ASAP7_75t_L g267 ( .A(n_268), .B(n_272), .C(n_273), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g280 ( .A(n_276), .Y(n_280) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_280), .B(n_281), .C(n_283), .Y(n_278) );
INVx1_ASAP7_75t_L g684 ( .A(n_282), .Y(n_684) );
INVx2_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_283), .B(n_653), .Y(n_652) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_285), .A2(n_306), .B(n_315), .Y(n_305) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_286), .A2(n_594), .A3(n_602), .B(n_606), .Y(n_593) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_293), .Y(n_288) );
AND2x4_ASAP7_75t_L g458 ( .A(n_289), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_290), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_513) );
AND2x4_ASAP7_75t_L g374 ( .A(n_291), .B(n_322), .Y(n_374) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g335 ( .A(n_292), .Y(n_335) );
AND2x2_ASAP7_75t_L g403 ( .A(n_293), .B(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_293), .Y(n_425) );
INVx2_ASAP7_75t_SL g437 ( .A(n_293), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_293), .B(n_464), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_294), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g359 ( .A(n_294), .Y(n_359) );
BUFx2_ASAP7_75t_SL g441 ( .A(n_294), .Y(n_441) );
AND2x2_ASAP7_75t_L g459 ( .A(n_294), .B(n_322), .Y(n_459) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_297), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g476 ( .A(n_297), .B(n_354), .Y(n_476) );
AND2x2_ASAP7_75t_L g498 ( .A(n_297), .B(n_361), .Y(n_498) );
INVx2_ASAP7_75t_R g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g427 ( .A(n_298), .Y(n_427) );
INVx1_ASAP7_75t_L g483 ( .A(n_299), .Y(n_483) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g501 ( .A(n_300), .B(n_368), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g345 ( .A(n_302), .B(n_304), .Y(n_345) );
AND2x2_ASAP7_75t_L g354 ( .A(n_302), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_SL g370 ( .A(n_303), .Y(n_370) );
INVx1_ASAP7_75t_L g394 ( .A(n_303), .Y(n_394) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_303), .Y(n_448) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g431 ( .A(n_304), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B(n_310), .Y(n_307) );
AND2x2_ASAP7_75t_L g597 ( .A(n_310), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g599 ( .A(n_310), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g372 ( .A(n_319), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_335), .Y(n_356) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_328), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_329), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g473 ( .A(n_330), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g496 ( .A(n_330), .B(n_346), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_336), .B1(n_342), .B2(n_347), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
INVx1_ASAP7_75t_L g464 ( .A(n_335), .Y(n_464) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_338), .B(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2x1_ASAP7_75t_SL g455 ( .A(n_339), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g474 ( .A(n_339), .Y(n_474) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_343), .A2(n_454), .B(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x2_ASAP7_75t_L g512 ( .A(n_345), .B(n_470), .Y(n_512) );
INVx2_ASAP7_75t_L g532 ( .A(n_345), .Y(n_532) );
AND2x2_ASAP7_75t_L g391 ( .A(n_346), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g406 ( .A(n_346), .Y(n_406) );
INVx2_ASAP7_75t_L g470 ( .A(n_346), .Y(n_470) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_346), .Y(n_541) );
OAI311xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_356), .A3(n_357), .B1(n_360), .C1(n_375), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x4_ASAP7_75t_L g389 ( .A(n_354), .B(n_369), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_354), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g445 ( .A(n_354), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g506 ( .A(n_354), .Y(n_506) );
AND2x2_ASAP7_75t_L g493 ( .A(n_355), .B(n_433), .Y(n_493) );
AND2x2_ASAP7_75t_L g511 ( .A(n_356), .B(n_359), .Y(n_511) );
INVx1_ASAP7_75t_L g521 ( .A(n_356), .Y(n_521) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_358), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_366), .B2(n_371), .Y(n_360) );
INVx2_ASAP7_75t_L g380 ( .A(n_361), .Y(n_380) );
AND2x2_ASAP7_75t_L g392 ( .A(n_361), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_361), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g528 ( .A(n_361), .B(n_431), .Y(n_528) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NOR2x1p5_ASAP7_75t_L g384 ( .A(n_364), .B(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2x2_ASAP7_75t_L g405 ( .A(n_367), .B(n_406), .Y(n_405) );
OR2x6_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g491 ( .A(n_369), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_372), .B(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g504 ( .A(n_373), .B(n_441), .Y(n_504) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g444 ( .A(n_374), .B(n_441), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_374), .B(n_385), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_381), .B2(n_386), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g400 ( .A(n_377), .Y(n_400) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
AND2x2_ASAP7_75t_L g543 ( .A(n_384), .B(n_409), .Y(n_543) );
INVx2_ASAP7_75t_L g399 ( .A(n_385), .Y(n_399) );
INVx2_ASAP7_75t_L g451 ( .A(n_385), .Y(n_451) );
INVx1_ASAP7_75t_L g510 ( .A(n_385), .Y(n_510) );
INVx1_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_395), .C(n_401), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_392), .A2(n_461), .B1(n_465), .B2(n_469), .C(n_472), .Y(n_460) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_397), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_397), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g487 ( .A(n_403), .Y(n_487) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g463 ( .A(n_410), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g529 ( .A1(n_413), .A2(n_530), .B(n_535), .Y(n_529) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g447 ( .A(n_416), .B(n_448), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_479), .C(n_507), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_460), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_428), .C(n_453), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_434), .B1(n_438), .B2(n_440), .C(n_443), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g439 ( .A(n_431), .Y(n_439) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_433), .B(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g442 ( .A(n_436), .Y(n_442) );
INVx1_ASAP7_75t_L g542 ( .A(n_438), .Y(n_542) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_447), .B2(n_449), .Y(n_443) );
INVx2_ASAP7_75t_L g517 ( .A(n_446), .Y(n_517) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g509 ( .A(n_452), .B(n_510), .Y(n_509) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g499 ( .A(n_468), .Y(n_499) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .B(n_477), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_494), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B1(n_486), .B2(n_490), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_484), .A2(n_538), .B1(n_542), .B2(n_543), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g516 ( .A(n_493), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_499), .B1(n_500), .B2(n_502), .C(n_505), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g527 ( .A(n_504), .Y(n_527) );
NAND3xp33_ASAP7_75t_SL g507 ( .A(n_508), .B(n_522), .C(n_537), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_511), .B(n_512), .C(n_513), .Y(n_508) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_525), .B(n_528), .C(n_529), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_SL g676 ( .A(n_545), .B(n_637), .Y(n_676) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx10_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx12f_ASAP7_75t_L g560 ( .A(n_548), .Y(n_560) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
OR2x6_ASAP7_75t_L g937 ( .A(n_551), .B(n_938), .Y(n_937) );
INVx8_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g941 ( .A(n_552), .B(n_942), .Y(n_941) );
OR2x6_ASAP7_75t_L g949 ( .A(n_552), .B(n_942), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_557), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_575), .B1(n_943), .B2(n_945), .C(n_946), .Y(n_565) );
INVx1_ASAP7_75t_L g945 ( .A(n_566), .Y(n_945) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_841), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_579), .B(n_737), .C(n_784), .D(n_816), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_721), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_694), .Y(n_580) );
OAI21xp33_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_618), .B(n_639), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_591), .Y(n_582) );
INVx1_ASAP7_75t_L g736 ( .A(n_583), .Y(n_736) );
AND2x2_ASAP7_75t_SL g741 ( .A(n_583), .B(n_622), .Y(n_741) );
AND2x2_ASAP7_75t_L g820 ( .A(n_583), .B(n_714), .Y(n_820) );
OR2x2_ASAP7_75t_L g844 ( .A(n_583), .B(n_845), .Y(n_844) );
AND2x2_ASAP7_75t_L g862 ( .A(n_583), .B(n_744), .Y(n_862) );
AND2x2_ASAP7_75t_L g884 ( .A(n_583), .B(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g900 ( .A(n_583), .Y(n_900) );
BUFx8_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g768 ( .A(n_584), .Y(n_768) );
AND2x2_ASAP7_75t_L g916 ( .A(n_584), .B(n_767), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_587), .B(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g678 ( .A(n_589), .Y(n_678) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_590), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g824 ( .A(n_591), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g905 ( .A(n_591), .B(n_761), .Y(n_905) );
INVxp67_ASAP7_75t_SL g921 ( .A(n_591), .Y(n_921) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_608), .Y(n_591) );
INVx1_ASAP7_75t_L g781 ( .A(n_592), .Y(n_781) );
INVx2_ASAP7_75t_SL g878 ( .A(n_592), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_592), .B(n_768), .Y(n_891) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g638 ( .A(n_593), .Y(n_638) );
OR2x2_ASAP7_75t_L g703 ( .A(n_593), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g714 ( .A(n_593), .B(n_623), .Y(n_714) );
AND2x2_ASAP7_75t_L g744 ( .A(n_593), .B(n_701), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_593), .B(n_704), .Y(n_797) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_608), .Y(n_727) );
INVx2_ASAP7_75t_L g760 ( .A(n_608), .Y(n_760) );
AND2x2_ASAP7_75t_L g927 ( .A(n_608), .B(n_701), .Y(n_927) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g621 ( .A(n_609), .Y(n_621) );
INVx1_ASAP7_75t_L g704 ( .A(n_609), .Y(n_704) );
AOI21x1_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_616), .Y(n_609) );
INVx1_ASAP7_75t_L g626 ( .A(n_615), .Y(n_626) );
INVx2_ASAP7_75t_L g849 ( .A(n_618), .Y(n_849) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g713 ( .A(n_619), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_619), .B(n_697), .Y(n_799) );
INVx4_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_SL g739 ( .A(n_620), .Y(n_739) );
AND2x2_ASAP7_75t_L g858 ( .A(n_620), .B(n_744), .Y(n_858) );
AND2x2_ASAP7_75t_L g871 ( .A(n_620), .B(n_622), .Y(n_871) );
INVx2_ASAP7_75t_L g874 ( .A(n_620), .Y(n_874) );
BUFx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g767 ( .A(n_621), .Y(n_767) );
INVx2_ASAP7_75t_L g845 ( .A(n_622), .Y(n_845) );
AND2x4_ASAP7_75t_L g622 ( .A(n_623), .B(n_638), .Y(n_622) );
INVx2_ASAP7_75t_L g701 ( .A(n_623), .Y(n_701) );
INVx1_ASAP7_75t_L g762 ( .A(n_623), .Y(n_762) );
BUFx3_ASAP7_75t_L g780 ( .A(n_623), .Y(n_780) );
AND2x4_ASAP7_75t_L g825 ( .A(n_623), .B(n_768), .Y(n_825) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AO31x2_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_629), .A3(n_633), .B(n_635), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_666), .Y(n_639) );
AND2x2_ASAP7_75t_L g887 ( .A(n_640), .B(n_719), .Y(n_887) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_655), .Y(n_640) );
INVx2_ASAP7_75t_L g711 ( .A(n_641), .Y(n_711) );
INVx1_ASAP7_75t_L g734 ( .A(n_641), .Y(n_734) );
AND2x2_ASAP7_75t_L g750 ( .A(n_641), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g813 ( .A(n_641), .Y(n_813) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_641), .Y(n_924) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B(n_654), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g710 ( .A(n_655), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g730 ( .A(n_655), .Y(n_730) );
INVx2_ASAP7_75t_L g748 ( .A(n_655), .Y(n_748) );
INVx1_ASAP7_75t_L g772 ( .A(n_655), .Y(n_772) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_656), .B(n_662), .Y(n_655) );
AND2x2_ASAP7_75t_SL g718 ( .A(n_656), .B(n_662), .Y(n_718) );
OA21x2_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B(n_661), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_660), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g798 ( .A(n_666), .Y(n_798) );
AND2x2_ASAP7_75t_L g847 ( .A(n_666), .B(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g935 ( .A(n_666), .B(n_710), .Y(n_935) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_677), .Y(n_666) );
OR2x2_ASAP7_75t_L g708 ( .A(n_667), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g720 ( .A(n_667), .Y(n_720) );
INVx2_ASAP7_75t_L g751 ( .A(n_667), .Y(n_751) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_667), .Y(n_777) );
INVx1_ASAP7_75t_L g811 ( .A(n_667), .Y(n_811) );
INVx1_ASAP7_75t_L g857 ( .A(n_667), .Y(n_857) );
AO31x2_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .A3(n_673), .B(n_676), .Y(n_667) );
OR2x2_ASAP7_75t_L g756 ( .A(n_677), .B(n_711), .Y(n_756) );
AND2x2_ASAP7_75t_L g812 ( .A(n_677), .B(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g880 ( .A(n_677), .B(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g903 ( .A(n_677), .B(n_748), .Y(n_903) );
AO21x2_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_692), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_687), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_705), .B1(n_712), .B2(n_715), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_702), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_696), .A2(n_833), .B1(n_898), .B2(n_901), .C(n_904), .Y(n_897) );
INVx4_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g839 ( .A(n_697), .B(n_840), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_697), .B(n_921), .Y(n_920) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g724 ( .A(n_698), .Y(n_724) );
INVx1_ASAP7_75t_L g763 ( .A(n_698), .Y(n_763) );
AND2x4_ASAP7_75t_L g791 ( .A(n_698), .B(n_780), .Y(n_791) );
AND2x2_ASAP7_75t_L g815 ( .A(n_702), .B(n_779), .Y(n_815) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g840 ( .A(n_703), .Y(n_840) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_704), .Y(n_792) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp67_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g806 ( .A(n_708), .B(n_771), .Y(n_806) );
AND2x2_ASAP7_75t_L g719 ( .A(n_709), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g749 ( .A(n_709), .Y(n_749) );
BUFx2_ASAP7_75t_L g783 ( .A(n_709), .Y(n_783) );
AND2x2_ASAP7_75t_L g827 ( .A(n_710), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_710), .B(n_783), .Y(n_837) );
AND2x2_ASAP7_75t_L g888 ( .A(n_710), .B(n_782), .Y(n_888) );
AND2x2_ASAP7_75t_L g911 ( .A(n_710), .B(n_801), .Y(n_911) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g723 ( .A(n_714), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g765 ( .A(n_714), .Y(n_765) );
INVx2_ASAP7_75t_L g831 ( .A(n_714), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_715), .A2(n_905), .B1(n_906), .B2(n_907), .Y(n_904) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2x1p5_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_717), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g856 ( .A(n_718), .B(n_734), .Y(n_856) );
INVx2_ASAP7_75t_L g881 ( .A(n_718), .Y(n_881) );
AND2x2_ASAP7_75t_L g914 ( .A(n_718), .B(n_734), .Y(n_914) );
AND2x4_ASAP7_75t_L g726 ( .A(n_719), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g853 ( .A(n_719), .Y(n_853) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_720), .Y(n_755) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_720), .Y(n_860) );
OAI32xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .A3(n_728), .B1(n_731), .B2(n_735), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_722), .A2(n_931), .B1(n_932), .B2(n_934), .Y(n_930) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_726), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g830 ( .A(n_727), .Y(n_830) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI311xp33_ASAP7_75t_L g816 ( .A1(n_729), .A2(n_817), .A3(n_818), .B(n_821), .C(n_832), .Y(n_816) );
BUFx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g809 ( .A(n_730), .B(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND5xp2_ASAP7_75t_L g775 ( .A(n_733), .B(n_776), .C(n_778), .D(n_781), .E(n_782), .Y(n_775) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_752), .C(n_774), .Y(n_737) );
AOI31xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .A3(n_742), .B(n_745), .Y(n_738) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g899 ( .A(n_744), .B(n_900), .Y(n_899) );
AND2x2_ASAP7_75t_L g915 ( .A(n_744), .B(n_916), .Y(n_915) );
AND2x2_ASAP7_75t_L g933 ( .A(n_744), .B(n_760), .Y(n_933) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_750), .Y(n_746) );
AND2x4_ASAP7_75t_L g922 ( .A(n_747), .B(n_923), .Y(n_922) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_748), .Y(n_835) );
BUFx2_ASAP7_75t_L g848 ( .A(n_748), .Y(n_848) );
AND2x4_ASAP7_75t_L g801 ( .A(n_749), .B(n_802), .Y(n_801) );
OR2x2_ASAP7_75t_L g861 ( .A(n_749), .B(n_813), .Y(n_861) );
AND2x2_ASAP7_75t_L g902 ( .A(n_750), .B(n_903), .Y(n_902) );
AND2x2_ASAP7_75t_L g908 ( .A(n_750), .B(n_772), .Y(n_908) );
INVx1_ASAP7_75t_L g802 ( .A(n_751), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_757), .B1(n_764), .B2(n_769), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g788 ( .A(n_754), .Y(n_788) );
OAI322xp33_ASAP7_75t_L g793 ( .A1(n_754), .A2(n_794), .A3(n_795), .B1(n_798), .B2(n_799), .C1(n_800), .C2(n_803), .Y(n_793) );
OR2x6_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVxp67_ASAP7_75t_L g773 ( .A(n_756), .Y(n_773) );
INVxp67_ASAP7_75t_SL g836 ( .A(n_756), .Y(n_836) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
BUFx3_ASAP7_75t_L g819 ( .A(n_760), .Y(n_819) );
AND2x2_ASAP7_75t_L g906 ( .A(n_760), .B(n_779), .Y(n_906) );
INVx1_ASAP7_75t_L g794 ( .A(n_761), .Y(n_794) );
AND2x4_ASAP7_75t_SL g761 ( .A(n_762), .B(n_763), .Y(n_761) );
OR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g804 ( .A(n_766), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AND2x2_ASAP7_75t_L g877 ( .A(n_768), .B(n_878), .Y(n_877) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
AND2x2_ASAP7_75t_L g776 ( .A(n_771), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g787 ( .A(n_771), .Y(n_787) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVxp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_779), .B(n_874), .Y(n_873) );
INVx2_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI211xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_789), .B(n_793), .C(n_805), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
OR2x2_ASAP7_75t_L g918 ( .A(n_792), .B(n_891), .Y(n_918) );
OAI211xp5_ASAP7_75t_L g909 ( .A1(n_794), .A2(n_910), .B(n_912), .C(n_919), .Y(n_909) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g885 ( .A(n_797), .Y(n_885) );
INVx1_ASAP7_75t_L g817 ( .A(n_801), .Y(n_817) );
AND2x2_ASAP7_75t_L g867 ( .A(n_801), .B(n_848), .Y(n_867) );
AND2x4_ASAP7_75t_L g894 ( .A(n_801), .B(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g913 ( .A(n_801), .B(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B(n_814), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AND2x4_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .Y(n_808) );
INVxp67_ASAP7_75t_L g828 ( .A(n_810), .Y(n_828) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_810), .Y(n_870) );
AND2x2_ASAP7_75t_L g929 ( .A(n_810), .B(n_924), .Y(n_929) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g822 ( .A(n_812), .Y(n_822) );
AND2x2_ASAP7_75t_L g865 ( .A(n_813), .B(n_857), .Y(n_865) );
INVx1_ASAP7_75t_L g895 ( .A(n_813), .Y(n_895) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .B1(n_826), .B2(n_829), .Y(n_821) );
INVx2_ASAP7_75t_SL g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OR2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_837), .B(n_838), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g893 ( .A(n_835), .Y(n_893) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_896), .Y(n_841) );
NOR3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_863), .C(n_882), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_846), .B1(n_849), .B2(n_850), .C(n_854), .Y(n_843) );
OAI211xp5_ASAP7_75t_L g863 ( .A1(n_844), .A2(n_864), .B(n_866), .C(n_872), .Y(n_863) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g852 ( .A(n_848), .Y(n_852) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
NOR2x1p5_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_858), .B1(n_859), .B2(n_862), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_856), .B(n_870), .Y(n_869) );
NOR2xp67_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AND2x4_ASAP7_75t_L g879 ( .A(n_865), .B(n_880), .Y(n_879) );
OAI21xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B(n_871), .Y(n_866) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_875), .B(n_879), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_876), .B(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI22xp33_ASAP7_75t_SL g882 ( .A1(n_883), .A2(n_886), .B1(n_889), .B2(n_892), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_888), .A2(n_913), .B1(n_915), .B2(n_917), .Y(n_912) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_909), .C(n_930), .Y(n_896) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
AND2x4_ASAP7_75t_L g928 ( .A(n_903), .B(n_929), .Y(n_928) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g931 ( .A(n_913), .Y(n_931) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_922), .B1(n_925), .B2(n_928), .Y(n_919) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_937), .Y(n_936) );
BUFx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_SL g944 ( .A(n_941), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
BUFx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
BUFx4_ASAP7_75t_SL g959 ( .A(n_951), .Y(n_959) );
OR2x2_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .Y(n_951) );
BUFx3_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
endmodule