module real_jpeg_23589_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_67),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_47),
.B(n_54),
.C(n_121),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_2),
.A2(n_39),
.B1(n_42),
.B2(n_47),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_26),
.C(n_90),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_71),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_82),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_87)
);

INVx8_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_39),
.B1(n_47),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_84),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_39),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_11),
.A2(n_39),
.B1(n_47),
.B2(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_61),
.B1(n_99),
.B2(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_61),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_24),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_14),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_14),
.A2(n_24),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_128),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_107),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_18),
.B(n_107),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_77),
.B2(n_78),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_48),
.B1(n_75),
.B2(n_76),
.Y(n_20)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_35),
.B2(n_36),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_25),
.A2(n_26),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_25),
.B(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_29),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_31),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B(n_41),
.C(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_37),
.A2(n_38),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_46),
.C(n_47),
.Y(n_45)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_41),
.A2(n_42),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_42),
.A2(n_51),
.B(n_55),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_42),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_42),
.B(n_88),
.Y(n_171)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_65),
.C(n_68),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_52),
.B1(n_89),
.B2(n_90),
.Y(n_94)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_52),
.B(n_150),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_62),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_60),
.B(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_63),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_71),
.A2(n_158),
.B(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_96),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_92),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_88),
.A2(n_92),
.B(n_138),
.Y(n_180)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_115),
.B1(n_117),
.B2(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_102),
.B(n_105),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_118),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_109),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_118),
.B1(n_119),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B(n_116),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_116),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_122),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_156),
.B(n_168),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_143),
.B(n_190),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_130),
.B(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.C(n_139),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_184),
.B(n_189),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_174),
.B(n_183),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_159),
.B(n_173),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_169),
.B(n_172),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_182),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_180),
.C(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_188),
.Y(n_189)
);


endmodule