module real_aes_11469_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_891, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_891;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_148;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_152;
wire n_836;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
wire n_869;
NAND2xp5_ASAP7_75t_L g182 ( .A(n_0), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g516 ( .A(n_1), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_2), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_3), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_4), .B(n_497), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_5), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_6), .B(n_189), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_7), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_8), .B(n_178), .Y(n_177) );
NOR2xp67_ASAP7_75t_L g844 ( .A(n_9), .B(n_92), .Y(n_844) );
INVx1_ASAP7_75t_L g882 ( .A(n_9), .Y(n_882) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_10), .B(n_162), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_11), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_12), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_13), .Y(n_858) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_14), .B(n_178), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_15), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_16), .B(n_165), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_17), .B(n_207), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_18), .B(n_178), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_19), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_20), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_21), .B(n_162), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_22), .B(n_189), .Y(n_222) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_23), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_24), .B(n_144), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_25), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_26), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_27), .B(n_144), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_28), .B(n_207), .Y(n_571) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_29), .Y(n_136) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_30), .A2(n_181), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_31), .B(n_162), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_32), .B(n_160), .Y(n_159) );
NAND2xp33_ASAP7_75t_SL g142 ( .A(n_33), .B(n_138), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_34), .B(n_162), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_35), .B(n_226), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_36), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_37), .B(n_135), .Y(n_269) );
INVx1_ASAP7_75t_L g843 ( .A(n_38), .Y(n_843) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_39), .A2(n_72), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_40), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_41), .B(n_162), .Y(n_505) );
AOI22xp5_ASAP7_75t_SL g850 ( .A1(n_42), .A2(n_101), .B1(n_851), .B2(n_852), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_42), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_43), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_44), .B(n_226), .Y(n_225) );
AND2x6_ASAP7_75t_L g149 ( .A(n_45), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_46), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_47), .B(n_126), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_48), .A2(n_86), .B1(n_497), .B2(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_49), .B(n_126), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_50), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_51), .B(n_156), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_52), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_53), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_54), .Y(n_534) );
INVx1_ASAP7_75t_L g150 ( .A(n_55), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_56), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_57), .B(n_212), .Y(n_211) );
OAI22xp5_ASAP7_75t_SL g835 ( .A1(n_58), .A2(n_91), .B1(n_836), .B2(n_837), .Y(n_835) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_58), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_59), .A2(n_114), .B1(n_115), .B2(n_477), .Y(n_113) );
INVxp33_ASAP7_75t_SL g477 ( .A(n_59), .Y(n_477) );
XOR2x1_ASAP7_75t_L g480 ( .A(n_59), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_60), .B(n_498), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_61), .B(n_498), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g137 ( .A(n_62), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_63), .B(n_226), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_64), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_65), .B(n_156), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_66), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g885 ( .A(n_67), .B(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g526 ( .A(n_68), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_69), .B(n_144), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_70), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_71), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_73), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_74), .B(n_178), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_75), .B(n_207), .Y(n_220) );
INVx1_ASAP7_75t_L g520 ( .A(n_76), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_77), .B(n_226), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_78), .Y(n_591) );
BUFx10_ASAP7_75t_L g841 ( .A(n_79), .Y(n_841) );
INVx1_ASAP7_75t_L g585 ( .A(n_80), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_81), .B(n_178), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_82), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_82), .B(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_83), .B(n_162), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_84), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_85), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_87), .B(n_156), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_88), .B(n_178), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_89), .A2(n_104), .B1(n_877), .B2(n_888), .Y(n_103) );
INVx1_ASAP7_75t_L g529 ( .A(n_90), .Y(n_529) );
INVx1_ASAP7_75t_L g836 ( .A(n_91), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_92), .B(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
BUFx2_ASAP7_75t_L g111 ( .A(n_94), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_94), .B(n_842), .Y(n_861) );
OR2x2_ASAP7_75t_L g866 ( .A(n_94), .B(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g887 ( .A(n_94), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_95), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_96), .B(n_160), .Y(n_267) );
INVx1_ASAP7_75t_L g886 ( .A(n_97), .Y(n_886) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_98), .B(n_189), .Y(n_197) );
NOR2xp67_ASAP7_75t_L g491 ( .A(n_99), .B(n_492), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_100), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_101), .Y(n_851) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_102), .B(n_156), .Y(n_595) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_838), .B(n_845), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_107), .B1(n_834), .B2(n_835), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_112), .B(n_478), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g479 ( .A(n_110), .Y(n_479) );
BUFx8_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_115), .Y(n_849) );
INVx1_ASAP7_75t_L g854 ( .A(n_115), .Y(n_854) );
NAND2x1p5_ASAP7_75t_L g115 ( .A(n_116), .B(n_398), .Y(n_115) );
NOR2x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_322), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_292), .Y(n_117) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_200), .B1(n_228), .B2(n_259), .C(n_272), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_152), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g351 ( .A(n_122), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_122), .B(n_350), .Y(n_416) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g300 ( .A(n_123), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g373 ( .A(n_123), .B(n_239), .Y(n_373) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g275 ( .A(n_124), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_124), .B(n_239), .Y(n_337) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_124), .Y(n_378) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g260 ( .A(n_125), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_125), .Y(n_345) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_131), .B(n_151), .Y(n_125) );
OAI21x1_ASAP7_75t_L g216 ( .A1(n_126), .A2(n_217), .B(n_225), .Y(n_216) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g199 ( .A(n_127), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_127), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx5_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g184 ( .A(n_129), .Y(n_184) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_141), .B(n_147), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_137), .C(n_139), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_134), .A2(n_535), .B1(n_541), .B2(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_135), .A2(n_162), .B1(n_174), .B2(n_175), .Y(n_173) );
INVx2_ASAP7_75t_L g497 ( .A(n_135), .Y(n_497) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_136), .Y(n_145) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx1_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
INVx2_ASAP7_75t_L g196 ( .A(n_138), .Y(n_196) );
INVx2_ASAP7_75t_L g493 ( .A(n_138), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_138), .Y(n_495) );
INVx2_ASAP7_75t_L g498 ( .A(n_138), .Y(n_498) );
INVx2_ASAP7_75t_SL g146 ( .A(n_139), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_139), .A2(n_159), .B(n_161), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_139), .A2(n_206), .B(n_208), .Y(n_205) );
INVx2_ASAP7_75t_SL g224 ( .A(n_139), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_139), .A2(n_505), .B(n_506), .Y(n_504) );
CKINVDCx6p67_ASAP7_75t_R g557 ( .A(n_139), .Y(n_557) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx12f_ASAP7_75t_L g181 ( .A(n_140), .Y(n_181) );
INVx5_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_144), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_144), .B(n_591), .Y(n_590) );
INVxp67_ASAP7_75t_L g602 ( .A(n_144), .Y(n_602) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g160 ( .A(n_145), .Y(n_160) );
INVx2_ASAP7_75t_L g180 ( .A(n_145), .Y(n_180) );
INVx2_ASAP7_75t_L g245 ( .A(n_145), .Y(n_245) );
INVx2_ASAP7_75t_L g535 ( .A(n_145), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_146), .A2(n_164), .B(n_166), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_146), .A2(n_149), .B(n_173), .C(n_176), .Y(n_172) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_146), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_146), .A2(n_508), .B(n_509), .Y(n_507) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_147), .A2(n_205), .B(n_209), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_147), .A2(n_243), .B(n_247), .Y(n_242) );
OAI21x1_ASAP7_75t_L g503 ( .A1(n_147), .A2(n_504), .B(n_507), .Y(n_503) );
INVx2_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
INVx8_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_148), .A2(n_226), .B(n_593), .Y(n_592) );
INVx8_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI21x1_ASAP7_75t_SL g186 ( .A1(n_149), .A2(n_187), .B(n_194), .Y(n_186) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_149), .A2(n_218), .B(n_221), .Y(n_217) );
AOI21xp33_ASAP7_75t_L g530 ( .A1(n_149), .A2(n_227), .B(n_528), .Y(n_530) );
INVx1_ASAP7_75t_L g538 ( .A(n_149), .Y(n_538) );
INVx1_ASAP7_75t_L g605 ( .A(n_149), .Y(n_605) );
INVx1_ASAP7_75t_SL g475 ( .A(n_152), .Y(n_475) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_170), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_153), .B(n_320), .Y(n_354) );
BUFx2_ASAP7_75t_L g376 ( .A(n_153), .Y(n_376) );
AND2x2_ASAP7_75t_L g391 ( .A(n_153), .B(n_234), .Y(n_391) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g285 ( .A(n_154), .Y(n_285) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g239 ( .A(n_155), .Y(n_239) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_168), .Y(n_155) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_156), .A2(n_172), .B(n_182), .Y(n_171) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_156), .A2(n_242), .B(n_251), .Y(n_241) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_156), .A2(n_264), .B(n_271), .Y(n_263) );
INVx2_ASAP7_75t_L g489 ( .A(n_156), .Y(n_489) );
NOR2x1p5_ASAP7_75t_SL g604 ( .A(n_156), .B(n_605), .Y(n_604) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_163), .B(n_167), .Y(n_157) );
INVx2_ASAP7_75t_L g518 ( .A(n_162), .Y(n_518) );
INVx2_ASAP7_75t_L g568 ( .A(n_162), .Y(n_568) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_167), .A2(n_265), .B(n_268), .Y(n_264) );
AO31x2_ASAP7_75t_L g488 ( .A1(n_167), .A2(n_489), .A3(n_490), .B(n_499), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_167), .A2(n_554), .B(n_558), .Y(n_553) );
OAI21x1_ASAP7_75t_SL g564 ( .A1(n_167), .A2(n_565), .B(n_570), .Y(n_564) );
AND2x2_ASAP7_75t_L g396 ( .A(n_170), .B(n_202), .Y(n_396) );
AND2x2_ASAP7_75t_L g472 ( .A(n_170), .B(n_298), .Y(n_472) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_185), .Y(n_170) );
INVx3_ASAP7_75t_L g234 ( .A(n_171), .Y(n_234) );
INVx2_ASAP7_75t_L g296 ( .A(n_171), .Y(n_296) );
AND2x2_ASAP7_75t_L g311 ( .A(n_171), .B(n_257), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_181), .Y(n_176) );
INVx5_ASAP7_75t_L g207 ( .A(n_178), .Y(n_207) );
OR2x2_ASAP7_75t_L g587 ( .A(n_178), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_181), .A2(n_195), .B(n_197), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_181), .A2(n_491), .B1(n_494), .B2(n_496), .Y(n_490) );
BUFx2_ASAP7_75t_L g521 ( .A(n_181), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_181), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_181), .B(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g569 ( .A(n_181), .Y(n_569) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_183), .A2(n_186), .B(n_198), .Y(n_185) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_183), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_183), .B(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g552 ( .A(n_183), .Y(n_552) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
INVx3_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .C(n_193), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_189), .A2(n_518), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g192 ( .A(n_190), .Y(n_192) );
INVx2_ASAP7_75t_L g212 ( .A(n_192), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_193), .A2(n_219), .B(n_220), .Y(n_218) );
O2A1O1Ixp5_ASAP7_75t_L g247 ( .A1(n_193), .A2(n_248), .B(n_249), .C(n_250), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_193), .A2(n_269), .B(n_270), .Y(n_268) );
OAI21xp33_ASAP7_75t_L g532 ( .A1(n_193), .A2(n_533), .B(n_537), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_193), .A2(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g573 ( .A(n_193), .Y(n_573) );
INVx2_ASAP7_75t_L g524 ( .A(n_196), .Y(n_524) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x6_ASAP7_75t_L g430 ( .A(n_201), .B(n_431), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g473 ( .A1(n_201), .A2(n_296), .A3(n_300), .B1(n_474), .B2(n_475), .B3(n_476), .Y(n_473) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_202), .B(n_367), .Y(n_420) );
INVx1_ASAP7_75t_L g443 ( .A(n_202), .Y(n_443) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_215), .Y(n_202) );
AND2x2_ASAP7_75t_L g230 ( .A(n_203), .B(n_216), .Y(n_230) );
BUFx2_ASAP7_75t_L g366 ( .A(n_203), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_213), .B(n_214), .Y(n_203) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_204), .A2(n_213), .B(n_214), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_207), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_207), .A2(n_497), .B1(n_598), .B2(n_599), .Y(n_597) );
OAI21x1_ASAP7_75t_L g502 ( .A1(n_213), .A2(n_503), .B(n_510), .Y(n_502) );
OAI21x1_ASAP7_75t_SL g563 ( .A1(n_213), .A2(n_564), .B(n_574), .Y(n_563) );
AND2x2_ASAP7_75t_L g253 ( .A(n_215), .B(n_233), .Y(n_253) );
INVx1_ASAP7_75t_L g291 ( .A(n_215), .Y(n_291) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_215), .Y(n_310) );
NOR2xp67_ASAP7_75t_L g347 ( .A(n_215), .B(n_288), .Y(n_347) );
INVx1_ASAP7_75t_L g364 ( .A(n_215), .Y(n_364) );
INVx1_ASAP7_75t_L g393 ( .A(n_215), .Y(n_393) );
AND2x2_ASAP7_75t_L g404 ( .A(n_215), .B(n_357), .Y(n_404) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_224), .A2(n_244), .B(n_246), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_224), .A2(n_266), .B(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_224), .A2(n_601), .B(n_602), .C(n_603), .Y(n_600) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_227), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_227), .B(n_585), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_235), .B1(n_240), .B2(n_252), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_230), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g327 ( .A(n_230), .Y(n_327) );
AND2x2_ASAP7_75t_L g355 ( .A(n_230), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g381 ( .A(n_230), .B(n_314), .Y(n_381) );
AND2x2_ASAP7_75t_L g418 ( .A(n_230), .B(n_329), .Y(n_418) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_232), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g288 ( .A(n_233), .Y(n_288) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_233), .Y(n_314) );
AND2x2_ASAP7_75t_L g329 ( .A(n_233), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_SL g357 ( .A(n_233), .Y(n_357) );
INVx1_ASAP7_75t_L g367 ( .A(n_233), .Y(n_367) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_233), .Y(n_409) );
AND2x2_ASAP7_75t_L g256 ( .A(n_234), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g330 ( .A(n_234), .Y(n_330) );
AND2x2_ASAP7_75t_L g356 ( .A(n_234), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g340 ( .A(n_236), .B(n_321), .Y(n_340) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g446 ( .A(n_237), .B(n_274), .Y(n_446) );
INVx1_ASAP7_75t_L g459 ( .A(n_237), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx2_ASAP7_75t_L g383 ( .A(n_238), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_238), .B(n_275), .Y(n_428) );
BUFx2_ASAP7_75t_L g453 ( .A(n_238), .Y(n_453) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g350 ( .A(n_240), .Y(n_350) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g279 ( .A(n_241), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x4_ASAP7_75t_L g297 ( .A(n_253), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g304 ( .A(n_253), .Y(n_304) );
AND2x2_ASAP7_75t_L g445 ( .A(n_253), .B(n_410), .Y(n_445) );
AND2x2_ASAP7_75t_L g467 ( .A(n_253), .B(n_295), .Y(n_467) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x6_ASAP7_75t_L g449 ( .A(n_255), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g346 ( .A(n_256), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g440 ( .A(n_256), .B(n_404), .Y(n_440) );
AND2x4_ASAP7_75t_L g290 ( .A(n_257), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g298 ( .A(n_257), .Y(n_298) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVxp67_ASAP7_75t_R g410 ( .A(n_258), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_259), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g470 ( .A(n_259), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_260), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_260), .B(n_318), .Y(n_387) );
AOI322xp5_ASAP7_75t_L g388 ( .A1(n_260), .A2(n_342), .A3(n_389), .B1(n_392), .B2(n_394), .C1(n_396), .C2(n_397), .Y(n_388) );
INVx1_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
AND2x2_ASAP7_75t_L g307 ( .A(n_262), .B(n_278), .Y(n_307) );
INVx1_ASAP7_75t_L g344 ( .A(n_262), .Y(n_344) );
AND2x2_ASAP7_75t_L g361 ( .A(n_262), .B(n_279), .Y(n_361) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AOI21xp33_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_281), .B(n_286), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_273), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
OR2x2_ASAP7_75t_L g353 ( .A(n_274), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g439 ( .A(n_274), .B(n_361), .Y(n_439) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g326 ( .A(n_275), .B(n_301), .Y(n_326) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g282 ( .A(n_277), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g432 ( .A(n_277), .B(n_376), .Y(n_432) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g305 ( .A(n_284), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g325 ( .A(n_284), .B(n_326), .Y(n_325) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_284), .B(n_360), .Y(n_359) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_284), .B(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g318 ( .A(n_285), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g397 ( .A(n_285), .B(n_350), .Y(n_397) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
OR2x2_ASAP7_75t_L g423 ( .A(n_287), .B(n_309), .Y(n_423) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g474 ( .A(n_290), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_299), .B(n_302), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g303 ( .A(n_295), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g442 ( .A(n_295), .B(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_296), .B(n_364), .Y(n_395) );
INVx2_ASAP7_75t_L g386 ( .A(n_298), .Y(n_386) );
BUFx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g425 ( .A(n_300), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_300), .B(n_453), .Y(n_452) );
NAND2xp67_ASAP7_75t_SL g476 ( .A(n_300), .B(n_383), .Y(n_476) );
OAI222xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_305), .B2(n_308), .C1(n_315), .C2(n_317), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_305), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g417 ( .A(n_306), .Y(n_417) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g377 ( .A(n_307), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
BUFx3_ASAP7_75t_L g332 ( .A(n_309), .Y(n_332) );
NAND2x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g403 ( .A(n_311), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND2x1_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_318), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g463 ( .A(n_318), .B(n_412), .Y(n_463) );
INVx1_ASAP7_75t_L g469 ( .A(n_318), .Y(n_469) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_348), .C(n_368), .Y(n_322) );
AOI322xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .A3(n_328), .B1(n_331), .B2(n_333), .C1(n_338), .C2(n_346), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_325), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g412 ( .A(n_326), .Y(n_412) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_326), .Y(n_426) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g438 ( .A(n_329), .B(n_390), .Y(n_438) );
AND2x2_ASAP7_75t_L g363 ( .A(n_330), .B(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_332), .A2(n_449), .B1(n_452), .B2(n_454), .Y(n_451) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g400 ( .A1(n_340), .A2(n_401), .B1(n_403), .B2(n_405), .C1(n_407), .C2(n_411), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_342), .B(n_383), .Y(n_406) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g382 ( .A(n_343), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_346), .A2(n_349), .B1(n_352), .B2(n_355), .C(n_358), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g437 ( .A(n_351), .B(n_361), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_354), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g471 ( .A(n_354), .Y(n_471) );
INVx2_ASAP7_75t_L g431 ( .A(n_356), .Y(n_431) );
AND2x2_ASAP7_75t_L g456 ( .A(n_356), .B(n_410), .Y(n_456) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g372 ( .A(n_361), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g464 ( .A(n_361), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_363), .Y(n_369) );
AND2x4_ASAP7_75t_L g407 ( .A(n_363), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx2_ASAP7_75t_L g390 ( .A(n_366), .Y(n_390) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_366), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_379), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx2_ASAP7_75t_L g434 ( .A(n_377), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B1(n_384), .B2(n_387), .C(n_388), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_383), .A2(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_393), .B(n_409), .Y(n_450) );
INVx1_ASAP7_75t_L g402 ( .A(n_396), .Y(n_402) );
INVxp67_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_399), .B(n_435), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_413), .C(n_421), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_412), .B(n_459), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_418), .C(n_419), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_420), .B(n_434), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B1(n_429), .B2(n_432), .C(n_433), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .C(n_427), .Y(n_424) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g465 ( .A(n_428), .Y(n_465) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
NAND4xp25_ASAP7_75t_SL g435 ( .A(n_436), .B(n_447), .C(n_455), .D(n_466), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_439), .B2(n_440), .C(n_441), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .B(n_446), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_460), .B2(n_463), .C1(n_464), .C2(n_891), .Y(n_455) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_470), .B2(n_472), .C(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NOR2x1p5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NOR2x1p5_ASAP7_75t_L g481 ( .A(n_482), .B(n_757), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_710), .Y(n_482) );
NOR4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_621), .C(n_652), .D(n_686), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_544), .B(n_612), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AOI322xp5_ASAP7_75t_L g724 ( .A1(n_486), .A2(n_613), .A3(n_635), .B1(n_725), .B2(n_726), .C1(n_727), .C2(n_728), .Y(n_724) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_511), .Y(n_486) );
INVx1_ASAP7_75t_L g669 ( .A(n_487), .Y(n_669) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_501), .Y(n_487) );
INVx2_ASAP7_75t_L g617 ( .A(n_488), .Y(n_617) );
INVx2_ASAP7_75t_SL g633 ( .A(n_488), .Y(n_633) );
AND2x2_ASAP7_75t_L g638 ( .A(n_488), .B(n_639), .Y(n_638) );
AND2x4_ASAP7_75t_L g662 ( .A(n_488), .B(n_618), .Y(n_662) );
INVx1_ASAP7_75t_L g678 ( .A(n_488), .Y(n_678) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_497), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_533) );
AND2x2_ASAP7_75t_L g636 ( .A(n_501), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g681 ( .A(n_501), .Y(n_681) );
AND2x2_ASAP7_75t_L g697 ( .A(n_501), .B(n_665), .Y(n_697) );
AND2x2_ASAP7_75t_L g709 ( .A(n_501), .B(n_531), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_501), .B(n_651), .Y(n_764) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_501), .Y(n_814) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g618 ( .A(n_502), .Y(n_618) );
BUFx3_ASAP7_75t_L g797 ( .A(n_511), .Y(n_797) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_531), .Y(n_511) );
OR2x2_ASAP7_75t_L g620 ( .A(n_512), .B(n_531), .Y(n_620) );
INVx2_ASAP7_75t_L g631 ( .A(n_512), .Y(n_631) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g637 ( .A(n_513), .Y(n_637) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_522), .B(n_530), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_519), .B(n_521), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_527), .B(n_528), .Y(n_522) );
AO21x1_ASAP7_75t_L g580 ( .A1(n_527), .A2(n_581), .B(n_584), .Y(n_580) );
AOI21x1_ASAP7_75t_L g586 ( .A1(n_527), .A2(n_587), .B(n_589), .Y(n_586) );
AND2x4_ASAP7_75t_L g632 ( .A(n_531), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g639 ( .A(n_531), .Y(n_639) );
INVx2_ASAP7_75t_SL g665 ( .A(n_531), .Y(n_665) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_531), .Y(n_668) );
AND2x2_ASAP7_75t_L g785 ( .A(n_531), .B(n_631), .Y(n_785) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_539), .B(n_543), .Y(n_531) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_606), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_546), .B(n_575), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_546), .B(n_677), .C(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g808 ( .A(n_547), .B(n_774), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_547), .B(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_562), .Y(n_548) );
INVx2_ASAP7_75t_L g646 ( .A(n_549), .Y(n_646) );
AND2x2_ASAP7_75t_L g703 ( .A(n_549), .B(n_609), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_549), .B(n_594), .Y(n_750) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g625 ( .A(n_550), .Y(n_625) );
OAI21x1_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_553), .B(n_561), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_557), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_557), .A2(n_597), .B(n_600), .C(n_604), .Y(n_596) );
AND2x4_ASAP7_75t_L g691 ( .A(n_562), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g701 ( .A(n_562), .B(n_594), .Y(n_701) );
INVx1_ASAP7_75t_L g756 ( .A(n_562), .Y(n_756) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx3_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
AOI21x1_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B(n_569), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B(n_573), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_575), .A2(n_824), .B1(n_826), .B2(n_827), .C(n_829), .Y(n_823) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g815 ( .A(n_576), .B(n_644), .Y(n_815) );
AND2x2_ASAP7_75t_L g831 ( .A(n_576), .B(n_703), .Y(n_831) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_594), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_577), .B(n_611), .Y(n_614) );
INVx2_ASAP7_75t_L g723 ( .A(n_577), .Y(n_723) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_578), .Y(n_706) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g608 ( .A(n_579), .Y(n_608) );
BUFx3_ASAP7_75t_L g643 ( .A(n_579), .Y(n_643) );
OAI21x1_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_586), .B(n_592), .Y(n_579) );
INVxp67_ASAP7_75t_L g593 ( .A(n_584), .Y(n_593) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g611 ( .A(n_594), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_594), .B(n_608), .Y(n_648) );
INVx1_ASAP7_75t_L g656 ( .A(n_594), .Y(n_656) );
INVx1_ASAP7_75t_L g692 ( .A(n_594), .Y(n_692) );
HB1xp67_ASAP7_75t_SL g716 ( .A(n_594), .Y(n_716) );
INVx1_ASAP7_75t_L g754 ( .A(n_594), .Y(n_754) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_606), .A2(n_613), .B(n_615), .Y(n_612) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_607), .B(n_610), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g655 ( .A(n_608), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g734 ( .A(n_608), .Y(n_734) );
INVx2_ASAP7_75t_L g626 ( .A(n_609), .Y(n_626) );
AND2x4_ASAP7_75t_L g644 ( .A(n_609), .B(n_624), .Y(n_644) );
BUFx2_ASAP7_75t_L g658 ( .A(n_609), .Y(n_658) );
AND2x2_ASAP7_75t_L g721 ( .A(n_609), .B(n_611), .Y(n_721) );
INVx1_ASAP7_75t_L g727 ( .A(n_610), .Y(n_727) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g672 ( .A(n_611), .B(n_624), .Y(n_672) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g782 ( .A(n_614), .B(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
AND2x4_ASAP7_75t_SL g649 ( .A(n_616), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_616), .B(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_SL g718 ( .A(n_616), .B(n_664), .Y(n_718) );
AOI32xp33_ASAP7_75t_L g767 ( .A1(n_616), .A2(n_629), .A3(n_745), .B1(n_768), .B2(n_769), .Y(n_767) );
INVxp67_ASAP7_75t_L g798 ( .A(n_616), .Y(n_798) );
AND2x4_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x4_ASAP7_75t_L g708 ( .A(n_617), .B(n_631), .Y(n_708) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_618), .Y(n_628) );
AND2x4_ASAP7_75t_L g736 ( .A(n_619), .B(n_662), .Y(n_736) );
AND2x4_ASAP7_75t_L g739 ( .A(n_619), .B(n_628), .Y(n_739) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g802 ( .A(n_620), .B(n_641), .Y(n_802) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_627), .B(n_634), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_622), .B(n_722), .Y(n_809) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI31xp33_ASAP7_75t_L g702 ( .A1(n_623), .A2(n_703), .A3(n_704), .B(n_707), .Y(n_702) );
OR4x1_ASAP7_75t_L g763 ( .A(n_623), .B(n_764), .C(n_765), .D(n_766), .Y(n_763) );
AND2x2_ASAP7_75t_L g768 ( .A(n_623), .B(n_722), .Y(n_768) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g700 ( .A(n_624), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_624), .B(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g783 ( .A(n_624), .Y(n_783) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g659 ( .A(n_625), .B(n_643), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g741 ( .A(n_628), .B(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g792 ( .A(n_628), .Y(n_792) );
AND2x2_ASAP7_75t_L g830 ( .A(n_628), .B(n_664), .Y(n_830) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g685 ( .A(n_630), .Y(n_685) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g725 ( .A(n_632), .B(n_636), .Y(n_725) );
INVx2_ASAP7_75t_L g742 ( .A(n_632), .Y(n_742) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_632), .Y(n_751) );
AND2x2_ASAP7_75t_L g828 ( .A(n_632), .B(n_685), .Y(n_828) );
INVx1_ASAP7_75t_L g696 ( .A(n_633), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_640), .B1(n_645), .B2(n_649), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx2_ASAP7_75t_L g651 ( .A(n_637), .Y(n_651) );
AND2x2_ASAP7_75t_L g664 ( .A(n_637), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g675 ( .A(n_637), .B(n_642), .Y(n_675) );
INVx1_ASAP7_75t_L g765 ( .A(n_638), .Y(n_765) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
AND2x2_ASAP7_75t_L g745 ( .A(n_641), .B(n_691), .Y(n_745) );
AND2x2_ASAP7_75t_L g762 ( .A(n_641), .B(n_721), .Y(n_762) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_644), .A2(n_674), .B1(n_676), .B2(n_682), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_644), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g726 ( .A(n_644), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_644), .B(n_683), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_645), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_737) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x4_ASAP7_75t_L g654 ( .A(n_646), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g693 ( .A(n_646), .Y(n_693) );
AND2x2_ASAP7_75t_L g775 ( .A(n_646), .B(n_701), .Y(n_775) );
INVx1_ASAP7_75t_L g800 ( .A(n_646), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_647), .B(n_703), .Y(n_788) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g795 ( .A(n_648), .Y(n_795) );
INVx1_ASAP7_75t_L g769 ( .A(n_650), .Y(n_769) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_651), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g771 ( .A(n_651), .B(n_696), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_660), .B1(n_666), .B2(n_670), .C(n_673), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
INVx2_ASAP7_75t_L g683 ( .A(n_655), .Y(n_683) );
AOI322xp5_ASAP7_75t_L g804 ( .A1(n_657), .A2(n_661), .A3(n_713), .B1(n_805), .B2(n_807), .C1(n_808), .C2(n_809), .Y(n_804) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x4_ASAP7_75t_L g671 ( .A(n_658), .B(n_672), .Y(n_671) );
OR2x6_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g714 ( .A(n_662), .B(n_667), .Y(n_714) );
AND2x2_ASAP7_75t_L g784 ( .A(n_662), .B(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_662), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g821 ( .A(n_662), .Y(n_821) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g791 ( .A(n_664), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g761 ( .A(n_666), .Y(n_761) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g688 ( .A(n_668), .Y(n_688) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI31xp33_ASAP7_75t_L g786 ( .A1(n_671), .A2(n_787), .A3(n_789), .B(n_791), .Y(n_786) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_672), .Y(n_728) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g684 ( .A(n_677), .Y(n_684) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g713 ( .A(n_680), .B(n_708), .Y(n_713) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .C(n_685), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_694), .B2(n_698), .C(n_702), .Y(n_686) );
INVx1_ASAP7_75t_L g746 ( .A(n_687), .Y(n_746) );
OR2x2_ASAP7_75t_L g820 ( .A(n_688), .B(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_690), .B(n_723), .Y(n_776) );
AND2x4_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
BUFx2_ASAP7_75t_L g780 ( .A(n_691), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
AND2x2_ASAP7_75t_L g807 ( .A(n_697), .B(n_708), .Y(n_807) );
AND2x4_ASAP7_75t_L g833 ( .A(n_697), .B(n_771), .Y(n_833) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g735 ( .A(n_701), .Y(n_735) );
BUFx2_ASAP7_75t_L g832 ( .A(n_703), .Y(n_832) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g790 ( .A(n_705), .B(n_735), .Y(n_790) );
INVx1_ASAP7_75t_L g774 ( .A(n_706), .Y(n_774) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_708), .B(n_709), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_729), .C(n_743), .Y(n_710) );
OAI221xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_724), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_713), .A2(n_748), .B1(n_751), .B2(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OR2x6_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g749 ( .A(n_723), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_726), .B(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_737), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_736), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g766 ( .A(n_733), .Y(n_766) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_734), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g818 ( .A(n_734), .Y(n_818) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_744), .B(n_747), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NAND4xp75_ASAP7_75t_L g757 ( .A(n_758), .B(n_777), .C(n_803), .D(n_822), .Y(n_757) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_770), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_763), .C(n_767), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g826 ( .A(n_775), .Y(n_826) );
NOR2x1_ASAP7_75t_L g777 ( .A(n_778), .B(n_793), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_786), .Y(n_778) );
OAI21xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B(n_784), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g806 ( .A(n_785), .Y(n_806) );
AND2x2_ASAP7_75t_L g825 ( .A(n_785), .B(n_792), .Y(n_825) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_796), .B1(n_798), .B2(n_799), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_797), .B(n_813), .Y(n_812) );
NAND2x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_810), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_815), .B1(n_816), .B2(n_819), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_829) );
INVxp67_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_839), .Y(n_838) );
OR2x6_ASAP7_75t_L g839 ( .A(n_840), .B(n_842), .Y(n_839) );
OR2x2_ASAP7_75t_L g860 ( .A(n_840), .B(n_861), .Y(n_860) );
BUFx2_ASAP7_75t_L g871 ( .A(n_840), .Y(n_871) );
INVx2_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g867 ( .A(n_842), .Y(n_867) );
AND2x4_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
NOR3xp33_ASAP7_75t_L g883 ( .A(n_843), .B(n_884), .C(n_887), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_868), .B(n_870), .Y(n_845) );
AOI21xp33_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_856), .B(n_857), .Y(n_846) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_847), .Y(n_869) );
AOI22x1_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_850), .B1(n_853), .B2(n_855), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_SL g855 ( .A(n_850), .Y(n_855) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_857), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B(n_862), .Y(n_857) );
BUFx12f_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g872 ( .A(n_862), .Y(n_872) );
INVx3_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
BUFx6f_ASAP7_75t_L g876 ( .A(n_865), .Y(n_876) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
BUFx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_879), .Y(n_878) );
INVx6_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_880), .Y(n_889) );
AND2x4_ASAP7_75t_L g880 ( .A(n_881), .B(n_883), .Y(n_880) );
INVx4_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
endmodule