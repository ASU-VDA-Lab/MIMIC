module fake_jpeg_30119_n_216 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_165;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_17),
.B(n_1),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_57),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_17),
.B(n_2),
.Y(n_58)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_31),
.B1(n_33),
.B2(n_22),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_81),
.B1(n_87),
.B2(n_48),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_22),
.B1(n_33),
.B2(n_18),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_80),
.B1(n_89),
.B2(n_24),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_6),
.C(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_10),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_32),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_36),
.B1(n_31),
.B2(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_7),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_85),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_43),
.A2(n_36),
.B1(n_50),
.B2(n_46),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_30),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_110),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_16),
.B(n_24),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_96),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_9),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_99),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_39),
.A3(n_56),
.B1(n_53),
.B2(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_63),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_47),
.B(n_38),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_85),
.B(n_63),
.C(n_68),
.Y(n_125)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_53),
.B1(n_48),
.B2(n_44),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_111),
.B1(n_87),
.B2(n_89),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_112),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_56),
.C(n_44),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_124),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_113),
.B1(n_111),
.B2(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_82),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_77),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_108),
.C(n_83),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_108),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_144),
.B1(n_130),
.B2(n_135),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_108),
.B1(n_83),
.B2(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_91),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_103),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_140),
.B(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_154),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_116),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_92),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_159),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_138),
.B(n_135),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_167),
.B(n_152),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_172),
.B1(n_141),
.B2(n_143),
.C(n_151),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_138),
.B(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_131),
.B1(n_130),
.B2(n_123),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_125),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_158),
.C(n_142),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_182),
.C(n_175),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_142),
.B1(n_141),
.B2(n_144),
.C(n_150),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_185),
.B(n_186),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_156),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_165),
.C(n_163),
.Y(n_182)
);

OAI322xp33_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_147),
.A3(n_146),
.B1(n_145),
.B2(n_121),
.C1(n_129),
.C2(n_12),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_121),
.B1(n_133),
.B2(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_12),
.C(n_133),
.Y(n_185)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_129),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_191),
.C(n_194),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_175),
.C(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_174),
.C(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_170),
.C(n_164),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_198),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_190),
.B1(n_186),
.B2(n_196),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_126),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_200),
.B1(n_184),
.B2(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_206),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_126),
.Y(n_206)
);

OAI221xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.C(n_98),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_78),
.B(n_86),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_66),
.B(n_104),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_211),
.B(n_68),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_78),
.B(n_86),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_213),
.C(n_210),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_68),
.Y(n_216)
);


endmodule