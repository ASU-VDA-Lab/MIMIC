module fake_jpeg_8138_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_42),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_18),
.B1(n_22),
.B2(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_62),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_25),
.B1(n_21),
.B2(n_33),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_25),
.B1(n_36),
.B2(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_70),
.A2(n_73),
.B1(n_18),
.B2(n_22),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_29),
.B1(n_23),
.B2(n_33),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_90),
.Y(n_98)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_33),
.B1(n_36),
.B2(n_35),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_82),
.B1(n_36),
.B2(n_53),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_39),
.B1(n_34),
.B2(n_35),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_85),
.B1(n_65),
.B2(n_68),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_68),
.B1(n_54),
.B2(n_62),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_105),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_59),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_31),
.B(n_49),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_67),
.B1(n_53),
.B2(n_39),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_90),
.B1(n_89),
.B2(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_53),
.B1(n_35),
.B2(n_54),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_32),
.B1(n_93),
.B2(n_17),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_66),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_120),
.B(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_119),
.B1(n_35),
.B2(n_74),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_37),
.B1(n_52),
.B2(n_45),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_37),
.B(n_14),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_22),
.B1(n_32),
.B2(n_28),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_86),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_124),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_94),
.C(n_71),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_128),
.C(n_110),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_71),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_132),
.B1(n_135),
.B2(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_137),
.B1(n_141),
.B2(n_145),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_74),
.B1(n_84),
.B2(n_87),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_84),
.B1(n_61),
.B2(n_47),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_123),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_47),
.B1(n_87),
.B2(n_88),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_91),
.B1(n_88),
.B2(n_17),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_28),
.B1(n_24),
.B2(n_16),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_149),
.B(n_98),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_122),
.Y(n_163)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_148),
.A2(n_103),
.B1(n_107),
.B2(n_99),
.Y(n_155)
);

NOR2x1_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_101),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_166),
.B(n_167),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_111),
.B1(n_108),
.B2(n_101),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_132),
.B1(n_136),
.B2(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_127),
.B1(n_130),
.B2(n_106),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_133),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_97),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_126),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_99),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

BUFx8_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_119),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_26),
.C(n_16),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_104),
.B(n_117),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_113),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_113),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_24),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_181),
.B1(n_183),
.B2(n_186),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_149),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_145),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_136),
.B1(n_130),
.B2(n_129),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_127),
.B1(n_124),
.B2(n_103),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_24),
.B1(n_66),
.B2(n_48),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_26),
.B1(n_19),
.B2(n_92),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_26),
.B1(n_19),
.B2(n_92),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_196),
.A2(n_197),
.B(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_19),
.B1(n_31),
.B2(n_3),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_19),
.C(n_31),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_161),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_150),
.CI(n_193),
.CON(n_200),
.SN(n_200)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_200),
.B(n_204),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_167),
.B(n_153),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_211),
.B(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_152),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_160),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_207),
.C(n_208),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_154),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_174),
.B(n_164),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_220),
.C(n_1),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_174),
.C(n_172),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_190),
.B1(n_198),
.B2(n_191),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_161),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_19),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_195),
.B(n_188),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_202),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_184),
.B(n_187),
.Y(n_226)
);

OAI22x1_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_229),
.B1(n_234),
.B2(n_200),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_181),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_190),
.B1(n_196),
.B2(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_197),
.B1(n_162),
.B2(n_13),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_232),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_1),
.C(n_2),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_12),
.B1(n_2),
.B2(n_4),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_201),
.B1(n_209),
.B2(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_1),
.C(n_4),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_215),
.C(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_207),
.C(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_247),
.C(n_249),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_225),
.B1(n_226),
.B2(n_233),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_248),
.B(n_231),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_243),
.B1(n_225),
.B2(n_240),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_206),
.C(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_4),
.C(n_5),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_257),
.B(n_6),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_230),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_228),
.C(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_241),
.C(n_7),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_242),
.B1(n_237),
.B2(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_261),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_249),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_247),
.B1(n_241),
.B2(n_8),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_257),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_257),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_8),
.C2(n_253),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_257),
.C(n_9),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_263),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_265),
.B1(n_11),
.B2(n_10),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_266),
.C1(n_259),
.C2(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

OAI311xp33_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_10),
.A3(n_271),
.B1(n_245),
.C1(n_251),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_277),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_276),
.Y(n_280)
);


endmodule