module fake_jpeg_22760_n_24 (n_3, n_2, n_1, n_0, n_4, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

INVx5_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_7),
.C(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_9),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_6),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_7),
.B(n_5),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_15),
.B(n_16),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_8),
.B1(n_11),
.B2(n_0),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_18),
.B1(n_14),
.B2(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_21),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_3),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_20),
.C(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_1),
.Y(n_24)
);


endmodule