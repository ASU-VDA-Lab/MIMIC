module real_aes_8920_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g449 ( .A(n_0), .Y(n_449) );
INVx1_ASAP7_75t_L g508 ( .A(n_1), .Y(n_508) );
INVx1_ASAP7_75t_L g265 ( .A(n_2), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_3), .A2(n_39), .B1(n_184), .B2(n_536), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g172 ( .A1(n_4), .A2(n_173), .B(n_174), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_5), .B(n_171), .Y(n_485) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_7), .A2(n_105), .B1(n_114), .B2(n_756), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_8), .A2(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_9), .B(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g181 ( .A(n_10), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_11), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
INVx1_ASAP7_75t_L g504 ( .A(n_13), .Y(n_504) );
INVx1_ASAP7_75t_L g247 ( .A(n_14), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_15), .B(n_149), .Y(n_542) );
AOI222xp33_ASAP7_75t_SL g453 ( .A1(n_16), .A2(n_454), .B1(n_455), .B2(n_464), .C1(n_751), .C2(n_752), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_17), .B(n_139), .Y(n_513) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_18), .B(n_122), .Y(n_121) );
AO32x2_ASAP7_75t_L g533 ( .A1(n_18), .A2(n_138), .A3(n_171), .B1(n_496), .B2(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_19), .B(n_184), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_20), .B(n_192), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_21), .B(n_139), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_22), .A2(n_51), .B1(n_184), .B2(n_536), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_23), .B(n_173), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_24), .A2(n_78), .B1(n_149), .B2(n_184), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_25), .B(n_184), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_26), .B(n_169), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_27), .A2(n_456), .B1(n_457), .B2(n_463), .Y(n_455) );
INVx1_ASAP7_75t_L g463 ( .A(n_27), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_28), .A2(n_245), .B(n_246), .C(n_248), .Y(n_244) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_29), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_30), .B(n_186), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_31), .B(n_179), .Y(n_266) );
INVx1_ASAP7_75t_L g157 ( .A(n_32), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_33), .B(n_186), .Y(n_530) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_35), .B(n_184), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_36), .B(n_186), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_37), .A2(n_43), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_37), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_38), .A2(n_146), .B(n_158), .C(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g155 ( .A(n_41), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_42), .B(n_179), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_43), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_44), .B(n_184), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_45), .A2(n_88), .B1(n_209), .B2(n_536), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_46), .B(n_184), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_47), .B(n_184), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_48), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_49), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_50), .B(n_173), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_52), .A2(n_61), .B1(n_149), .B2(n_184), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_53), .A2(n_149), .B1(n_152), .B2(n_158), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_54), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_55), .B(n_184), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_56), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_57), .B(n_184), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_58), .A2(n_178), .B(n_180), .C(n_183), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_59), .Y(n_222) );
INVx1_ASAP7_75t_L g175 ( .A(n_60), .Y(n_175) );
INVx1_ASAP7_75t_L g147 ( .A(n_62), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_63), .B(n_184), .Y(n_509) );
INVx1_ASAP7_75t_L g142 ( .A(n_64), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
AO32x2_ASAP7_75t_L g553 ( .A1(n_66), .A2(n_171), .A3(n_227), .B1(n_496), .B2(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g493 ( .A(n_67), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_68), .A2(n_125), .B1(n_126), .B2(n_129), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_68), .Y(n_129) );
INVx1_ASAP7_75t_L g525 ( .A(n_69), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_SL g191 ( .A1(n_70), .A2(n_183), .B(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_71), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_72), .B(n_149), .Y(n_526) );
INVx1_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_74), .Y(n_166) );
INVx1_ASAP7_75t_L g215 ( .A(n_75), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_76), .A2(n_102), .B1(n_461), .B2(n_462), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_76), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_77), .B(n_451), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_79), .A2(n_146), .B(n_158), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_80), .B(n_536), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_81), .B(n_149), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_82), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_84), .B(n_192), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_85), .B(n_149), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_86), .A2(n_146), .B(n_158), .C(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g108 ( .A(n_87), .Y(n_108) );
OR2x2_ASAP7_75t_L g446 ( .A(n_87), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g467 ( .A(n_87), .B(n_448), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_89), .A2(n_103), .B1(n_149), .B2(n_150), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_90), .B(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_91), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_92), .A2(n_146), .B(n_158), .C(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_93), .Y(n_237) );
INVx1_ASAP7_75t_L g190 ( .A(n_94), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_95), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_96), .B(n_205), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_97), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_97), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_98), .B(n_149), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_99), .B(n_171), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_100), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_101), .A2(n_173), .B(n_189), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_102), .Y(n_462) );
INVx1_ASAP7_75t_SL g757 ( .A(n_105), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_112), .Y(n_106) );
OR2x2_ASAP7_75t_L g750 ( .A(n_108), .B(n_448), .Y(n_750) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_108), .B(n_447), .Y(n_751) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g448 ( .A(n_113), .B(n_449), .Y(n_448) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_452), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g755 ( .A(n_119), .Y(n_755) );
OAI21x1_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_443), .B(n_450), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_130), .B2(n_131), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_130), .A2(n_465), .B1(n_468), .B2(n_748), .Y(n_464) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_131), .A2(n_465), .B1(n_753), .B2(n_754), .Y(n_752) );
AND3x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_368), .C(n_417), .Y(n_131) );
NOR3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_275), .C(n_313), .Y(n_132) );
OAI222xp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_196), .B1(n_250), .B2(n_256), .C1(n_270), .C2(n_273), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_167), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_135), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_135), .B(n_318), .Y(n_409) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g286 ( .A(n_136), .B(n_187), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_136), .B(n_168), .Y(n_294) );
AND2x2_ASAP7_75t_L g329 ( .A(n_136), .B(n_306), .Y(n_329) );
OR2x2_ASAP7_75t_L g353 ( .A(n_136), .B(n_168), .Y(n_353) );
OR2x2_ASAP7_75t_L g361 ( .A(n_136), .B(n_260), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_136), .B(n_187), .Y(n_364) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g258 ( .A(n_137), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_137), .B(n_187), .Y(n_272) );
AND2x2_ASAP7_75t_L g322 ( .A(n_137), .B(n_260), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_137), .B(n_168), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_137), .B(n_421), .Y(n_442) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_165), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_138), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_138), .A2(n_261), .B(n_268), .Y(n_260) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_140), .B(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B1(n_161), .B2(n_162), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_145), .A2(n_175), .B(n_176), .C(n_177), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_145), .A2(n_176), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_145), .A2(n_176), .B(n_243), .C(n_244), .Y(n_242) );
INVx4_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_146), .B(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g173 ( .A(n_146), .B(n_163), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_146), .A2(n_477), .B(n_480), .Y(n_476) );
BUFx3_ASAP7_75t_L g496 ( .A(n_146), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_146), .A2(n_503), .B(n_507), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_146), .A2(n_524), .B(n_527), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_146), .A2(n_540), .B(n_544), .Y(n_539) );
INVx2_ASAP7_75t_L g267 ( .A(n_149), .Y(n_267) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx1_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g152 ( .A1(n_153), .A2(n_155), .B1(n_156), .B2(n_157), .Y(n_152) );
INVx2_ASAP7_75t_L g156 ( .A(n_153), .Y(n_156) );
INVx4_ASAP7_75t_L g245 ( .A(n_153), .Y(n_245) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
AND2x2_ASAP7_75t_L g163 ( .A(n_154), .B(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx3_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx5_ASAP7_75t_L g176 ( .A(n_158), .Y(n_176) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
BUFx3_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
INVx1_ASAP7_75t_L g536 ( .A(n_159), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_162), .A2(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_162), .A2(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g483 ( .A(n_164), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_167), .A2(n_361), .B(n_362), .C(n_365), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_167), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_167), .B(n_305), .Y(n_427) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_187), .Y(n_167) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_168), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g285 ( .A(n_168), .Y(n_285) );
AND2x2_ASAP7_75t_L g312 ( .A(n_168), .B(n_306), .Y(n_312) );
INVx1_ASAP7_75t_SL g320 ( .A(n_168), .Y(n_320) );
AND2x2_ASAP7_75t_L g343 ( .A(n_168), .B(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g421 ( .A(n_168), .Y(n_421) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_185), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_170), .B(n_212), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_170), .B(n_496), .C(n_515), .Y(n_514) );
AO21x1_ASAP7_75t_L g559 ( .A1(n_170), .A2(n_515), .B(n_560), .Y(n_559) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_171), .A2(n_188), .B(n_195), .Y(n_187) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_171), .A2(n_476), .B(n_485), .Y(n_475) );
BUFx2_ASAP7_75t_L g241 ( .A(n_173), .Y(n_241) );
O2A1O1Ixp5_ASAP7_75t_L g492 ( .A1(n_178), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_178), .A2(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_179), .A2(n_484), .B1(n_516), .B2(n_517), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_179), .A2(n_484), .B1(n_535), .B2(n_537), .Y(n_534) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_179), .A2(n_182), .B1(n_555), .B2(n_556), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_182), .B(n_194), .Y(n_193) );
INVx5_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
O2A1O1Ixp5_ASAP7_75t_SL g524 ( .A1(n_183), .A2(n_205), .B(n_525), .C(n_526), .Y(n_524) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
INVx1_ASAP7_75t_L g223 ( .A(n_186), .Y(n_223) );
INVx2_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_186), .A2(n_240), .B(n_249), .Y(n_239) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_186), .A2(n_523), .B(n_530), .Y(n_522) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_186), .A2(n_539), .B(n_547), .Y(n_538) );
BUFx2_ASAP7_75t_L g257 ( .A(n_187), .Y(n_257) );
INVx1_ASAP7_75t_L g319 ( .A(n_187), .Y(n_319) );
INVx3_ASAP7_75t_L g344 ( .A(n_187), .Y(n_344) );
INVx1_ASAP7_75t_L g543 ( .A(n_192), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_196), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_224), .Y(n_196) );
INVx1_ASAP7_75t_L g340 ( .A(n_197), .Y(n_340) );
OAI32xp33_ASAP7_75t_L g346 ( .A1(n_197), .A2(n_285), .A3(n_347), .B1(n_348), .B2(n_349), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_197), .A2(n_351), .B1(n_354), .B2(n_359), .Y(n_350) );
INVx4_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g288 ( .A(n_198), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g366 ( .A(n_198), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g436 ( .A(n_198), .B(n_382), .Y(n_436) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
AND2x2_ASAP7_75t_L g251 ( .A(n_199), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g281 ( .A(n_199), .Y(n_281) );
INVx1_ASAP7_75t_L g300 ( .A(n_199), .Y(n_300) );
OR2x2_ASAP7_75t_L g308 ( .A(n_199), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_199), .B(n_289), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_199), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g336 ( .A(n_199), .B(n_254), .Y(n_336) );
INVx3_ASAP7_75t_L g358 ( .A(n_199), .Y(n_358) );
AND2x2_ASAP7_75t_L g383 ( .A(n_199), .B(n_255), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_199), .B(n_348), .Y(n_431) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_211), .Y(n_199) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_202), .B(n_210), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B(n_207), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_205), .A2(n_265), .B(n_266), .C(n_267), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_205), .A2(n_478), .B(n_479), .Y(n_477) );
INVx2_ASAP7_75t_L g484 ( .A(n_205), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_205), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_207), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
INVx1_ASAP7_75t_L g220 ( .A(n_210), .Y(n_220) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_210), .A2(n_488), .B(n_497), .Y(n_487) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_210), .A2(n_502), .B(n_510), .Y(n_501) );
INVx2_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
AND2x2_ASAP7_75t_L g387 ( .A(n_213), .B(n_225), .Y(n_387) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_223), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_223), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g429 ( .A(n_224), .Y(n_429) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_238), .Y(n_224) );
INVx1_ASAP7_75t_L g274 ( .A(n_225), .Y(n_274) );
AND2x2_ASAP7_75t_L g301 ( .A(n_225), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_225), .B(n_255), .Y(n_309) );
AND2x2_ASAP7_75t_L g367 ( .A(n_225), .B(n_290), .Y(n_367) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g253 ( .A(n_226), .Y(n_253) );
AND2x2_ASAP7_75t_L g280 ( .A(n_226), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g289 ( .A(n_226), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_226), .B(n_255), .Y(n_355) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_236), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_234), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_238), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_238), .B(n_255), .Y(n_348) );
AND2x2_ASAP7_75t_L g357 ( .A(n_238), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g382 ( .A(n_238), .Y(n_382) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g254 ( .A(n_239), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g290 ( .A(n_239), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_245), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g506 ( .A(n_245), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_245), .A2(n_528), .B(n_529), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_250), .A2(n_260), .B1(n_419), .B2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_252), .A2(n_363), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_253), .B(n_358), .Y(n_375) );
INVx1_ASAP7_75t_L g400 ( .A(n_253), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_254), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g327 ( .A(n_254), .B(n_280), .Y(n_327) );
INVx2_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
INVx1_ASAP7_75t_L g333 ( .A(n_255), .Y(n_333) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_256), .A2(n_408), .B1(n_425), .B2(n_428), .C(n_430), .Y(n_424) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_257), .B(n_306), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_258), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g349 ( .A(n_258), .B(n_295), .Y(n_349) );
INVx3_ASAP7_75t_SL g390 ( .A(n_258), .Y(n_390) );
AND2x2_ASAP7_75t_L g334 ( .A(n_259), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g363 ( .A(n_259), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_259), .B(n_272), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_259), .B(n_318), .Y(n_404) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g306 ( .A(n_260), .Y(n_306) );
OAI322xp33_ASAP7_75t_L g401 ( .A1(n_260), .A2(n_332), .A3(n_354), .B1(n_402), .B2(n_404), .C1(n_405), .C2(n_406), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_267), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_271), .A2(n_274), .B(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_272), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g373 ( .A(n_272), .B(n_285), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_272), .B(n_312), .Y(n_388) );
INVxp67_ASAP7_75t_L g339 ( .A(n_274), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_274), .A2(n_346), .B(n_350), .C(n_360), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_284), .B1(n_287), .B2(n_291), .C(n_296), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g299 ( .A(n_283), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g416 ( .A(n_283), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_284), .A2(n_433), .B1(n_438), .B2(n_439), .C(n_441), .Y(n_432) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g332 ( .A(n_285), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_285), .B(n_363), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_285), .B(n_390), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_286), .B(n_311), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_286), .A2(n_298), .B1(n_408), .B2(n_409), .Y(n_407) );
OR2x2_ASAP7_75t_L g438 ( .A(n_286), .B(n_306), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g415 ( .A(n_289), .Y(n_415) );
AND2x2_ASAP7_75t_L g440 ( .A(n_289), .B(n_383), .Y(n_440) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g304 ( .A(n_294), .B(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_303), .B1(n_307), .B2(n_310), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g371 ( .A(n_299), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_299), .B(n_339), .Y(n_406) );
AOI322xp5_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_331), .A3(n_333), .B1(n_334), .B2(n_336), .C1(n_337), .C2(n_341), .Y(n_330) );
INVxp67_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_304), .A2(n_309), .B1(n_326), .B2(n_328), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_305), .B(n_318), .Y(n_405) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_306), .B(n_344), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_306), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g402 ( .A(n_308), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NAND3xp33_ASAP7_75t_SL g313 ( .A(n_314), .B(n_330), .C(n_345), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_321), .B2(n_323), .C(n_325), .Y(n_314) );
AND2x2_ASAP7_75t_L g321 ( .A(n_317), .B(n_322), .Y(n_321) );
INVx3_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_324), .Y(n_403) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_329), .B(n_343), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_332), .B(n_390), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_333), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g408 ( .A(n_336), .Y(n_408) );
AND2x2_ASAP7_75t_L g423 ( .A(n_336), .B(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_347), .A2(n_418), .B(n_424), .C(n_432), .Y(n_417) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g386 ( .A(n_357), .B(n_387), .Y(n_386) );
NAND2x1_ASAP7_75t_SL g428 ( .A(n_358), .B(n_429), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g393 ( .A(n_367), .Y(n_393) );
AND2x2_ASAP7_75t_L g397 ( .A(n_367), .B(n_383), .Y(n_397) );
NOR5xp2_ASAP7_75t_L g368 ( .A(n_369), .B(n_384), .C(n_401), .D(n_407), .E(n_410), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_372), .B2(n_374), .C(n_376), .Y(n_369) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_373), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g399 ( .A(n_383), .B(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_388), .B1(n_389), .B2(n_391), .C(n_394), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
AOI211xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_413), .B(n_415), .C(n_416), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
CKINVDCx14_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g451 ( .A(n_446), .Y(n_451) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_450), .B(n_453), .C(n_755), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
CKINVDCx14_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g753 ( .A(n_468), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_469), .B(n_672), .Y(n_468) );
AND2x2_ASAP7_75t_SL g469 ( .A(n_470), .B(n_630), .Y(n_469) );
NOR4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_570), .C(n_606), .D(n_620), .Y(n_470) );
OAI221xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_518), .B1(n_548), .B2(n_557), .C(n_561), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_472), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_498), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_486), .Y(n_474) );
AND2x2_ASAP7_75t_L g567 ( .A(n_475), .B(n_487), .Y(n_567) );
INVx3_ASAP7_75t_L g575 ( .A(n_475), .Y(n_575) );
AND2x2_ASAP7_75t_L g629 ( .A(n_475), .B(n_501), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_475), .B(n_500), .Y(n_665) );
AND2x2_ASAP7_75t_L g723 ( .A(n_475), .B(n_585), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_484), .Y(n_480) );
INVx2_ASAP7_75t_L g494 ( .A(n_483), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_484), .A2(n_494), .B(n_508), .C(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g558 ( .A(n_486), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g572 ( .A(n_486), .B(n_501), .Y(n_572) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_487), .B(n_501), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_487), .B(n_575), .Y(n_599) );
OR2x2_ASAP7_75t_L g601 ( .A(n_487), .B(n_559), .Y(n_601) );
AND2x2_ASAP7_75t_L g636 ( .A(n_487), .B(n_559), .Y(n_636) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_487), .Y(n_681) );
INVx1_ASAP7_75t_L g689 ( .A(n_487), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B(n_496), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_498), .A2(n_607), .B1(n_611), .B2(n_615), .C(n_616), .Y(n_606) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g566 ( .A(n_499), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
INVx2_ASAP7_75t_L g565 ( .A(n_500), .Y(n_565) );
AND2x2_ASAP7_75t_L g618 ( .A(n_500), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g637 ( .A(n_500), .B(n_575), .Y(n_637) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g700 ( .A(n_501), .B(n_575), .Y(n_700) );
AND2x2_ASAP7_75t_L g622 ( .A(n_511), .B(n_567), .Y(n_622) );
OAI322xp33_ASAP7_75t_L g690 ( .A1(n_511), .A2(n_646), .A3(n_691), .B1(n_693), .B2(n_696), .C1(n_698), .C2(n_702), .Y(n_690) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_512), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g586 ( .A(n_512), .Y(n_586) );
AND2x2_ASAP7_75t_L g695 ( .A(n_512), .B(n_575), .Y(n_695) );
AND2x2_ASAP7_75t_L g727 ( .A(n_512), .B(n_599), .Y(n_727) );
OR2x2_ASAP7_75t_L g730 ( .A(n_512), .B(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g560 ( .A(n_513), .Y(n_560) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
INVx1_ASAP7_75t_L g743 ( .A(n_520), .Y(n_743) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_538), .Y(n_550) );
INVx2_ASAP7_75t_L g583 ( .A(n_521), .Y(n_583) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g605 ( .A(n_522), .Y(n_605) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
OR2x2_ASAP7_75t_L g737 ( .A(n_522), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g562 ( .A(n_531), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g602 ( .A(n_531), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g654 ( .A(n_531), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_538), .Y(n_531) );
AND2x2_ASAP7_75t_L g551 ( .A(n_532), .B(n_552), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g609 ( .A(n_532), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g663 ( .A(n_532), .B(n_553), .Y(n_663) );
OR2x2_ASAP7_75t_L g671 ( .A(n_532), .B(n_605), .Y(n_671) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g580 ( .A(n_533), .Y(n_580) );
AND2x2_ASAP7_75t_L g590 ( .A(n_533), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g614 ( .A(n_533), .B(n_538), .Y(n_614) );
AND2x2_ASAP7_75t_L g678 ( .A(n_533), .B(n_553), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_538), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_538), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g591 ( .A(n_538), .Y(n_591) );
INVx1_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
AND2x2_ASAP7_75t_L g608 ( .A(n_538), .B(n_609), .Y(n_608) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_538), .Y(n_686) );
INVx1_ASAP7_75t_L g738 ( .A(n_538), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g715 ( .A(n_549), .B(n_624), .Y(n_715) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g642 ( .A(n_551), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g741 ( .A(n_551), .B(n_676), .Y(n_741) );
INVx1_ASAP7_75t_L g563 ( .A(n_552), .Y(n_563) );
AND2x2_ASAP7_75t_L g589 ( .A(n_552), .B(n_583), .Y(n_589) );
BUFx2_ASAP7_75t_L g648 ( .A(n_552), .Y(n_648) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_553), .Y(n_569) );
INVx1_ASAP7_75t_L g579 ( .A(n_553), .Y(n_579) );
NOR2xp67_ASAP7_75t_L g717 ( .A(n_557), .B(n_564), .Y(n_717) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI32xp33_ASAP7_75t_L g561 ( .A1(n_558), .A2(n_562), .A3(n_564), .B1(n_566), .B2(n_568), .Y(n_561) );
AND2x2_ASAP7_75t_L g701 ( .A(n_558), .B(n_574), .Y(n_701) );
AND2x2_ASAP7_75t_L g739 ( .A(n_558), .B(n_637), .Y(n_739) );
INVx1_ASAP7_75t_L g619 ( .A(n_559), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_563), .B(n_625), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_564), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_564), .B(n_567), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_564), .B(n_636), .Y(n_718) );
OR2x2_ASAP7_75t_L g732 ( .A(n_564), .B(n_601), .Y(n_732) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g659 ( .A(n_565), .B(n_567), .Y(n_659) );
OR2x2_ASAP7_75t_L g668 ( .A(n_565), .B(n_655), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_567), .B(n_618), .Y(n_640) );
INVx2_ASAP7_75t_L g655 ( .A(n_569), .Y(n_655) );
OR2x2_ASAP7_75t_L g670 ( .A(n_569), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g685 ( .A(n_569), .B(n_686), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_569), .A2(n_662), .B(n_743), .C(n_744), .Y(n_742) );
OAI321xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_576), .A3(n_581), .B1(n_584), .B2(n_588), .C(n_592), .Y(n_570) );
INVx1_ASAP7_75t_L g683 ( .A(n_571), .Y(n_683) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g694 ( .A(n_572), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g646 ( .A(n_574), .Y(n_646) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_575), .B(n_689), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_576), .A2(n_714), .B1(n_716), .B2(n_718), .C(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
AND2x2_ASAP7_75t_L g651 ( .A(n_578), .B(n_625), .Y(n_651) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_579), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g666 ( .A1(n_581), .A2(n_622), .B(n_667), .C(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g633 ( .A(n_583), .B(n_590), .Y(n_633) );
BUFx2_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
INVx1_ASAP7_75t_L g658 ( .A(n_583), .Y(n_658) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
OR2x2_ASAP7_75t_L g664 ( .A(n_586), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g747 ( .A(n_586), .Y(n_747) );
INVx1_ASAP7_75t_L g740 ( .A(n_587), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g593 ( .A(n_589), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g697 ( .A(n_589), .B(n_614), .Y(n_697) );
INVx1_ASAP7_75t_L g626 ( .A(n_590), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_597), .B1(n_600), .B2(n_602), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_594), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g662 ( .A(n_595), .B(n_663), .Y(n_662) );
BUFx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_596), .B(n_605), .Y(n_625) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g617 ( .A(n_599), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g627 ( .A(n_601), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_604), .A2(n_722), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_721) );
INVx1_ASAP7_75t_L g610 ( .A(n_605), .Y(n_610) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_605), .Y(n_676) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_608), .B(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_609), .A2(n_614), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_612), .B(n_622), .Y(n_719) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g688 ( .A(n_613), .Y(n_688) );
AND2x2_ASAP7_75t_L g647 ( .A(n_614), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g736 ( .A(n_614), .Y(n_736) );
INVx1_ASAP7_75t_L g652 ( .A(n_617), .Y(n_652) );
INVx1_ASAP7_75t_L g707 ( .A(n_618), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B1(n_626), .B2(n_627), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_624), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g692 ( .A(n_625), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_625), .B(n_663), .Y(n_729) );
OR2x2_ASAP7_75t_L g702 ( .A(n_626), .B(n_655), .Y(n_702) );
INVx1_ASAP7_75t_L g641 ( .A(n_627), .Y(n_641) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_629), .B(n_680), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_649), .C(n_660), .Y(n_630) );
OAI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_638), .C(n_644), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_633), .A2(n_704), .B1(n_708), .B2(n_711), .C(n_713), .Y(n_703) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g645 ( .A(n_636), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g699 ( .A(n_636), .B(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_637), .A2(n_685), .B(n_687), .C(n_689), .Y(n_684) );
INVx2_ASAP7_75t_L g731 ( .A(n_637), .Y(n_731) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_641), .B(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g710 ( .A(n_643), .B(n_663), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_652), .B(n_653), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B(n_659), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_654), .B(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_659), .B(n_746), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_666), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g687 ( .A(n_663), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND4x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_703), .C(n_720), .D(n_742), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_690), .Y(n_673) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_679), .B(n_682), .C(n_684), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_678), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_689), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g724 ( .A(n_699), .Y(n_724) );
INVx2_ASAP7_75t_SL g712 ( .A(n_700), .Y(n_712) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g725 ( .A(n_710), .Y(n_725) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_SL g720 ( .A(n_721), .B(n_728), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
OAI221xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_730), .B1(n_732), .B2(n_733), .C(n_734), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g754 ( .A(n_749), .Y(n_754) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
BUFx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
endmodule