module fake_jpeg_14130_n_29 (n_3, n_2, n_1, n_0, n_4, n_5, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_0),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_3),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

O2A1O1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_17),
.B(n_8),
.C(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.C(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_11),
.B(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_3),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_21),
.C(n_19),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_22),
.C(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_17),
.B1(n_12),
.B2(n_18),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

OAI31xp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_0),
.A3(n_2),
.B(n_27),
.Y(n_29)
);


endmodule