module fake_netlist_1_9895_n_21 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
INVx3_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
AOI22xp5_ASAP7_75t_L g12 ( .A1(n_8), .A2(n_0), .B1(n_7), .B2(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx5_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_11), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_14), .Y(n_17) );
OAI221xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_13), .B1(n_12), .B2(n_15), .C(n_2), .Y(n_18) );
O2A1O1Ixp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_15), .B(n_3), .C(n_6), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI22xp5_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_2), .B1(n_10), .B2(n_15), .Y(n_21) );
endmodule