module real_jpeg_23879_n_27 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_156, n_24, n_165, n_6, n_159, n_161, n_162, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_155, n_27);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_156;
input n_24;
input n_165;
input n_6;
input n_159;
input n_161;
input n_162;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_80;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_0),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_1),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_3),
.B(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_56),
.C(n_135),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_7),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_8),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_9),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_10),
.B(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_11),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_138),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_12),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_13),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_14),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_15),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_15),
.B(n_125),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_16),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_16),
.B(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_17),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_17),
.B(n_89),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_19),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_19),
.B(n_58),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_21),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_22),
.B(n_51),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_26),
.B(n_107),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_148),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_42),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_32),
.B(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_35),
.B(n_136),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_36),
.B(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_40),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_40),
.B(n_151),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_41),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_59),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_46),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_147),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_141),
.B(n_146),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_137),
.B(n_140),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_134),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_129),
.B(n_133),
.Y(n_60)
);

OAI321xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_119),
.A3(n_124),
.B1(n_127),
.B2(n_128),
.C(n_155),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_111),
.B(n_118),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_106),
.B(n_110),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_100),
.B(n_105),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B(n_99),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_92),
.B(n_98),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_88),
.B(n_91),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_81),
.B(n_87),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_102),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_145),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_156),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_157),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_158),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_159),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_160),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_161),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_162),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_163),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_164),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_165),
.Y(n_126)
);


endmodule