module fake_jpeg_31697_n_222 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx2_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_40),
.B(n_47),
.Y(n_75)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_25),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_27),
.B2(n_34),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_57),
.B1(n_68),
.B2(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_71),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_34),
.B1(n_21),
.B2(n_25),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_36),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_69),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_18),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_35),
.B(n_29),
.C(n_31),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_21),
.B1(n_35),
.B2(n_22),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_48),
.B1(n_43),
.B2(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_37),
.A2(n_33),
.B1(n_22),
.B2(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_19),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_49),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_85),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_44),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_66),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_50),
.B1(n_42),
.B2(n_48),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_49),
.B(n_16),
.C(n_15),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_98),
.B(n_6),
.C(n_9),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_91),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_45),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_66),
.B1(n_64),
.B2(n_10),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_14),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_0),
.B(n_4),
.C(n_5),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_103),
.B(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_14),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_11),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_60),
.B(n_10),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_64),
.B1(n_65),
.B2(n_63),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_112),
.B1(n_125),
.B2(n_128),
.Y(n_139)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_88),
.B(n_95),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_124),
.B(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_51),
.B1(n_70),
.B2(n_9),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_51),
.B1(n_70),
.B2(n_83),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_77),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_141),
.C(n_85),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_144),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_106),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_148),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_143),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_92),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_84),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_98),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_98),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_154),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_122),
.B1(n_113),
.B2(n_115),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_130),
.B1(n_133),
.B2(n_115),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_122),
.B(n_114),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_159),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_116),
.B1(n_110),
.B2(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_109),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_175),
.B1(n_178),
.B2(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_166),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_161),
.B(n_167),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_164),
.C(n_154),
.Y(n_190)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_132),
.A3(n_139),
.B1(n_141),
.B2(n_137),
.C(n_93),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_129),
.C(n_130),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_183),
.C(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_129),
.C(n_96),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_120),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_179),
.C(n_162),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_189),
.A2(n_195),
.B(n_174),
.C(n_183),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_191),
.B(n_192),
.C(n_193),
.D(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_139),
.B1(n_152),
.B2(n_168),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_200),
.C(n_202),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_165),
.C(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_192),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_159),
.C(n_165),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_156),
.C(n_142),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_186),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_208),
.B(n_207),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_120),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_R g206 ( 
.A(n_196),
.B(n_187),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_117),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_133),
.B1(n_80),
.B2(n_100),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_204),
.B(n_203),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_104),
.C(n_70),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_221),
.Y(n_222)
);


endmodule