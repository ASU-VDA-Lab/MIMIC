module fake_jpeg_18955_n_335 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_13),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_43),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_51),
.Y(n_103)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_14),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_19),
.B1(n_35),
.B2(n_14),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_86),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_59),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_70),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_71),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_82),
.Y(n_116)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_110),
.Y(n_120)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_44),
.B1(n_35),
.B2(n_45),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_106),
.B1(n_98),
.B2(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_41),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_83),
.A2(n_97),
.B1(n_104),
.B2(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_39),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_84),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_29),
.B1(n_19),
.B2(n_48),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_49),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_95),
.B1(n_111),
.B2(n_113),
.Y(n_127)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_89),
.Y(n_121)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_39),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_22),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_93),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_17),
.B(n_1),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_99),
.B(n_0),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_29),
.B1(n_19),
.B2(n_33),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_29),
.B1(n_23),
.B2(n_33),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_101),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_17),
.B(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_17),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_17),
.B1(n_30),
.B2(n_28),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_46),
.B1(n_38),
.B2(n_36),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_32),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_46),
.B1(n_38),
.B2(n_36),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_17),
.B1(n_21),
.B2(n_30),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_32),
.C(n_15),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_118),
.C(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_27),
.C(n_15),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_15),
.B1(n_16),
.B2(n_27),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_136),
.B1(n_138),
.B2(n_152),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_99),
.B(n_95),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_21),
.B(n_30),
.C(n_28),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_95),
.B(n_79),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_18),
.B1(n_27),
.B2(n_16),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_73),
.B1(n_110),
.B2(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_151),
.B1(n_74),
.B2(n_101),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_16),
.C(n_18),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_31),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_111),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_81),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_158),
.Y(n_197)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_173),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_181),
.B(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_160),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_115),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_166),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_88),
.B1(n_96),
.B2(n_75),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_168),
.B1(n_172),
.B2(n_177),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_87),
.B1(n_109),
.B2(n_75),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_127),
.B1(n_149),
.B2(n_135),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_78),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_170),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_77),
.B1(n_90),
.B2(n_72),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_71),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_80),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_80),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_72),
.B1(n_89),
.B2(n_114),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_116),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_31),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_119),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_0),
.B(n_3),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_0),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_148),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_0),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_137),
.B1(n_128),
.B2(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_164),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_200),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_199),
.B(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_118),
.C(n_132),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_196),
.C(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_195),
.B1(n_208),
.B2(n_213),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_124),
.B1(n_147),
.B2(n_130),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_133),
.C(n_146),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_124),
.C(n_138),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_125),
.B1(n_139),
.B2(n_119),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_139),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_205),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_121),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_7),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_125),
.B1(n_121),
.B2(n_122),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_122),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_157),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_5),
.C(n_6),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_7),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_5),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_217),
.A2(n_170),
.B(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_242),
.B1(n_243),
.B2(n_193),
.Y(n_248)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_238),
.C(n_241),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_181),
.B(n_178),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

AO21x1_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_176),
.B(n_174),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_R g245 ( 
.A1(n_228),
.A2(n_186),
.B(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_233),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_183),
.B(n_159),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_231),
.A2(n_234),
.B1(n_244),
.B2(n_199),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_158),
.B(n_154),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_180),
.B(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_175),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_156),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_171),
.B(n_8),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_213),
.C(n_215),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_201),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_248),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_239),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_192),
.C(n_196),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_261),
.C(n_263),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_186),
.B1(n_191),
.B2(n_188),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_255),
.B1(n_258),
.B2(n_260),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_191),
.B1(n_212),
.B2(n_198),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_199),
.B1(n_205),
.B2(n_204),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_202),
.B1(n_211),
.B2(n_9),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_202),
.C(n_9),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_11),
.C(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_233),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_274),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_255),
.C(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_281),
.C(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_279),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_221),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_228),
.B1(n_222),
.B2(n_219),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_248),
.B1(n_251),
.B2(n_259),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_247),
.A2(n_226),
.B(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_257),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_235),
.C(n_236),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_220),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_227),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_266),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_219),
.C(n_220),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_285),
.B1(n_281),
.B2(n_269),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_282),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_295),
.C(n_269),
.Y(n_307)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_229),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

O2A1O1Ixp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_279),
.B(n_262),
.C(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.C(n_310),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_278),
.B1(n_260),
.B2(n_265),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_273),
.C(n_282),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_304),
.A2(n_290),
.B(n_299),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_289),
.C(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_316),
.Y(n_323)
);

XOR2x2_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_286),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_300),
.B(n_303),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_293),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_309),
.B1(n_306),
.B2(n_302),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_241),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_307),
.C(n_292),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_324),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_323),
.C(n_324),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_329),
.B(n_321),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_326),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_327),
.B(n_318),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_320),
.B(n_317),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_316),
.B(n_234),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);


endmodule