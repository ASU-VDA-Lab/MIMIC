module fake_jpeg_24313_n_283 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_25),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_19),
.B1(n_15),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_55),
.B1(n_24),
.B2(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_15),
.B1(n_20),
.B2(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_22),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_22),
.B1(n_24),
.B2(n_32),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_38),
.B1(n_47),
.B2(n_16),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_33),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_35),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_35),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_31),
.B(n_34),
.C(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_33),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_37),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_101),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_61),
.B(n_59),
.C(n_52),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_105),
.B(n_26),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_91),
.B1(n_57),
.B2(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_94),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_54),
.A3(n_37),
.B1(n_72),
.B2(n_79),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_32),
.Y(n_128)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_99),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_40),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_83),
.C(n_64),
.Y(n_116)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_37),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_21),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_34),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_0),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_107),
.B1(n_114),
.B2(n_124),
.Y(n_130)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_47),
.B(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_76),
.B1(n_80),
.B2(n_77),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_120),
.B1(n_122),
.B2(n_86),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_0),
.Y(n_111)
);

NAND2xp67_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_121),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_119),
.C(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_14),
.B(n_17),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_76),
.B1(n_80),
.B2(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_74),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_34),
.A3(n_31),
.B1(n_81),
.B2(n_14),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_16),
.B1(n_25),
.B2(n_54),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_31),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_96),
.C(n_85),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_63),
.C(n_32),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_81),
.Y(n_142)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_137),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_103),
.B1(n_105),
.B2(n_101),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_135),
.B1(n_147),
.B2(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_101),
.B1(n_86),
.B2(n_63),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_140),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_81),
.B1(n_34),
.B2(n_31),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_147),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_145),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_28),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_152),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_98),
.B1(n_94),
.B2(n_32),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_25),
.B1(n_84),
.B2(n_17),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_149),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_90),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_116),
.C(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_172),
.C(n_18),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_163),
.B1(n_137),
.B2(n_131),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_112),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_84),
.B1(n_32),
.B2(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_29),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_140),
.B1(n_139),
.B2(n_134),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_173),
.B1(n_27),
.B2(n_4),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_127),
.B(n_119),
.C(n_106),
.D(n_111),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_114),
.B1(n_127),
.B2(n_118),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_127),
.B(n_124),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_175),
.B(n_177),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_17),
.B(n_26),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_21),
.B(n_28),
.C(n_18),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_153),
.B1(n_152),
.B2(n_145),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_183),
.B1(n_187),
.B2(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_138),
.B1(n_146),
.B2(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_181),
.B(n_164),
.CI(n_156),
.CON(n_212),
.SN(n_212)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_90),
.B1(n_67),
.B2(n_62),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_90),
.C(n_67),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_194),
.C(n_198),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_62),
.B1(n_29),
.B2(n_27),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_0),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_29),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_168),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_29),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_174),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_29),
.C(n_27),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_195),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_27),
.C(n_2),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_159),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_167),
.C(n_172),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_209),
.C(n_213),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_206),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_171),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_210),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_164),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_192),
.B1(n_189),
.B2(n_182),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_156),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_216),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_201),
.C(n_200),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_215),
.B(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_177),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_231),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_227),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_186),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_228),
.B(n_229),
.CI(n_13),
.CON(n_243),
.SN(n_243)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_183),
.B1(n_196),
.B2(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_168),
.B1(n_189),
.B2(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_1),
.C(n_4),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_217),
.C(n_209),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_228),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_226),
.B1(n_240),
.B2(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_1),
.C(n_4),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_4),
.C(n_5),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_5),
.C(n_6),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_10),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_234),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_245),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_13),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_222),
.B1(n_229),
.B2(n_224),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_253),
.C(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_256),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_219),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_10),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_10),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_5),
.Y(n_257)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_11),
.B(n_13),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_262),
.A2(n_263),
.B(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_11),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_11),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_250),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_272),
.B(n_6),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_12),
.C(n_7),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_258),
.B(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_274),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_6),
.B(n_7),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_276),
.B(n_268),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_267),
.B(n_277),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_7),
.C(n_8),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_8),
.B(n_264),
.Y(n_283)
);


endmodule