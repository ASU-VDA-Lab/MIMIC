module fake_jpeg_31845_n_537 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_537);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx2_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2x1_ASAP7_75t_SL g135 ( 
.A(n_57),
.B(n_79),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_61),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_20),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_74),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_86),
.Y(n_131)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_28),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_91),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_1),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_16),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_105),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_34),
.Y(n_143)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_46),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_102),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_37),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_49),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_39),
.B(n_15),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_106),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_30),
.B(n_26),
.C(n_43),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_109),
.B(n_141),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_57),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_120),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_125),
.A2(n_95),
.B1(n_49),
.B2(n_35),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

BUFx4f_ASAP7_75t_SL g132 ( 
.A(n_53),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_132),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_91),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_140),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_97),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_30),
.B(n_26),
.C(n_43),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_164),
.Y(n_173)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_151),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_168),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_80),
.A2(n_87),
.B1(n_99),
.B2(n_101),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_103),
.B1(n_71),
.B2(n_92),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_82),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_72),
.B(n_52),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_45),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_94),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_169),
.B(n_156),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_50),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_171),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_174),
.A2(n_175),
.B1(n_186),
.B2(n_198),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_109),
.A2(n_90),
.B1(n_81),
.B2(n_77),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_179),
.A2(n_202),
.B1(n_167),
.B2(n_145),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

BUFx2_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_70),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_183),
.B(n_177),
.Y(n_264)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_135),
.A2(n_73),
.B1(n_85),
.B2(n_78),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_59),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_188),
.B(n_189),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_124),
.B(n_55),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g271 ( 
.A(n_190),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_139),
.B(n_52),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_199),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_194),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_197),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_35),
.B1(n_32),
.B2(n_47),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_111),
.B(n_45),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_50),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_216),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_107),
.A2(n_67),
.B1(n_63),
.B2(n_58),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_48),
.B1(n_47),
.B2(n_37),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_158),
.B1(n_154),
.B2(n_128),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_209),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_115),
.B(n_37),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_212),
.C(n_129),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_37),
.C(n_106),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_40),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_157),
.A2(n_48),
.B1(n_35),
.B2(n_32),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_125),
.B1(n_165),
.B2(n_155),
.Y(n_232)
);

CKINVDCx12_ASAP7_75t_R g220 ( 
.A(n_151),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_126),
.B(n_40),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_226),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_147),
.B(n_14),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_121),
.B(n_14),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_228),
.A2(n_255),
.B1(n_267),
.B2(n_175),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_232),
.A2(n_202),
.B1(n_214),
.B2(n_133),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_170),
.A2(n_167),
.B1(n_155),
.B2(n_154),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_236),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_243),
.A2(n_272),
.B(n_224),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_158),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_256),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_181),
.A2(n_163),
.B1(n_162),
.B2(n_128),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_173),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_171),
.B(n_121),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_257),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_191),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_136),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_213),
.A2(n_174),
.B1(n_186),
.B2(n_222),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_183),
.A2(n_113),
.B1(n_149),
.B2(n_127),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_187),
.A2(n_113),
.B(n_133),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_127),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

INVx4_ASAP7_75t_SL g311 ( 
.A(n_274),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_198),
.B(n_225),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_310),
.B1(n_254),
.B2(n_232),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_212),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_276),
.B(n_280),
.Y(n_337)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_250),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_182),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_284),
.A2(n_229),
.B1(n_246),
.B2(n_271),
.Y(n_324)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_286),
.A2(n_232),
.B1(n_228),
.B2(n_255),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_200),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_196),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_296),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_194),
.C(n_221),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_303),
.C(n_267),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_191),
.C(n_205),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_299),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_205),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_291),
.B(n_292),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_295),
.B(n_301),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_236),
.B(n_197),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_302),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_233),
.B(n_149),
.C(n_219),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_244),
.B(n_214),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_236),
.B(n_258),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_307),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_156),
.Y(n_307)
);

AOI22x1_ASAP7_75t_SL g308 ( 
.A1(n_233),
.A2(n_224),
.B1(n_132),
.B2(n_210),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_308),
.A2(n_246),
.B(n_274),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_210),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_232),
.A2(n_204),
.B1(n_209),
.B2(n_193),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_313),
.A2(n_314),
.B1(n_271),
.B2(n_311),
.Y(n_320)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_263),
.B(n_225),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_315),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_316),
.A2(n_325),
.B1(n_341),
.B2(n_350),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_320),
.A2(n_330),
.B(n_351),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_321),
.A2(n_324),
.B1(n_339),
.B2(n_129),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_299),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_310),
.B1(n_279),
.B2(n_277),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_326),
.A2(n_344),
.B(n_346),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_242),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_313),
.C(n_300),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_302),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_329),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_249),
.B1(n_230),
.B2(n_259),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_247),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_290),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_284),
.A2(n_190),
.B1(n_195),
.B2(n_206),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_279),
.A2(n_265),
.B1(n_268),
.B2(n_237),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_277),
.A2(n_268),
.B1(n_237),
.B2(n_231),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_311),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_306),
.A2(n_234),
.B(n_230),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_234),
.B(n_253),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_291),
.A2(n_231),
.B1(n_165),
.B2(n_253),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_351),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_307),
.A2(n_248),
.B1(n_207),
.B2(n_251),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_348),
.B(n_281),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_353),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_332),
.B(n_287),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_356),
.B(n_366),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_298),
.Y(n_357)
);

NOR4xp25_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_360),
.C(n_362),
.D(n_361),
.Y(n_398)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_292),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_289),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_368),
.C(n_373),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_334),
.B(n_309),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_324),
.A2(n_339),
.B1(n_316),
.B2(n_347),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_369),
.A2(n_328),
.B(n_338),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_303),
.Y(n_370)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_336),
.Y(n_371)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_297),
.B1(n_314),
.B2(n_294),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_372),
.A2(n_375),
.B1(n_329),
.B2(n_322),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_285),
.C(n_312),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_374),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_325),
.A2(n_278),
.B1(n_283),
.B2(n_293),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_381),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

OAI21xp33_ASAP7_75t_SL g391 ( 
.A1(n_378),
.A2(n_358),
.B(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_224),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_380),
.A2(n_323),
.B(n_326),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_319),
.A2(n_42),
.B1(n_123),
.B2(n_32),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_386),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_333),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_383),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_344),
.B(n_14),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_384),
.Y(n_389)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_388),
.A2(n_390),
.B(n_391),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_350),
.B(n_341),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_392),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_370),
.B(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_393),
.B(n_398),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_327),
.B1(n_352),
.B2(n_335),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_395),
.A2(n_401),
.B1(n_383),
.B2(n_355),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_363),
.A2(n_338),
.B(n_352),
.Y(n_402)
);

AO22x1_ASAP7_75t_L g436 ( 
.A1(n_402),
.A2(n_385),
.B1(n_379),
.B2(n_374),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_409),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_363),
.A2(n_327),
.B(n_345),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_403),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_365),
.A2(n_322),
.B1(n_345),
.B2(n_42),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_375),
.A2(n_136),
.B1(n_123),
.B2(n_12),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_355),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_419),
.A2(n_435),
.B1(n_436),
.B2(n_415),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_420),
.A2(n_443),
.B1(n_417),
.B2(n_405),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_364),
.C(n_376),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_425),
.C(n_404),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_368),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_430),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_373),
.C(n_371),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_353),
.Y(n_427)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_427),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_382),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_437),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_386),
.Y(n_429)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_393),
.B(n_408),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_396),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_434),
.B(n_438),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_395),
.A2(n_381),
.B1(n_378),
.B2(n_380),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_2),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_439),
.B(n_441),
.Y(n_452)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

AO22x1_ASAP7_75t_SL g442 ( 
.A1(n_394),
.A2(n_414),
.B1(n_400),
.B2(n_402),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_442),
.B(n_444),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_29),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_394),
.B(n_2),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_427),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_447),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_428),
.A2(n_405),
.B1(n_404),
.B2(n_390),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_448),
.A2(n_454),
.B1(n_456),
.B2(n_460),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_389),
.B1(n_409),
.B2(n_406),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_461),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_421),
.Y(n_470)
);

OAI22x1_ASAP7_75t_L g454 ( 
.A1(n_436),
.A2(n_402),
.B1(n_407),
.B2(n_413),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_425),
.B(n_416),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_443),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_413),
.B1(n_415),
.B2(n_416),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_465),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_422),
.A2(n_411),
.B1(n_397),
.B2(n_12),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_435),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_29),
.Y(n_465)
);

INVx11_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_479),
.Y(n_497)
);

INVx13_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_480),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_478),
.C(n_482),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_466),
.A2(n_419),
.B1(n_418),
.B2(n_420),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_464),
.B1(n_465),
.B2(n_462),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_446),
.A2(n_436),
.B(n_418),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_460),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_459),
.A2(n_456),
.B(n_448),
.Y(n_476)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_476),
.Y(n_494)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_430),
.C(n_437),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_451),
.B(n_442),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_458),
.B(n_442),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_439),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_429),
.C(n_423),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_485),
.B(n_486),
.Y(n_511)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_469),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_489),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_452),
.B1(n_450),
.B2(n_444),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_482),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_493),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_464),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_495),
.B(n_472),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_476),
.A2(n_471),
.B(n_481),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_499),
.Y(n_507)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_470),
.C(n_490),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_504),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_484),
.A2(n_467),
.B1(n_480),
.B2(n_483),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_492),
.A2(n_467),
.B(n_477),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_509),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_472),
.C(n_457),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_508),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_494),
.A2(n_479),
.B1(n_473),
.B2(n_431),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_475),
.C(n_469),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_475),
.C(n_29),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_475),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_501),
.A2(n_488),
.B1(n_498),
.B2(n_4),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_519),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_511),
.Y(n_519)
);

AOI31xp67_ASAP7_75t_L g521 ( 
.A1(n_502),
.A2(n_2),
.A3(n_3),
.B(n_5),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_507),
.C(n_510),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_525),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_503),
.C(n_506),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_523),
.B(n_524),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_509),
.C(n_6),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_5),
.C(n_6),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_5),
.C(n_10),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_516),
.B(n_519),
.Y(n_528)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_528),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_527),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_531),
.B(n_529),
.Y(n_533)
);

INVxp33_ASAP7_75t_L g534 ( 
.A(n_533),
.Y(n_534)
);

AOI322xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_5),
.A3(n_10),
.B1(n_11),
.B2(n_520),
.C1(n_532),
.C2(n_533),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_10),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_11),
.Y(n_537)
);


endmodule