module fake_netlist_6_148_n_1031 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1031);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1031;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_608;
wire n_261;
wire n_474;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_964;
wire n_802;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_267;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_37),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_9),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_216),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_178),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_119),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_126),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_180),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_102),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_195),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_9),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_12),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_37),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_123),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_122),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_114),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_108),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_170),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_116),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_90),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_152),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_192),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_124),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_87),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_117),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_32),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_13),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_155),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_147),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_199),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

HB1xp67_ASAP7_75t_SL g276 ( 
.A(n_157),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_187),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_68),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_109),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_112),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_105),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_135),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_31),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_42),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_46),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_38),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_72),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_36),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_164),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_98),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_113),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_104),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_83),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_137),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_226),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_145),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_140),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_33),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_121),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_130),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_221),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_85),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_88),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_210),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_156),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_131),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_94),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_7),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_215),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_111),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_163),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_166),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_107),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_21),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_133),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_158),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_151),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_40),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_211),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_22),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_63),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_230),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_243),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_228),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_244),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_233),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_235),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_284),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_236),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_234),
.B(n_0),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_0),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_238),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_247),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

INVx4_ASAP7_75t_R g346 ( 
.A(n_276),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_244),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_253),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_259),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_255),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_255),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_237),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_239),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_261),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_234),
.B(n_1),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_284),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_240),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_256),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_229),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_270),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_241),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_275),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_232),
.B(n_1),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_231),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_242),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_293),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_249),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_273),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_273),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_250),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_252),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_280),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_254),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_309),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_280),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_350),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_328),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_232),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_335),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_372),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_277),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_360),
.B(n_257),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_352),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_314),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_353),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_359),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_363),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_374),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_325),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g420 ( 
.A1(n_339),
.A2(n_282),
.B(n_277),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

AND2x4_ASAP7_75t_SL g422 ( 
.A(n_333),
.B(n_286),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_361),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_282),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_374),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_347),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_351),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_365),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_371),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_357),
.B(n_321),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_293),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_398),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_262),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_405),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_390),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_297),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_397),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_246),
.B1(n_248),
.B2(n_245),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_409),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_285),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_435),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_346),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_290),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_385),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_302),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_402),
.B(n_303),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_386),
.B(n_293),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_387),
.B(n_295),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_381),
.B(n_286),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_396),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_392),
.B(n_258),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_386),
.B(n_295),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_419),
.B(n_268),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_381),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_433),
.B(n_413),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_422),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_420),
.B(n_295),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_420),
.B(n_260),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_421),
.B(n_299),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_394),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_425),
.B(n_299),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_401),
.B(n_295),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_432),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_401),
.B(n_287),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_403),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_404),
.A2(n_289),
.B1(n_300),
.B2(n_316),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_422),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_425),
.B(n_377),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_445),
.B(n_423),
.Y(n_514)
);

AND2x6_ASAP7_75t_SL g515 ( 
.A(n_512),
.B(n_326),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_496),
.A2(n_305),
.B1(n_265),
.B2(n_311),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_463),
.A2(n_377),
.B1(n_380),
.B2(n_423),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_445),
.A2(n_418),
.B1(n_267),
.B2(n_312),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_269),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_439),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_440),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_448),
.B(n_271),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_446),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_461),
.B(n_272),
.Y(n_527)
);

O2A1O1Ixp5_ASAP7_75t_L g528 ( 
.A1(n_494),
.A2(n_305),
.B(n_323),
.C(n_319),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_457),
.A2(n_380),
.B1(n_326),
.B2(n_358),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_461),
.B(n_274),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_443),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_454),
.B(n_279),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_498),
.A2(n_313),
.B1(n_283),
.B2(n_288),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_SL g535 ( 
.A(n_459),
.B(n_429),
.C(n_291),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_451),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_511),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_443),
.B(n_281),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_476),
.A2(n_331),
.B1(n_336),
.B2(n_358),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_441),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_484),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_462),
.B(n_292),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_466),
.B(n_449),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_464),
.B(n_305),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_480),
.B(n_429),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_496),
.A2(n_305),
.B1(n_294),
.B2(n_315),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_480),
.B(n_331),
.Y(n_552)
);

A2O1A1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_469),
.A2(n_450),
.B(n_458),
.C(n_452),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_469),
.A2(n_318),
.B(n_304),
.C(n_306),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_487),
.A2(n_296),
.B1(n_307),
.B2(n_317),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_467),
.A2(n_336),
.B1(n_417),
.B2(n_408),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_475),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_470),
.B(n_428),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_493),
.B(n_43),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_493),
.B(n_44),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_504),
.B(n_428),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_455),
.B(n_45),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_504),
.B(n_397),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_493),
.A2(n_417),
.B1(n_408),
.B2(n_4),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_493),
.B(n_47),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_492),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_472),
.B(n_2),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_497),
.A2(n_100),
.B1(n_224),
.B2(n_223),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_472),
.B(n_2),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_493),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_493),
.B(n_48),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_444),
.B(n_49),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

NOR2x1p5_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_3),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_L g579 ( 
.A(n_444),
.B(n_50),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_444),
.B(n_51),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_468),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_484),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_482),
.B(n_52),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_486),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_486),
.Y(n_585)
);

AO221x1_ASAP7_75t_L g586 ( 
.A1(n_507),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_444),
.B(n_53),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_485),
.B(n_6),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_482),
.B(n_54),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_477),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_502),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_444),
.B(n_55),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_502),
.B(n_56),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_481),
.A2(n_125),
.B(n_222),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_444),
.B(n_57),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_453),
.A2(n_127),
.B(n_220),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_488),
.B(n_58),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_499),
.A2(n_120),
.B1(n_219),
.B2(n_218),
.Y(n_599)
);

NAND2x1p5_ASAP7_75t_L g600 ( 
.A(n_532),
.B(n_513),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_564),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_568),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_552),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_SL g604 ( 
.A(n_517),
.B(n_485),
.C(n_503),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_545),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_518),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_522),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_548),
.B(n_483),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_544),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_SL g610 ( 
.A(n_517),
.B(n_557),
.C(n_529),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_584),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_550),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_514),
.B(n_532),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_544),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_540),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_519),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_556),
.B(n_533),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

NOR2x1_ASAP7_75t_R g619 ( 
.A(n_537),
.B(n_511),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_582),
.B(n_509),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_533),
.B(n_483),
.Y(n_621)
);

BUFx5_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_577),
.B(n_509),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_545),
.B(n_508),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_546),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_SL g627 ( 
.A(n_559),
.B(n_505),
.C(n_501),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_545),
.B(n_508),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_545),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_540),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx3_ASAP7_75t_SL g632 ( 
.A(n_559),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_569),
.B(n_483),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_553),
.B(n_511),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_585),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_563),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_547),
.B(n_525),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_526),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_566),
.B(n_506),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_578),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_576),
.B(n_513),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_596),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_521),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_588),
.B(n_510),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_569),
.B(n_479),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_515),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_536),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_538),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_SL g650 ( 
.A(n_562),
.B(n_457),
.C(n_500),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_447),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_539),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_541),
.Y(n_654)
);

NOR2x1p5_ASAP7_75t_L g655 ( 
.A(n_527),
.B(n_491),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_581),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_566),
.B(n_475),
.C(n_489),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_535),
.Y(n_658)
);

NOR2x1_ASAP7_75t_L g659 ( 
.A(n_583),
.B(n_447),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_R g660 ( 
.A(n_525),
.B(n_447),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_565),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_590),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_516),
.B(n_460),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_460),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_575),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_531),
.Y(n_666)
);

NOR2x1_ASAP7_75t_L g667 ( 
.A(n_629),
.B(n_562),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_617),
.A2(n_551),
.B1(n_572),
.B2(n_520),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_621),
.A2(n_561),
.B(n_560),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_659),
.A2(n_528),
.B(n_567),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_605),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_549),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_606),
.Y(n_673)
);

NAND2x1_ASAP7_75t_L g674 ( 
.A(n_638),
.B(n_489),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_620),
.B(n_609),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_621),
.A2(n_574),
.B(n_558),
.Y(n_676)
);

NAND4xp25_ASAP7_75t_L g677 ( 
.A(n_623),
.B(n_542),
.C(n_572),
.D(n_555),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_652),
.A2(n_554),
.B(n_549),
.Y(n_678)
);

AO31x2_ASAP7_75t_L g679 ( 
.A1(n_633),
.A2(n_591),
.A3(n_570),
.B(n_594),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_612),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_657),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_637),
.B(n_571),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_608),
.A2(n_579),
.B(n_489),
.Y(n_683)
);

AO31x2_ASAP7_75t_L g684 ( 
.A1(n_633),
.A2(n_597),
.A3(n_592),
.B(n_587),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_625),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_666),
.B(n_534),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_608),
.A2(n_589),
.B(n_583),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_605),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_616),
.Y(n_689)
);

CKINVDCx11_ASAP7_75t_R g690 ( 
.A(n_646),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_643),
.B(n_535),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_613),
.A2(n_593),
.B(n_589),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_622),
.B(n_593),
.Y(n_693)
);

BUFx2_ASAP7_75t_SL g694 ( 
.A(n_618),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_614),
.B(n_586),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_654),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_622),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_610),
.B(n_599),
.C(n_598),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_652),
.A2(n_598),
.B(n_595),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_632),
.B(n_603),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_622),
.B(n_580),
.Y(n_701)
);

CKINVDCx12_ASAP7_75t_R g702 ( 
.A(n_619),
.Y(n_702)
);

AOI21x1_ASAP7_75t_L g703 ( 
.A1(n_645),
.A2(n_460),
.B(n_475),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_SL g704 ( 
.A1(n_636),
.A2(n_475),
.B(n_474),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_605),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_639),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_644),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_663),
.A2(n_474),
.B(n_456),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_605),
.A2(n_474),
.B(n_456),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_607),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_618),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_643),
.B(n_456),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_622),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_624),
.B(n_456),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_615),
.B(n_59),
.Y(n_715)
);

OAI21x1_ASAP7_75t_SL g716 ( 
.A1(n_663),
.A2(n_132),
.B(n_225),
.Y(n_716)
);

OAI21x1_ASAP7_75t_L g717 ( 
.A1(n_664),
.A2(n_474),
.B(n_473),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_664),
.A2(n_473),
.B(n_128),
.Y(n_718)
);

AOI211x1_ASAP7_75t_L g719 ( 
.A1(n_626),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_630),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_631),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_697),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_691),
.B(n_644),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_668),
.A2(n_657),
.B1(n_651),
.B2(n_600),
.Y(n_725)
);

AO31x2_ASAP7_75t_L g726 ( 
.A1(n_706),
.A2(n_645),
.A3(n_602),
.B(n_601),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_710),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_720),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_680),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_689),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_720),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_697),
.Y(n_733)
);

AOI221xp5_ASAP7_75t_L g734 ( 
.A1(n_677),
.A2(n_604),
.B1(n_706),
.B2(n_698),
.C(n_707),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_671),
.Y(n_735)
);

AO31x2_ASAP7_75t_L g736 ( 
.A1(n_669),
.A2(n_648),
.A3(n_647),
.B(n_653),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_695),
.A2(n_658),
.B1(n_661),
.B2(n_641),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_667),
.B(n_625),
.Y(n_738)
);

OAI222xp33_ASAP7_75t_L g739 ( 
.A1(n_682),
.A2(n_640),
.B1(n_642),
.B2(n_600),
.C1(n_634),
.C2(n_662),
.Y(n_739)
);

AOI21x1_ASAP7_75t_L g740 ( 
.A1(n_703),
.A2(n_634),
.B(n_656),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_689),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_681),
.B(n_650),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_696),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_687),
.A2(n_662),
.A3(n_622),
.B(n_627),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_708),
.A2(n_638),
.B(n_649),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_696),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_708),
.A2(n_649),
.B(n_635),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_686),
.A2(n_651),
.B1(n_636),
.B2(n_641),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_713),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_690),
.Y(n_750)
);

OAI22x1_ASAP7_75t_L g751 ( 
.A1(n_681),
.A2(n_655),
.B1(n_628),
.B2(n_611),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_717),
.A2(n_635),
.B(n_611),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_675),
.A2(n_628),
.B1(n_636),
.B2(n_646),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_672),
.B(n_660),
.Y(n_754)
);

NOR2x1_ASAP7_75t_R g755 ( 
.A(n_690),
.B(n_694),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_707),
.A2(n_665),
.B(n_18),
.C(n_19),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_713),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_700),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_712),
.B(n_711),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_671),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_692),
.B(n_665),
.Y(n_761)
);

AOI21x1_ASAP7_75t_L g762 ( 
.A1(n_676),
.A2(n_665),
.B(n_473),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_685),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_714),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_688),
.B(n_61),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_685),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_678),
.B(n_17),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_685),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_693),
.A2(n_473),
.B1(n_18),
.B2(n_19),
.Y(n_769)
);

NOR2x1_ASAP7_75t_SL g770 ( 
.A(n_693),
.B(n_64),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_688),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_702),
.B(n_17),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_679),
.B(n_20),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_732),
.Y(n_774)
);

NAND2x1_ASAP7_75t_L g775 ( 
.A(n_735),
.B(n_704),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_723),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_722),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_724),
.B(n_715),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_727),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_728),
.B(n_705),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_730),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_728),
.B(n_768),
.Y(n_782)
);

INVx3_ASAP7_75t_SL g783 ( 
.A(n_750),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_759),
.B(n_719),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_768),
.B(n_705),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_722),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_767),
.A2(n_718),
.B1(n_683),
.B2(n_701),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_749),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_734),
.A2(n_716),
.B1(n_701),
.B2(n_674),
.C(n_679),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_731),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_758),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_767),
.A2(n_699),
.B1(n_670),
.B2(n_679),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_742),
.A2(n_670),
.B1(n_679),
.B2(n_473),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_741),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_749),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_742),
.B(n_20),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_SL g797 ( 
.A1(n_754),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_773),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_737),
.B(n_684),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_729),
.B(n_684),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_771),
.Y(n_801)
);

BUFx8_ASAP7_75t_L g802 ( 
.A(n_766),
.Y(n_802)
);

OAI211xp5_ASAP7_75t_L g803 ( 
.A1(n_756),
.A2(n_709),
.B(n_26),
.C(n_27),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_762),
.A2(n_684),
.B(n_473),
.Y(n_804)
);

AOI221xp5_ASAP7_75t_SL g805 ( 
.A1(n_756),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.C(n_29),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_771),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_739),
.B(n_28),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_SL g808 ( 
.A1(n_725),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_769),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_753),
.B(n_35),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_743),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_751),
.B(n_684),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_761),
.A2(n_35),
.B(n_36),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_748),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_751),
.B(n_65),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_773),
.A2(n_39),
.B1(n_41),
.B2(n_66),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_757),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_764),
.B(n_41),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_757),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_735),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_733),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_750),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_738),
.A2(n_217),
.B1(n_69),
.B2(n_71),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_763),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_738),
.B(n_67),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_765),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_733),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_738),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_761),
.A2(n_77),
.B(n_78),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_812),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_787),
.A2(n_740),
.B(n_745),
.Y(n_832)
);

AOI221xp5_ASAP7_75t_L g833 ( 
.A1(n_798),
.A2(n_772),
.B1(n_765),
.B2(n_763),
.C(n_760),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_808),
.A2(n_807),
.B1(n_809),
.B2(n_816),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_808),
.A2(n_765),
.B1(n_760),
.B2(n_735),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_823),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_798),
.A2(n_733),
.B1(n_726),
.B2(n_770),
.C(n_755),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_807),
.A2(n_752),
.B(n_747),
.C(n_745),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_783),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_812),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_827),
.A2(n_726),
.B(n_744),
.C(n_736),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_777),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_800),
.B(n_726),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_812),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_791),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_799),
.B(n_726),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_809),
.A2(n_752),
.B1(n_747),
.B2(n_744),
.Y(n_847)
);

OR2x2_ASAP7_75t_SL g848 ( 
.A(n_784),
.B(n_726),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_822),
.B(n_736),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_816),
.A2(n_744),
.B1(n_736),
.B2(n_82),
.Y(n_850)
);

OAI211xp5_ASAP7_75t_L g851 ( 
.A1(n_813),
.A2(n_744),
.B(n_736),
.C(n_84),
.Y(n_851)
);

INVx5_ASAP7_75t_SL g852 ( 
.A(n_815),
.Y(n_852)
);

AOI221xp5_ASAP7_75t_L g853 ( 
.A1(n_797),
.A2(n_736),
.B1(n_744),
.B2(n_86),
.C(n_89),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_791),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_778),
.A2(n_796),
.B1(n_824),
.B2(n_815),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_822),
.B(n_80),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_814),
.A2(n_81),
.B1(n_91),
.B2(n_92),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_824),
.A2(n_93),
.B1(n_99),
.B2(n_101),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_774),
.Y(n_859)
);

OA21x2_ASAP7_75t_L g860 ( 
.A1(n_793),
.A2(n_792),
.B(n_804),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_790),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_794),
.B(n_214),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_777),
.Y(n_863)
);

AOI221xp5_ASAP7_75t_L g864 ( 
.A1(n_805),
.A2(n_103),
.B1(n_106),
.B2(n_110),
.C(n_115),
.Y(n_864)
);

AND2x4_ASAP7_75t_SL g865 ( 
.A(n_815),
.B(n_118),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_818),
.A2(n_129),
.B1(n_134),
.B2(n_136),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_786),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_792),
.A2(n_138),
.B(n_139),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_786),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_810),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_803),
.A2(n_148),
.B1(n_150),
.B2(n_153),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_811),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_819),
.B(n_781),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_829),
.B(n_793),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_842),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_861),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_861),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_872),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_846),
.B(n_776),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_846),
.B(n_779),
.Y(n_880)
);

OAI21xp33_ASAP7_75t_L g881 ( 
.A1(n_834),
.A2(n_827),
.B(n_830),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_843),
.B(n_828),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_843),
.B(n_828),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_848),
.B(n_787),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_873),
.B(n_820),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_855),
.A2(n_826),
.B(n_789),
.Y(n_886)
);

NAND2x1_ASAP7_75t_L g887 ( 
.A(n_831),
.B(n_821),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_831),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_849),
.B(n_788),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_872),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_863),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_849),
.B(n_788),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_863),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_840),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_840),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_863),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_867),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_844),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_844),
.B(n_795),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_873),
.B(n_817),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_867),
.B(n_782),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_867),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_845),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_836),
.B(n_859),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_869),
.Y(n_905)
);

AND2x4_ASAP7_75t_SL g906 ( 
.A(n_854),
.B(n_782),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_876),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_906),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_881),
.A2(n_852),
.B1(n_858),
.B2(n_871),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_903),
.B(n_852),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_876),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_877),
.Y(n_912)
);

OAI221xp5_ASAP7_75t_L g913 ( 
.A1(n_881),
.A2(n_833),
.B1(n_870),
.B2(n_864),
.C(n_853),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_879),
.B(n_860),
.Y(n_914)
);

OAI221xp5_ASAP7_75t_L g915 ( 
.A1(n_886),
.A2(n_857),
.B1(n_837),
.B2(n_850),
.C(n_866),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_886),
.A2(n_852),
.B1(n_865),
.B2(n_835),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_879),
.B(n_852),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_875),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_904),
.B(n_839),
.Y(n_919)
);

AOI222xp33_ASAP7_75t_L g920 ( 
.A1(n_880),
.A2(n_865),
.B1(n_852),
.B2(n_851),
.C1(n_862),
.C2(n_783),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_L g921 ( 
.A1(n_884),
.A2(n_874),
.B1(n_839),
.B2(n_865),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_906),
.Y(n_922)
);

NAND3xp33_ASAP7_75t_SL g923 ( 
.A(n_884),
.B(n_806),
.C(n_862),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_901),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_877),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_880),
.B(n_848),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_926),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_910),
.B(n_917),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_907),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_914),
.B(n_894),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_914),
.B(n_894),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_918),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_924),
.B(n_895),
.Y(n_933)
);

NOR4xp25_ASAP7_75t_SL g934 ( 
.A(n_915),
.B(n_895),
.C(n_841),
.D(n_878),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_918),
.B(n_888),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_922),
.B(n_825),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_911),
.B(n_901),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_919),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_912),
.B(n_882),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_925),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_923),
.B(n_882),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_929),
.B(n_878),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_L g943 ( 
.A(n_941),
.B(n_908),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_927),
.B(n_908),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_933),
.B(n_883),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_937),
.B(n_889),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_928),
.A2(n_909),
.B1(n_913),
.B2(n_916),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_930),
.B(n_898),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_929),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_947),
.B(n_930),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_943),
.A2(n_920),
.B1(n_921),
.B2(n_936),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_949),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_942),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_944),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_948),
.B(n_931),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_948),
.B(n_931),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_952),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_951),
.A2(n_934),
.B1(n_950),
.B2(n_954),
.Y(n_958)
);

AOI222xp33_ASAP7_75t_L g959 ( 
.A1(n_954),
.A2(n_938),
.B1(n_921),
.B2(n_933),
.C1(n_942),
.C2(n_940),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_953),
.B(n_946),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_957),
.B(n_955),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_960),
.Y(n_962)
);

AOI211xp5_ASAP7_75t_L g963 ( 
.A1(n_958),
.A2(n_919),
.B(n_953),
.C(n_955),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_959),
.Y(n_964)
);

OAI321xp33_ASAP7_75t_L g965 ( 
.A1(n_963),
.A2(n_964),
.A3(n_962),
.B1(n_961),
.B2(n_956),
.C(n_934),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_964),
.B(n_956),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_962),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_964),
.B(n_802),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_962),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_966),
.A2(n_939),
.B1(n_940),
.B2(n_945),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_SL g971 ( 
.A1(n_967),
.A2(n_935),
.B(n_932),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_935),
.Y(n_972)
);

AOI211xp5_ASAP7_75t_L g973 ( 
.A1(n_965),
.A2(n_868),
.B(n_856),
.C(n_780),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_969),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_966),
.B(n_932),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_967),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_968),
.B(n_802),
.C(n_801),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_973),
.A2(n_976),
.B1(n_974),
.B2(n_975),
.C(n_972),
.Y(n_978)
);

OAI211xp5_ASAP7_75t_L g979 ( 
.A1(n_977),
.A2(n_887),
.B(n_868),
.C(n_856),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_SL g980 ( 
.A(n_970),
.B(n_887),
.Y(n_980)
);

XNOR2x2_ASAP7_75t_L g981 ( 
.A(n_971),
.B(n_885),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_972),
.A2(n_906),
.B(n_898),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_L g983 ( 
.A1(n_972),
.A2(n_898),
.B(n_900),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_SL g984 ( 
.A1(n_973),
.A2(n_838),
.B(n_847),
.C(n_874),
.Y(n_984)
);

AOI211xp5_ASAP7_75t_L g985 ( 
.A1(n_973),
.A2(n_780),
.B(n_801),
.C(n_785),
.Y(n_985)
);

AOI31xp33_ASAP7_75t_L g986 ( 
.A1(n_978),
.A2(n_785),
.A3(n_900),
.B(n_890),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_SL g987 ( 
.A(n_985),
.B(n_979),
.C(n_982),
.Y(n_987)
);

NOR2x1_ASAP7_75t_R g988 ( 
.A(n_981),
.B(n_801),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_888),
.Y(n_990)
);

AOI221x1_ASAP7_75t_L g991 ( 
.A1(n_984),
.A2(n_801),
.B1(n_890),
.B2(n_888),
.C(n_821),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_981),
.B(n_899),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_978),
.A2(n_775),
.B(n_899),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_980),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_986),
.B(n_905),
.C(n_891),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_994),
.B(n_883),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_987),
.B(n_154),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_SL g998 ( 
.A1(n_989),
.A2(n_992),
.B(n_990),
.Y(n_998)
);

AND2x2_ASAP7_75t_SL g999 ( 
.A(n_988),
.B(n_888),
.Y(n_999)
);

AND3x2_ASAP7_75t_L g1000 ( 
.A(n_991),
.B(n_159),
.C(n_160),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_905),
.C(n_891),
.Y(n_1001)
);

NAND3x2_ASAP7_75t_L g1002 ( 
.A(n_994),
.B(n_892),
.C(n_889),
.Y(n_1002)
);

OAI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_986),
.A2(n_888),
.B1(n_897),
.B2(n_902),
.C(n_896),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_996),
.A2(n_888),
.B1(n_892),
.B2(n_897),
.Y(n_1004)
);

NAND5xp2_ASAP7_75t_L g1005 ( 
.A(n_1001),
.B(n_161),
.C(n_162),
.D(n_165),
.E(n_167),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_998),
.B(n_168),
.Y(n_1006)
);

NAND5xp2_ASAP7_75t_L g1007 ( 
.A(n_997),
.B(n_169),
.C(n_171),
.D(n_172),
.E(n_173),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_SL g1008 ( 
.A(n_995),
.B(n_174),
.C(n_175),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_SL g1009 ( 
.A(n_1003),
.B(n_176),
.C(n_177),
.Y(n_1009)
);

OAI211xp5_ASAP7_75t_L g1010 ( 
.A1(n_1002),
.A2(n_902),
.B(n_896),
.C(n_893),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_1007),
.B(n_1000),
.Y(n_1011)
);

AOI211xp5_ASAP7_75t_L g1012 ( 
.A1(n_1006),
.A2(n_999),
.B(n_183),
.C(n_184),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_1008),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_1005),
.B(n_893),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_1009),
.Y(n_1015)
);

OAI22x1_ASAP7_75t_L g1016 ( 
.A1(n_1014),
.A2(n_1011),
.B1(n_1015),
.B2(n_1013),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_1004),
.B1(n_1010),
.B2(n_832),
.Y(n_1017)
);

NOR4xp25_ASAP7_75t_L g1018 ( 
.A(n_1015),
.B(n_182),
.C(n_185),
.D(n_186),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_1011),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_1019),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_1016),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1021),
.A2(n_1018),
.B(n_1017),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_1020),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_1023),
.A2(n_188),
.B(n_189),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1022),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1025),
.Y(n_1026)
);

AOI222xp33_ASAP7_75t_L g1027 ( 
.A1(n_1024),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.C1(n_194),
.C2(n_198),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_1027),
.B(n_200),
.C(n_201),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_SL g1029 ( 
.A1(n_1026),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1028),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.C(n_209),
.Y(n_1030)
);

AOI211xp5_ASAP7_75t_L g1031 ( 
.A1(n_1030),
.A2(n_1029),
.B(n_212),
.C(n_213),
.Y(n_1031)
);


endmodule