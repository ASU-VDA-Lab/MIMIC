module fake_jpeg_7383_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_0),
.C(n_1),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_20),
.B(n_4),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_10),
.B1(n_7),
.B2(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_28),
.B(n_31),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_18),
.C(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_23),
.B1(n_24),
.B2(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_20),
.B1(n_22),
.B2(n_12),
.Y(n_36)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_9),
.B(n_29),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_20),
.B1(n_9),
.B2(n_5),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_36),
.B(n_35),
.C(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_33),
.Y(n_41)
);

AOI21x1_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B(n_38),
.Y(n_43)
);


endmodule