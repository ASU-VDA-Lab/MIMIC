module fake_jpeg_7121_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_58),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_31),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_20),
.B1(n_25),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_63),
.B1(n_23),
.B2(n_30),
.Y(n_74)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_61),
.Y(n_86)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_16),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_75),
.B1(n_84),
.B2(n_16),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_52),
.B(n_55),
.C(n_38),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_80),
.B(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_85),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_37),
.B1(n_35),
.B2(n_46),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_36),
.B1(n_32),
.B2(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_68),
.B1(n_54),
.B2(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_30),
.B1(n_40),
.B2(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_98),
.B1(n_67),
.B2(n_34),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_35),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_0),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_21),
.B1(n_18),
.B2(n_32),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_107),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_110),
.B1(n_122),
.B2(n_76),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_113),
.Y(n_151)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_47),
.B1(n_59),
.B2(n_18),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_123),
.B1(n_93),
.B2(n_99),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_36),
.B(n_21),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_73),
.B(n_86),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_67),
.C(n_26),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_76),
.C(n_84),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_67),
.B1(n_34),
.B2(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_78),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_0),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_156),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_131),
.B(n_143),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_74),
.B1(n_78),
.B2(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_154),
.B1(n_126),
.B2(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_140),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_139),
.B1(n_148),
.B2(n_121),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_95),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_90),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_71),
.C(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_97),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_33),
.B1(n_34),
.B2(n_17),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_89),
.B1(n_87),
.B2(n_85),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_81),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_157),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_82),
.B1(n_72),
.B2(n_77),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_72),
.C(n_70),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_109),
.Y(n_184)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_139),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_112),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_161),
.B(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

OAI22x1_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_127),
.B1(n_152),
.B2(n_128),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_168),
.B1(n_174),
.B2(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_188),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_107),
.B1(n_108),
.B2(n_100),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_185),
.B1(n_135),
.B2(n_131),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_100),
.B1(n_106),
.B2(n_115),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_179),
.B1(n_159),
.B2(n_103),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_115),
.B1(n_118),
.B2(n_113),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_142),
.C(n_83),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_141),
.Y(n_186)
);

AO21x2_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_103),
.B(n_32),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_143),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_33),
.B(n_1),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_0),
.B(n_1),
.Y(n_221)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_198),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_130),
.B1(n_147),
.B2(n_138),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_196),
.A2(n_212),
.B1(n_163),
.B2(n_3),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_140),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_210),
.C(n_219),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_142),
.B(n_33),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_221),
.B(n_162),
.Y(n_223)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_213),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_170),
.B(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_183),
.Y(n_225)
);

BUFx24_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_17),
.B1(n_83),
.B2(n_2),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_17),
.B1(n_83),
.B2(n_3),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_186),
.B1(n_176),
.B2(n_182),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_189),
.C(n_188),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_15),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_189),
.C(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_1),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_196),
.B(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_228),
.B(n_227),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_172),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_232),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_181),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_190),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_191),
.C(n_173),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_209),
.B(n_178),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_247),
.B1(n_203),
.B2(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_216),
.B1(n_201),
.B2(n_200),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_163),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_248),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_15),
.Y(n_248)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_211),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_259),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_194),
.B(n_221),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_269),
.B(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_263),
.C(n_268),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_266),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_194),
.B1(n_201),
.B2(n_217),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_270),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_227),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_206),
.B(n_207),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_277),
.B(n_4),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_245),
.C(n_228),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_5),
.C(n_7),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_223),
.B(n_233),
.C(n_247),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_248),
.C(n_206),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_7),
.C(n_8),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_226),
.B1(n_244),
.B2(n_198),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_286),
.B1(n_287),
.B2(n_265),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_257),
.B(n_215),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_264),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_249),
.A2(n_204),
.B1(n_5),
.B2(n_6),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_264),
.B1(n_251),
.B2(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_293),
.B1(n_285),
.B2(n_276),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_252),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_291),
.C(n_296),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_268),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_271),
.B(n_10),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_9),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_272),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_279),
.B1(n_277),
.B2(n_274),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_307),
.C(n_310),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_289),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_276),
.B1(n_273),
.B2(n_11),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_11),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_303),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_290),
.C(n_299),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_319),
.B(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_13),
.C(n_14),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_7),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_13),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_7),
.B(n_8),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_310),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_311),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_15),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_333),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_324),
.C(n_325),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_327),
.B(n_332),
.C(n_329),
.D(n_320),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_330),
.B(n_8),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_8),
.Y(n_338)
);


endmodule