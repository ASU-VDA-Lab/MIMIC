module fake_ariane_1076_n_777 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_777);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_777;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_84),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_5),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_64),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_57),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_30),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_76),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_77),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_65),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_89),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_35),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_26),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_10),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_22),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_21),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_101),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_55),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_81),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_41),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_102),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_12),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_91),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_118),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_23),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_73),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_6),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_56),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

OAI21x1_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_69),
.B(n_156),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_0),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_167),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_171),
.A2(n_1),
.B(n_2),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_3),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_211),
.Y(n_242)
);

OAI22x1_ASAP7_75t_SL g243 ( 
.A1(n_189),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_7),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_8),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

OAI22x1_ASAP7_75t_R g249 ( 
.A1(n_189),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_163),
.B(n_9),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_163),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_193),
.A2(n_79),
.B(n_155),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_194),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_230),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_219),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_197),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_219),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVxp67_ASAP7_75t_R g277 ( 
.A(n_249),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_R g280 ( 
.A(n_226),
.B(n_164),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_236),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_251),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_242),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_225),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_246),
.B(n_241),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_218),
.B(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_250),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_199),
.B1(n_198),
.B2(n_202),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_251),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_255),
.B(n_170),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_251),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_254),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_224),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_241),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_223),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_244),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_244),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_253),
.C(n_246),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_252),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_262),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_266),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_221),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_285),
.B(n_246),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_286),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_269),
.B(n_221),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_255),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_261),
.B(n_255),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_228),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_275),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_259),
.B(n_228),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_229),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_229),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_234),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_283),
.B(n_222),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_260),
.B(n_222),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_263),
.B(n_222),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_290),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_273),
.B(n_234),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_245),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_245),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_272),
.B(n_227),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_272),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_297),
.A2(n_235),
.B1(n_253),
.B2(n_247),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_247),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_276),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_276),
.B(n_247),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_264),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_265),
.B(n_248),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_248),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_274),
.B(n_256),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_282),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_277),
.B(n_172),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_303),
.B(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_292),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_268),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_221),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_288),
.B(n_248),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_288),
.B(n_248),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_288),
.B(n_180),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_332),
.Y(n_373)
);

NOR2x2_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_243),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_312),
.A2(n_235),
.B1(n_187),
.B2(n_207),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_315),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_258),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_347),
.A2(n_235),
.B1(n_205),
.B2(n_258),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_181),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_217),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_368),
.Y(n_384)
);

NOR2x2_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_11),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_310),
.B(n_184),
.Y(n_388)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_347),
.A2(n_206),
.B1(n_214),
.B2(n_213),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_308),
.B(n_14),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_313),
.B(n_188),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_309),
.A2(n_217),
.B(n_210),
.C(n_209),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_313),
.B(n_196),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_309),
.B(n_201),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

NAND2x2_ASAP7_75t_L g404 ( 
.A(n_323),
.B(n_14),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_203),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

AND2x6_ASAP7_75t_SL g410 ( 
.A(n_358),
.B(n_15),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_204),
.Y(n_411)
);

NAND2x2_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_15),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_345),
.A2(n_321),
.B1(n_318),
.B2(n_365),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_157),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_340),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_327),
.B(n_19),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_20),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_343),
.Y(n_421)
);

AOI21x1_ASAP7_75t_L g422 ( 
.A1(n_339),
.A2(n_24),
.B(n_25),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_340),
.B(n_154),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_355),
.B(n_27),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_324),
.B(n_153),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_345),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_325),
.B(n_152),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_325),
.B(n_32),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_369),
.B(n_33),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_326),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_344),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_346),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_370),
.B(n_151),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_L g439 ( 
.A1(n_363),
.A2(n_38),
.B(n_39),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_362),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_328),
.B(n_40),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_391),
.A2(n_360),
.B1(n_338),
.B2(n_337),
.Y(n_443)
);

BUFx4f_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_390),
.A2(n_330),
.B1(n_354),
.B2(n_348),
.Y(n_446)
);

AO32x1_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_421),
.A3(n_437),
.B1(n_406),
.B2(n_415),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_330),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_330),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_409),
.A2(n_330),
.B1(n_43),
.B2(n_44),
.Y(n_450)
);

BUFx12f_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_438),
.A2(n_330),
.B(n_45),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_42),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_389),
.B(n_46),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_47),
.B(n_48),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_49),
.B(n_50),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_51),
.C(n_52),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_54),
.B(n_59),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_414),
.A2(n_60),
.B(n_61),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_423),
.A2(n_425),
.B(n_442),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_377),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_403),
.B(n_62),
.C(n_63),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_382),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_413),
.B(n_71),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_72),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_407),
.B(n_74),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_428),
.A2(n_75),
.B(n_78),
.C(n_80),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_389),
.B(n_384),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_389),
.B(n_83),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_424),
.A2(n_85),
.B(n_86),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_393),
.B(n_88),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_388),
.B(n_92),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_428),
.A2(n_93),
.B(n_94),
.C(n_96),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_411),
.A2(n_97),
.B1(n_99),
.B2(n_103),
.Y(n_480)
);

O2A1O1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_400),
.A2(n_105),
.B(n_106),
.C(n_109),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_434),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_440),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_436),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_376),
.A2(n_394),
.B(n_395),
.Y(n_486)
);

O2A1O1Ixp5_ASAP7_75t_L g487 ( 
.A1(n_431),
.A2(n_119),
.B(n_120),
.C(n_121),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_376),
.A2(n_125),
.B(n_126),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_379),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_380),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_373),
.A2(n_131),
.B(n_132),
.C(n_133),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_379),
.Y(n_494)
);

BUFx4f_ASAP7_75t_SL g495 ( 
.A(n_418),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_SL g496 ( 
.A(n_439),
.B(n_134),
.C(n_135),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_386),
.B(n_139),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_408),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_452),
.A2(n_422),
.B(n_375),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_399),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_456),
.Y(n_503)
);

INVx3_ASAP7_75t_SL g504 ( 
.A(n_462),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_472),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

AOI22x1_ASAP7_75t_L g508 ( 
.A1(n_461),
.A2(n_435),
.B1(n_398),
.B2(n_397),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_490),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_490),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_486),
.A2(n_375),
.B(n_398),
.Y(n_511)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_496),
.A2(n_378),
.B(n_383),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_445),
.Y(n_514)
);

AO21x1_ASAP7_75t_SL g515 ( 
.A1(n_470),
.A2(n_416),
.B(n_433),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_475),
.A2(n_383),
.B(n_378),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_457),
.A2(n_459),
.B(n_460),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_453),
.A2(n_378),
.B(n_383),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

CKINVDCx12_ASAP7_75t_R g520 ( 
.A(n_477),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_465),
.A2(n_378),
.B1(n_383),
.B2(n_404),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_443),
.B(n_397),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_467),
.B(n_435),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_471),
.A2(n_435),
.B(n_397),
.Y(n_525)
);

OAI21x1_ASAP7_75t_SL g526 ( 
.A1(n_468),
.A2(n_412),
.B(n_410),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_477),
.Y(n_527)
);

AOI21x1_ASAP7_75t_L g528 ( 
.A1(n_478),
.A2(n_140),
.B(n_141),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_492),
.A2(n_144),
.B(n_148),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_494),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_494),
.Y(n_531)
);

BUFx2_ASAP7_75t_R g532 ( 
.A(n_473),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_448),
.A2(n_449),
.B(n_479),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_485),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_487),
.A2(n_150),
.B(n_374),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_485),
.Y(n_536)
);

BUFx4f_ASAP7_75t_L g537 ( 
.A(n_495),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_454),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_469),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_446),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_541),
.A2(n_497),
.B1(n_450),
.B2(n_484),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_541),
.A2(n_482),
.B1(n_463),
.B2(n_466),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_506),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_501),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_540),
.A2(n_458),
.B1(n_480),
.B2(n_493),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_505),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_SL g549 ( 
.A1(n_527),
.A2(n_455),
.B1(n_489),
.B2(n_447),
.Y(n_549)
);

BUFx8_ASAP7_75t_L g550 ( 
.A(n_507),
.Y(n_550)
);

AOI21x1_ASAP7_75t_L g551 ( 
.A1(n_500),
.A2(n_447),
.B(n_481),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_514),
.B(n_523),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_503),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_521),
.Y(n_554)
);

NOR2x1p5_ASAP7_75t_L g555 ( 
.A(n_498),
.B(n_527),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_537),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_506),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_500),
.A2(n_518),
.B(n_533),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_499),
.A2(n_519),
.B1(n_524),
.B2(n_515),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_499),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_522),
.A2(n_499),
.B1(n_538),
.B2(n_537),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_536),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_524),
.A2(n_502),
.B1(n_507),
.B2(n_504),
.Y(n_565)
);

CKINVDCx6p67_ASAP7_75t_R g566 ( 
.A(n_504),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_506),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_506),
.B(n_531),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_530),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_537),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_511),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_525),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_534),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_508),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_536),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_525),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_531),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_530),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_539),
.Y(n_582)
);

OA21x2_ASAP7_75t_L g583 ( 
.A1(n_517),
.A2(n_516),
.B(n_529),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_520),
.A2(n_538),
.B1(n_498),
.B2(n_510),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_532),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_550),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_570),
.B(n_509),
.Y(n_587)
);

CKINVDCx9p33_ASAP7_75t_R g588 ( 
.A(n_550),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_550),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_564),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_566),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_548),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_555),
.B(n_509),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_543),
.A2(n_539),
.B1(n_526),
.B2(n_518),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_556),
.B(n_510),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_539),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_513),
.Y(n_599)
);

NOR2x1p5_ASAP7_75t_L g600 ( 
.A(n_556),
.B(n_528),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_548),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_563),
.B(n_513),
.Y(n_602)
);

AO31x2_ASAP7_75t_L g603 ( 
.A1(n_573),
.A2(n_512),
.A3(n_516),
.B(n_517),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_544),
.A2(n_535),
.B1(n_561),
.B2(n_565),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_SL g605 ( 
.A(n_547),
.B(n_566),
.C(n_579),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_584),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_564),
.B(n_535),
.Y(n_608)
);

AOI221xp5_ASAP7_75t_L g609 ( 
.A1(n_549),
.A2(n_552),
.B1(n_574),
.B2(n_579),
.C(n_572),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_580),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_575),
.B(n_572),
.C(n_583),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_559),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_578),
.B(n_576),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_542),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_568),
.B(n_581),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_R g616 ( 
.A(n_568),
.B(n_567),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_542),
.A2(n_546),
.B1(n_582),
.B2(n_558),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_582),
.A2(n_545),
.B1(n_567),
.B2(n_557),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_568),
.B(n_567),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_582),
.A2(n_558),
.B1(n_577),
.B2(n_571),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_582),
.B(n_545),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_557),
.B(n_560),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_560),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_560),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_582),
.A2(n_545),
.B1(n_557),
.B2(n_569),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_569),
.B(n_558),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_569),
.A2(n_551),
.B1(n_583),
.B2(n_230),
.Y(n_629)
);

AOI211xp5_ASAP7_75t_L g630 ( 
.A1(n_569),
.A2(n_309),
.B(n_540),
.C(n_253),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_569),
.B(n_583),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_R g632 ( 
.A(n_551),
.B(n_353),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_591),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_610),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_628),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_631),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_594),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_608),
.B(n_590),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_593),
.B(n_599),
.Y(n_639)
);

AO31x2_ASAP7_75t_L g640 ( 
.A1(n_604),
.A2(n_614),
.A3(n_612),
.B(n_601),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_624),
.B(n_598),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_606),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_598),
.B(n_623),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_620),
.B(n_613),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_615),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_611),
.B(n_621),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_629),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_603),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_609),
.A2(n_604),
.B1(n_607),
.B2(n_596),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_622),
.B(n_602),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_611),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_630),
.B(n_626),
.Y(n_652)
);

INVx4_ASAP7_75t_SL g653 ( 
.A(n_602),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_617),
.B(n_605),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_627),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_602),
.B(n_627),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_630),
.B(n_597),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_587),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_622),
.B(n_600),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_618),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_622),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_592),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_618),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_595),
.B(n_585),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_662),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_636),
.B(n_586),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_641),
.B(n_589),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_650),
.B(n_616),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_633),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_637),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_657),
.B(n_632),
.C(n_588),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_636),
.B(n_638),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_636),
.B(n_638),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_652),
.B(n_662),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_641),
.B(n_643),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_643),
.B(n_644),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_644),
.B(n_645),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_642),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_639),
.B(n_663),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_662),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_634),
.B(n_655),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_642),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_640),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_650),
.B(n_659),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_640),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_650),
.B(n_659),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_640),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_660),
.B(n_647),
.Y(n_688)
);

NAND2x1_ASAP7_75t_L g689 ( 
.A(n_659),
.B(n_658),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_656),
.B(n_653),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_647),
.B(n_654),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_640),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_654),
.B(n_662),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_634),
.B(n_664),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_672),
.B(n_651),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_672),
.B(n_651),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_678),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_693),
.B(n_662),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_670),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_675),
.B(n_646),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_673),
.B(n_648),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_678),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_677),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_673),
.B(n_648),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_669),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_676),
.B(n_646),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_682),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_675),
.B(n_635),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_666),
.B(n_664),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_676),
.B(n_656),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_681),
.B(n_653),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_666),
.B(n_653),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_694),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_686),
.B(n_653),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_679),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_682),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_715),
.Y(n_718)
);

OAI33xp33_ASAP7_75t_L g719 ( 
.A1(n_700),
.A2(n_691),
.A3(n_688),
.B1(n_671),
.B2(n_687),
.B3(n_683),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_697),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_706),
.B(n_665),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_699),
.Y(n_722)
);

NAND2x2_ASAP7_75t_L g723 ( 
.A(n_708),
.B(n_689),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_713),
.Y(n_724)
);

NAND2x1_ASAP7_75t_L g725 ( 
.A(n_710),
.B(n_684),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_706),
.B(n_674),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_709),
.A2(n_649),
.B(n_674),
.C(n_668),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_699),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_722),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_728),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_727),
.A2(n_705),
.B(n_703),
.Y(n_731)
);

XOR2x2_ASAP7_75t_L g732 ( 
.A(n_725),
.B(n_667),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_718),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_729),
.B(n_724),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_732),
.B(n_717),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_730),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_733),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_735),
.B(n_724),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_737),
.Y(n_739)
);

AOI221xp5_ASAP7_75t_L g740 ( 
.A1(n_734),
.A2(n_719),
.B1(n_731),
.B2(n_695),
.C(n_696),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_734),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_740),
.A2(n_731),
.B(n_738),
.Y(n_742)
);

AO22x1_ASAP7_75t_L g743 ( 
.A1(n_741),
.A2(n_736),
.B1(n_712),
.B2(n_711),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_739),
.A2(n_726),
.B(n_698),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_742),
.B(n_721),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_L g746 ( 
.A1(n_744),
.A2(n_695),
.B(n_696),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_743),
.B(n_712),
.C(n_711),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_742),
.A2(n_723),
.B1(n_701),
.B2(n_704),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_745),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_748),
.B(n_701),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_746),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_747),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_745),
.Y(n_753)
);

AO22x2_ASAP7_75t_L g754 ( 
.A1(n_753),
.A2(n_720),
.B1(n_704),
.B2(n_668),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_749),
.A2(n_752),
.B(n_751),
.Y(n_755)
);

AOI211xp5_ASAP7_75t_L g756 ( 
.A1(n_750),
.A2(n_680),
.B(n_668),
.C(n_714),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_749),
.B(n_716),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_749),
.B(n_707),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_749),
.B(n_707),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_755),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_757),
.B(n_714),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_686),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_754),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_764),
.A2(n_754),
.B1(n_756),
.B2(n_686),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_760),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_762),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_761),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_766),
.A2(n_763),
.B1(n_680),
.B2(n_684),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_768),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_765),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_767),
.B1(n_714),
.B2(n_690),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_772),
.Y(n_773)
);

AOI21x1_ASAP7_75t_L g774 ( 
.A1(n_773),
.A2(n_771),
.B(n_769),
.Y(n_774)
);

OAI211xp5_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_661),
.B(n_692),
.C(n_685),
.Y(n_775)
);

AOI22x1_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_690),
.B1(n_661),
.B2(n_692),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_L g777 ( 
.A1(n_776),
.A2(n_702),
.B1(n_697),
.B2(n_685),
.Y(n_777)
);


endmodule